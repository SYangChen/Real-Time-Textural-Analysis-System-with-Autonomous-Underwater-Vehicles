`timescale 1ns/10ps

module nnctrl_tb ;
	reg			clock, reset ;
	reg			input_signal ;
	reg[31:0]	in ;
	wire		category ;
	// wire[15:0]	cur ;
	
	reg[15:0]	i ;
	
	nnctrl nn ( reset, clock, input_signal, in, category ) ;

	initial // reset、clock
	begin
		clock = 1'b0 ;
		reset = 1'b0 ;
		input_signal = 1'b0 ;
		i = 16'd0 ;
		#10
		reset = 1'b1 ;
		#10
		reset = 1'b0 ;
		
		#100 ;
		in = 32'h003EB2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0046C3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005351 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00559E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005330 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004F54 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004CC4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004BA8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0043D6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003A50 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003E29 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004795 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005430 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00599A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004BFB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00424B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0039C4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0041E1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004C3C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004DAE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003D08 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0039FA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004625 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005922 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005D95 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005D9B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00587E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004F90 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00468F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004304 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00438B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004FFF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0051F5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00559F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006344 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00691B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006504 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006176 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0066C2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00713C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0075F5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006CC4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006AA3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005962 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005A68 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00604B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0060F2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00563F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005585 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006A89 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006ADF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006F5E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007430 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007706 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006B06 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006341 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00655A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00646B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0061C4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006279 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005C86 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005DCA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005860 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00577C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006284 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006480 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0062C7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0068F7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006755 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004BF1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004B86 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0052F8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0056BA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005F0D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005E5F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005A2D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0061BA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0065C1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005D58 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00521E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005235 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0051EC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005A44 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006585 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00690A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00681A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006A1F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005E03 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005CFB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005D65 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005AFC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005B14 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006F1A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0075B9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007859 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00710D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006104 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0054E4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004FD3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005E60 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006C8C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007C98 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008236 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0090D7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008F6A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0098DB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009DE4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A25C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A6A8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AE4F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B7D3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BB88 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B70F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AAAA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0099DA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007922 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006733 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007EE5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009CFE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B104 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B470 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A5E2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00979B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008E48 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008A01 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0079F9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0073A6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007669 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006516 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006BFD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006FB7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0074B6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007987 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007CB9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0074DF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007158 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007255 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007E90 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007FAA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007C63 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0081FE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008456 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008B5D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00862A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007614 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0067E8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007081 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007254 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006CC7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005F43 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00737E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007994 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0083F6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009507 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00969C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009780 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009648 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00929F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008C19 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007E81 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007971 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007348 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006221 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006829 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00753D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00814C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008318 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007BC9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00595D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006373 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007B1F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00811F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009049 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009AB7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00946F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009557 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A24A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A931 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AB01 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0098C5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00959A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009BA6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00997B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0096A2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AE87 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CAF9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CE70 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D3B5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C19F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B3C2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BF71 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C80A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D006 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CD34 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BD58 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A77C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BD5B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BE8F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C79A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CA31 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D3F6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D48B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D1A5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CCFA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B772 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A4D9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00976B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0097A4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008FFB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009A73 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00ADE9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00ADFE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00922A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00794D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0081BF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B1C1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C153 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BE98 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B550 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A754 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A8B0 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AF98 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B0AD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AED4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AD02 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009F51 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008641 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008A93 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008BCE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0089C9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007EFD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007A36 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008580 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A0A4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BA42 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C48A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BA4C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009BE7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009D99 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009859 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009845 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A2C3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B82E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D1B8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D15C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C3B6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A886 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009A6C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007959 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008E27 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008EEC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0082B7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007CCA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009842 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009051 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008331 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0082E6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00821E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00979B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C605 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00DAA1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D1B5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BD23 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BB98 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D002 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D791 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00E570 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00F26C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00F57D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00EA71 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00E098 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D378 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CC61 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B92E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BD34 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C9BA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BFAE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A75F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008774 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00797F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00897D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009415 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00937D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008426 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008975 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009A1D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BA12 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BEBE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BA69 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C06E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C254 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CB3D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CFD4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D3CE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CCBA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B91E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C37A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00DCD4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00FFD2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h01699F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h011930 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h010AA7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00FF32 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0109B8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h010B05 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00FC48 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D0BE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B8BA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BF03 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00DB2D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0105A6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h011D13 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h012179 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h010E4F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D22A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00981F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008001 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009389 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A24A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A12C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A4D8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009769 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008638 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A320 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BE51 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C976 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C2A2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C567 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B0B5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009B5F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0091AC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0096EA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008B1B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0070A2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007D15 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008936 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008F9A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A062 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C6E2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00E4BF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00EEB6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00ED92 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00E580 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00DFE6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C0FF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A57A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A2F5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B1D5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C342 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BE56 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C963 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CE08 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C9DF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AE84 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B459 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BB54 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B252 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AA32 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A61B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008D0C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0084A2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A459 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BACF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BFC3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A8E0 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A965 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AD3D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AA52 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AF8C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B99D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D1BD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00EC7F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00F2E2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00ED45 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D715 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B2FF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009822 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0092B8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008E1D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A09B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A450 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A45D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A598 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A46B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009C78 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009EF6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B258 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D185 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D331 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CE2F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C236 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CEBE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C8E4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C6B8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C7F5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C41C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AD1D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00786F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007F9D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009BCC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AC36 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A9A9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009A09 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006B9E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0076C4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009886 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B258 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AF25 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A97C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A345 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B05B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C82F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00DC36 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00DFAD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D59A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00CCE3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C741 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00DB83 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00F2B5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00F354 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00F134 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00E087 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D5AA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BE86 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009836 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006FE3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00834D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0088BE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0081E7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007FA5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0099AA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AF2E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00ACD7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A1B3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00993A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0097F7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A543 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B4BD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B608 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A421 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008C40 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008664 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009659 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A24D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B3C7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00BEC0 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B819 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A4C5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A584 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A983 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AF98 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00ADA8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009D91 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008102 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007445 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0070B1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007F5A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008888 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008D0B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008ACD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008BFA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00807E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00961B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h014C58 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00915D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00813F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00688E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005B47 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0060B3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0070BA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00861E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0094C8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009969 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B664 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009018 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00883C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008135 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007B8A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0074B8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00746F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0093D4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0098D5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009003 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008368 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007992 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008913 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00955B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A843 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B4F5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00B629 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AC92 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AB7E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AE18 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A99D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AA5A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A00F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A62A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A775 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0095D4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008795 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007F6F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0089F3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009AC8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009D7A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009E81 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009651 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009667 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00911C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008D9C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0089B6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007D1D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006BFB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006E1E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0072AF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007E13 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0085F4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00833E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007888 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006A65 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0079D8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007E99 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008291 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007BE1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00828D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007338 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005958 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006A89 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007C3A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00748A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006EA6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007E00 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008749 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008FBC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00832F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007D93 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008839 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0083F7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007FDB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008A11 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008F10 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0084DD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006937 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005E08 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005921 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00542A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00545D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005BA1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005886 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0045CA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004556 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004564 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0048CE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00527D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005CFD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006721 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007561 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0078C2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008694 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009638 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009FF7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009E0E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0091B5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008841 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007B8A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006CC1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0068E9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006D2F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0059C0 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004E29 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0046B4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005C53 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005F97 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0066F6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00702E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006366 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00516E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0045EC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004778 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004E59 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005717 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0053A5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004FCA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0044E1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003E6A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0038D1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004254 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004CB0 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004EBA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004D49 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004F26 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004406 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003D5E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0037A1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00368F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003C60 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005819 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005F16 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0065A7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0069DD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006576 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005D65 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00663C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006D67 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007320 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00785F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007E78 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007515 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007097 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00595C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0052E4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004C79 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004BAF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003FFE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00475A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0053EB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005D57 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0066C7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006D9D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0065D5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00661E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0066C7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0062F2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00607D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005858 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004238 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003AF5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00379B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0038C2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00336C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004196 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0044D3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0041B2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0037A1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0038AC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003365 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00312E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003894 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003AF7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00382C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003C17 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0035CC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00345B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00363C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003753 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002CFB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00261C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002785 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0013C8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001C9D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002F85 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003AF8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00498C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004974 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004237 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0040DF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00326D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002D8D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002EFB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003F75 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004310 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00422B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003A45 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003477 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003652 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003E2E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0040AA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004911 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004AB5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004FBD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004A80 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004828 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003DCE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004120 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003D2C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003390 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00325A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0038A3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003B78 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003B2A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0032A1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003251 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0028BB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002669 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002F5D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003586 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0038B1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003524 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002F32 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002B8A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001B0F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0015C4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0016CA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001323 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h000DF3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001860 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002390 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002814 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002777 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0023D4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002279 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001DA8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0024DC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002A5E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003236 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0035CE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0030B6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0023DB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001B68 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001D4D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001BA4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001C1F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0022DD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002515 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0025D8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002566 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002E4D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00301F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002BFD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002E2F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002D71 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002C6C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002889 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002B23 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0030DA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002E82 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0026AE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00247D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001F42 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002087 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002E58 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003802 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004301 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0029FE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0026F5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002D27 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003900 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0032BB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003B28 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005BA6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003A6D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00226C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002CA2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0034D9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002D96 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001D95 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0035A2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00274D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00226F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002A82 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004C7F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002A5E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0022ED ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0022BF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0034CD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001880 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0017DF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001CC0 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00105C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001014 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001105 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0014D4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001C85 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0019CD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001AB3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002B47 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00255C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002E11 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003B1A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005087 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002D99 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001D5E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00198D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00168B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001F7D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001D70 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001C38 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001C93 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002000 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0019ED ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001386 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0015FE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00134C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0012BB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0010C1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001187 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0010D5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001CB7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001ACA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001C5F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001B72 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0021E1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h000D7A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001030 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0016E2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h000E5B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001268 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00152A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002413 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0017E0 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0012FE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001B19 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001610 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001719 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00194F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00220B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0019BF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001949 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0012CA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001870 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001DAD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001E33 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002357 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00265F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002B1E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0019BD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002424 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002BD3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002B17 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0025CF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002F5C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00212E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001B34 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001C82 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0023D1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001F04 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0014ED ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00268C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0038E1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00216E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0022A5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003633 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0048FC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003FAB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003065 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003035 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002944 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002346 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001F57 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0021F9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001BD6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001799 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001AB4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002527 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0028DD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001DE2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001BE0 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h001F86 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002A46 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002E13 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002361 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002254 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0033F6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00264E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002F5B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003287 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0029D5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003B1A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002402 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002C03 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002DD5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002742 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004888 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002BD4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003278 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00338A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003598 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004123 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00382D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0055CB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00745B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005B4F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00401B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00294D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003263 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002D02 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00341B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00301F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0033FE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0023A6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002EC1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004885 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0041E3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004057 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003A42 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0043AB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00274E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0041B5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0030DB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003816 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00286A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003740 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0055FE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004AC1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004325 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004FFC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007058 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005DF8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00579B ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008812 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007DA9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007246 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0097C6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0075F7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AE4D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009E2A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006993 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h009301 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005D39 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005223 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00890D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AC02 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0097BC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0072B4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008741 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0084E8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008AE3 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00942C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A695 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C3FB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A095 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A181 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A059 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AD08 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00C482 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00AB14 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00D9FB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00F418 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007B5E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A60A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0079DA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h008B52 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0085A4 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0077AC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00A710 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006C35 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00621A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006ADB ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006CA7 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005DB2 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00642D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006211 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005379 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004BCC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004A87 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00343F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0055CA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0052BF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0064DF ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006CDC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006E38 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0068BA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006225 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007813 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007282 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0074DD ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007813 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006FF6 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0057E8 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h007A99 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0058BA ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0061F5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0063D9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005D65 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0053E5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004670 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004FD5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0051A5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00405C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004424 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006400 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006441 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00687F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005B7C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h006392 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005732 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004954 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00394C ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00510A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004A3E ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00480F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003A6D ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0042D0 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00545F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005A43 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h005572 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003BCC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002800 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0037F1 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003C72 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0035E5 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h0047A9 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004886 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002D9F ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002B31 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h002BAE ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003AAC ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003004 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h00403A ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h004881 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;

		in = 32'h003F60 ;
		input_signal = 1'b1 ;
		#40 ;
		input_signal = 1'b0 ;
		#40 ;


		/*for ( i = 0 ; i < 1000 ; i = i+1 ) begin
			in = 32'hi ;
			input_signal = 1'b1 ;
			#40 ;
			input_signal = 1'b0 ;
			#40 ;
		end*/
		#1000 ;
		// $stop ;
	end
	always #10 clock = clock + 1'b1; 


endmodule