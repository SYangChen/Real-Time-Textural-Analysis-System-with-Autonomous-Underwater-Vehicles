module ROM50( rst, addr, dataOUT1, dataOUT2, dataOUT3, dataOUT4, dataOUT5, dataOUT6, dataOUT7, dataOUT8, dataOUT9, dataOUT10, dataOUT11, dataOUT12, dataOUT13, dataOUT14, dataOUT15, dataOUT16, dataOUT17, dataOUT18, dataOUT19,  dataOUT20, dataOUT21, dataOUT22, dataOUT23, dataOUT24, dataOUT25, dataOUT26, dataOUT27, dataOUT28, dataOUT29, dataOUT30, dataOUT31, dataOUT32, dataOUT33, dataOUT34, dataOUT35, dataOUT36, dataOUT37, dataOUT38, dataOUT39, dataOUT40, dataOUT41, dataOUT42, dataOUT43, dataOUT44, dataOUT45, dataOUT46, dataOUT47, dataOUT48, dataOUT49, dataOUT50, enRead ) ;

	input rst ;
	input [31:0] addr ;	// address to access
	input enRead ;		// enable to read
	output reg [7:0] dataOUT1, dataOUT2, dataOUT3, dataOUT4, dataOUT5, dataOUT6, dataOUT7, dataOUT8, dataOUT9, dataOUT10, dataOUT11, dataOUT12, dataOUT13, dataOUT14, dataOUT15, dataOUT16, dataOUT17, dataOUT18, dataOUT19,  dataOUT20, dataOUT21, dataOUT22, dataOUT23, dataOUT24, dataOUT25, dataOUT26, dataOUT27, dataOUT28, dataOUT29, dataOUT30, dataOUT31, dataOUT32, dataOUT33, dataOUT34, dataOUT35, dataOUT36, dataOUT37, dataOUT38, dataOUT39, dataOUT40, dataOUT41, dataOUT42, dataOUT43, dataOUT44, dataOUT45, dataOUT46, dataOUT47, dataOUT48, dataOUT49, dataOUT50 ;	// output data
	reg[7:0] data [131071:0] ;	// weight
 
	always @(*) begin
		if ( rst ) begin
			data[0] <= 8'h10 ;
			data[1] <= 8'h10 ;
			data[2] <= 8'h10 ;
			data[3] <= 8'h10 ;
			data[4] <= 8'h10 ;
			data[5] <= 8'h10 ;
			data[6] <= 8'h10 ;
			data[7] <= 8'h10 ;
			data[8] <= 8'h10 ;
			data[9] <= 8'h10 ;
			data[10] <= 8'h10 ;
			data[11] <= 8'h10 ;
			data[12] <= 8'h10 ;
			data[13] <= 8'h10 ;
			data[14] <= 8'h10 ;
			data[15] <= 8'h10 ;
			data[16] <= 8'h10 ;
			data[17] <= 8'h10 ;
			data[18] <= 8'h10 ;
			data[19] <= 8'h10 ;
			data[20] <= 8'h10 ;
			data[21] <= 8'h10 ;
			data[22] <= 8'h10 ;
			data[23] <= 8'h10 ;
			data[24] <= 8'h10 ;
			data[25] <= 8'h10 ;
			data[26] <= 8'h10 ;
			data[27] <= 8'h10 ;
			data[28] <= 8'h10 ;
			data[29] <= 8'h10 ;
			data[30] <= 8'h10 ;
			data[31] <= 8'h10 ;
			data[32] <= 8'h10 ;
			data[33] <= 8'h10 ;
			data[34] <= 8'h10 ;
			data[35] <= 8'h10 ;
			data[36] <= 8'h10 ;
			data[37] <= 8'h10 ;
			data[38] <= 8'h10 ;
			data[39] <= 8'h10 ;
			data[40] <= 8'h10 ;
			data[41] <= 8'h10 ;
			data[42] <= 8'h10 ;
			data[43] <= 8'h10 ;
			data[44] <= 8'h10 ;
			data[45] <= 8'h10 ;
			data[46] <= 8'h10 ;
			data[47] <= 8'h10 ;
			data[48] <= 8'h10 ;
			data[49] <= 8'h10 ;
			data[50] <= 8'h10 ;
			data[51] <= 8'h10 ;
			data[52] <= 8'h10 ;
			data[53] <= 8'h10 ;
			data[54] <= 8'h10 ;
			data[55] <= 8'h10 ;
			data[56] <= 8'h10 ;
			data[57] <= 8'h10 ;
			data[58] <= 8'h10 ;
			data[59] <= 8'h10 ;
			data[60] <= 8'h10 ;
			data[61] <= 8'h10 ;
			data[62] <= 8'h10 ;
			data[63] <= 8'h10 ;
			data[64] <= 8'h10 ;
			data[65] <= 8'h10 ;
			data[66] <= 8'h10 ;
			data[67] <= 8'h10 ;
			data[68] <= 8'h10 ;
			data[69] <= 8'h10 ;
			data[70] <= 8'h10 ;
			data[71] <= 8'h10 ;
			data[72] <= 8'h10 ;
			data[73] <= 8'h10 ;
			data[74] <= 8'h10 ;
			data[75] <= 8'h10 ;
			data[76] <= 8'h10 ;
			data[77] <= 8'h10 ;
			data[78] <= 8'h10 ;
			data[79] <= 8'h10 ;
			data[80] <= 8'h10 ;
			data[81] <= 8'h10 ;
			data[82] <= 8'h10 ;
			data[83] <= 8'h10 ;
			data[84] <= 8'h10 ;
			data[85] <= 8'h10 ;
			data[86] <= 8'h10 ;
			data[87] <= 8'h10 ;
			data[88] <= 8'h10 ;
			data[89] <= 8'h10 ;
			data[90] <= 8'h10 ;
			data[91] <= 8'h10 ;
			data[92] <= 8'h10 ;
			data[93] <= 8'h10 ;
			data[94] <= 8'h10 ;
			data[95] <= 8'h10 ;
			data[96] <= 8'h10 ;
			data[97] <= 8'h10 ;
			data[98] <= 8'h10 ;
			data[99] <= 8'h10 ;
			data[100] <= 8'h10 ;
			data[101] <= 8'h10 ;
			data[102] <= 8'h10 ;
			data[103] <= 8'h10 ;
			data[104] <= 8'h10 ;
			data[105] <= 8'h10 ;
			data[106] <= 8'h10 ;
			data[107] <= 8'h10 ;
			data[108] <= 8'h10 ;
			data[109] <= 8'h10 ;
			data[110] <= 8'h10 ;
			data[111] <= 8'h10 ;
			data[112] <= 8'h10 ;
			data[113] <= 8'h10 ;
			data[114] <= 8'h10 ;
			data[115] <= 8'h10 ;
			data[116] <= 8'h10 ;
			data[117] <= 8'h10 ;
			data[118] <= 8'h10 ;
			data[119] <= 8'h10 ;
			data[120] <= 8'h10 ;
			data[121] <= 8'h10 ;
			data[122] <= 8'h10 ;
			data[123] <= 8'h10 ;
			data[124] <= 8'h10 ;
			data[125] <= 8'h10 ;
			data[126] <= 8'h10 ;
			data[127] <= 8'h10 ;
			data[128] <= 8'h10 ;
			data[129] <= 8'h10 ;
			data[130] <= 8'h10 ;
			data[131] <= 8'h10 ;
			data[132] <= 8'h10 ;
			data[133] <= 8'h10 ;
			data[134] <= 8'h10 ;
			data[135] <= 8'h10 ;
			data[136] <= 8'h10 ;
			data[137] <= 8'h10 ;
			data[138] <= 8'h10 ;
			data[139] <= 8'h10 ;
			data[140] <= 8'h10 ;
			data[141] <= 8'h10 ;
			data[142] <= 8'h10 ;
			data[143] <= 8'h10 ;
			data[144] <= 8'h10 ;
			data[145] <= 8'h10 ;
			data[146] <= 8'h10 ;
			data[147] <= 8'h10 ;
			data[148] <= 8'h10 ;
			data[149] <= 8'h10 ;
			data[150] <= 8'h10 ;
			data[151] <= 8'h10 ;
			data[152] <= 8'h10 ;
			data[153] <= 8'h10 ;
			data[154] <= 8'h10 ;
			data[155] <= 8'h10 ;
			data[156] <= 8'h10 ;
			data[157] <= 8'h10 ;
			data[158] <= 8'h10 ;
			data[159] <= 8'h10 ;
			data[160] <= 8'h10 ;
			data[161] <= 8'h10 ;
			data[162] <= 8'h10 ;
			data[163] <= 8'h10 ;
			data[164] <= 8'h10 ;
			data[165] <= 8'h10 ;
			data[166] <= 8'h10 ;
			data[167] <= 8'h10 ;
			data[168] <= 8'h10 ;
			data[169] <= 8'h10 ;
			data[170] <= 8'h10 ;
			data[171] <= 8'h10 ;
			data[172] <= 8'h10 ;
			data[173] <= 8'h10 ;
			data[174] <= 8'h10 ;
			data[175] <= 8'h10 ;
			data[176] <= 8'h10 ;
			data[177] <= 8'h10 ;
			data[178] <= 8'h10 ;
			data[179] <= 8'h10 ;
			data[180] <= 8'h10 ;
			data[181] <= 8'h10 ;
			data[182] <= 8'h10 ;
			data[183] <= 8'h10 ;
			data[184] <= 8'h10 ;
			data[185] <= 8'h10 ;
			data[186] <= 8'h10 ;
			data[187] <= 8'h10 ;
			data[188] <= 8'h10 ;
			data[189] <= 8'h10 ;
			data[190] <= 8'h10 ;
			data[191] <= 8'h10 ;
			data[192] <= 8'h10 ;
			data[193] <= 8'h10 ;
			data[194] <= 8'h10 ;
			data[195] <= 8'h10 ;
			data[196] <= 8'h10 ;
			data[197] <= 8'h10 ;
			data[198] <= 8'h10 ;
			data[199] <= 8'h10 ;
			data[200] <= 8'h10 ;
			data[201] <= 8'h10 ;
			data[202] <= 8'h10 ;
			data[203] <= 8'h10 ;
			data[204] <= 8'h10 ;
			data[205] <= 8'h10 ;
			data[206] <= 8'h10 ;
			data[207] <= 8'h10 ;
			data[208] <= 8'h10 ;
			data[209] <= 8'h10 ;
			data[210] <= 8'h10 ;
			data[211] <= 8'h10 ;
			data[212] <= 8'h10 ;
			data[213] <= 8'h10 ;
			data[214] <= 8'h10 ;
			data[215] <= 8'h10 ;
			data[216] <= 8'h10 ;
			data[217] <= 8'h10 ;
			data[218] <= 8'h10 ;
			data[219] <= 8'h10 ;
			data[220] <= 8'h10 ;
			data[221] <= 8'h10 ;
			data[222] <= 8'h10 ;
			data[223] <= 8'h10 ;
			data[224] <= 8'h10 ;
			data[225] <= 8'h10 ;
			data[226] <= 8'h10 ;
			data[227] <= 8'h10 ;
			data[228] <= 8'h10 ;
			data[229] <= 8'h10 ;
			data[230] <= 8'h10 ;
			data[231] <= 8'h10 ;
			data[232] <= 8'h10 ;
			data[233] <= 8'h10 ;
			data[234] <= 8'h10 ;
			data[235] <= 8'h10 ;
			data[236] <= 8'h10 ;
			data[237] <= 8'h10 ;
			data[238] <= 8'h10 ;
			data[239] <= 8'h10 ;
			data[240] <= 8'h10 ;
			data[241] <= 8'h10 ;
			data[242] <= 8'h10 ;
			data[243] <= 8'h10 ;
			data[244] <= 8'h10 ;
			data[245] <= 8'h10 ;
			data[246] <= 8'h10 ;
			data[247] <= 8'h10 ;
			data[248] <= 8'h10 ;
			data[249] <= 8'h10 ;
			data[250] <= 8'h10 ;
			data[251] <= 8'h10 ;
			data[252] <= 8'h10 ;
			data[253] <= 8'h10 ;
			data[254] <= 8'h10 ;
			data[255] <= 8'h10 ;
			data[256] <= 8'h10 ;
			data[257] <= 8'h10 ;
			data[258] <= 8'h10 ;
			data[259] <= 8'h10 ;
			data[260] <= 8'h10 ;
			data[261] <= 8'h10 ;
			data[262] <= 8'h10 ;
			data[263] <= 8'h10 ;
			data[264] <= 8'h10 ;
			data[265] <= 8'h10 ;
			data[266] <= 8'h10 ;
			data[267] <= 8'h10 ;
			data[268] <= 8'h10 ;
			data[269] <= 8'h10 ;
			data[270] <= 8'h10 ;
			data[271] <= 8'h10 ;
			data[272] <= 8'h10 ;
			data[273] <= 8'h10 ;
			data[274] <= 8'h10 ;
			data[275] <= 8'h10 ;
			data[276] <= 8'h10 ;
			data[277] <= 8'h10 ;
			data[278] <= 8'h10 ;
			data[279] <= 8'h10 ;
			data[280] <= 8'h10 ;
			data[281] <= 8'h10 ;
			data[282] <= 8'h10 ;
			data[283] <= 8'h10 ;
			data[284] <= 8'h10 ;
			data[285] <= 8'h10 ;
			data[286] <= 8'h10 ;
			data[287] <= 8'h10 ;
			data[288] <= 8'h10 ;
			data[289] <= 8'h10 ;
			data[290] <= 8'h10 ;
			data[291] <= 8'h10 ;
			data[292] <= 8'h10 ;
			data[293] <= 8'h10 ;
			data[294] <= 8'h10 ;
			data[295] <= 8'h10 ;
			data[296] <= 8'h10 ;
			data[297] <= 8'h10 ;
			data[298] <= 8'h10 ;
			data[299] <= 8'h10 ;
			data[300] <= 8'h10 ;
			data[301] <= 8'h10 ;
			data[302] <= 8'h10 ;
			data[303] <= 8'h10 ;
			data[304] <= 8'h10 ;
			data[305] <= 8'h10 ;
			data[306] <= 8'h10 ;
			data[307] <= 8'h10 ;
			data[308] <= 8'h10 ;
			data[309] <= 8'h10 ;
			data[310] <= 8'h10 ;
			data[311] <= 8'h10 ;
			data[312] <= 8'h10 ;
			data[313] <= 8'h10 ;
			data[314] <= 8'h10 ;
			data[315] <= 8'h10 ;
			data[316] <= 8'h10 ;
			data[317] <= 8'h10 ;
			data[318] <= 8'h10 ;
			data[319] <= 8'h10 ;
			data[320] <= 8'h10 ;
			data[321] <= 8'h10 ;
			data[322] <= 8'h10 ;
			data[323] <= 8'h10 ;
			data[324] <= 8'h10 ;
			data[325] <= 8'h10 ;
			data[326] <= 8'h10 ;
			data[327] <= 8'h10 ;
			data[328] <= 8'h10 ;
			data[329] <= 8'h10 ;
			data[330] <= 8'h10 ;
			data[331] <= 8'h10 ;
			data[332] <= 8'h10 ;
			data[333] <= 8'h10 ;
			data[334] <= 8'h10 ;
			data[335] <= 8'h10 ;
			data[336] <= 8'h10 ;
			data[337] <= 8'h10 ;
			data[338] <= 8'h10 ;
			data[339] <= 8'h10 ;
			data[340] <= 8'h10 ;
			data[341] <= 8'h10 ;
			data[342] <= 8'h10 ;
			data[343] <= 8'h10 ;
			data[344] <= 8'h10 ;
			data[345] <= 8'h10 ;
			data[346] <= 8'h10 ;
			data[347] <= 8'h10 ;
			data[348] <= 8'h10 ;
			data[349] <= 8'h10 ;
			data[350] <= 8'h10 ;
			data[351] <= 8'h10 ;
			data[352] <= 8'h10 ;
			data[353] <= 8'h10 ;
			data[354] <= 8'h10 ;
			data[355] <= 8'h10 ;
			data[356] <= 8'h10 ;
			data[357] <= 8'h10 ;
			data[358] <= 8'h10 ;
			data[359] <= 8'h10 ;
			data[360] <= 8'h10 ;
			data[361] <= 8'h10 ;
			data[362] <= 8'h10 ;
			data[363] <= 8'h10 ;
			data[364] <= 8'h10 ;
			data[365] <= 8'h10 ;
			data[366] <= 8'h10 ;
			data[367] <= 8'h10 ;
			data[368] <= 8'h10 ;
			data[369] <= 8'h10 ;
			data[370] <= 8'h10 ;
			data[371] <= 8'h10 ;
			data[372] <= 8'h10 ;
			data[373] <= 8'h10 ;
			data[374] <= 8'h10 ;
			data[375] <= 8'h10 ;
			data[376] <= 8'h10 ;
			data[377] <= 8'h10 ;
			data[378] <= 8'h10 ;
			data[379] <= 8'h10 ;
			data[380] <= 8'h10 ;
			data[381] <= 8'h10 ;
			data[382] <= 8'h10 ;
			data[383] <= 8'h10 ;
			data[384] <= 8'h10 ;
			data[385] <= 8'h10 ;
			data[386] <= 8'h10 ;
			data[387] <= 8'h10 ;
			data[388] <= 8'h10 ;
			data[389] <= 8'h10 ;
			data[390] <= 8'h10 ;
			data[391] <= 8'h10 ;
			data[392] <= 8'h10 ;
			data[393] <= 8'h10 ;
			data[394] <= 8'h10 ;
			data[395] <= 8'h10 ;
			data[396] <= 8'h10 ;
			data[397] <= 8'h10 ;
			data[398] <= 8'h10 ;
			data[399] <= 8'h10 ;
			data[400] <= 8'h10 ;
			data[401] <= 8'h10 ;
			data[402] <= 8'h10 ;
			data[403] <= 8'h10 ;
			data[404] <= 8'h10 ;
			data[405] <= 8'h10 ;
			data[406] <= 8'h10 ;
			data[407] <= 8'h10 ;
			data[408] <= 8'h10 ;
			data[409] <= 8'h10 ;
			data[410] <= 8'h10 ;
			data[411] <= 8'h10 ;
			data[412] <= 8'h10 ;
			data[413] <= 8'h10 ;
			data[414] <= 8'h10 ;
			data[415] <= 8'h10 ;
			data[416] <= 8'h10 ;
			data[417] <= 8'h10 ;
			data[418] <= 8'h10 ;
			data[419] <= 8'h10 ;
			data[420] <= 8'h10 ;
			data[421] <= 8'h10 ;
			data[422] <= 8'h10 ;
			data[423] <= 8'h10 ;
			data[424] <= 8'h10 ;
			data[425] <= 8'h10 ;
			data[426] <= 8'h10 ;
			data[427] <= 8'h10 ;
			data[428] <= 8'h10 ;
			data[429] <= 8'h10 ;
			data[430] <= 8'h10 ;
			data[431] <= 8'h10 ;
			data[432] <= 8'h10 ;
			data[433] <= 8'h10 ;
			data[434] <= 8'h10 ;
			data[435] <= 8'h10 ;
			data[436] <= 8'h10 ;
			data[437] <= 8'h10 ;
			data[438] <= 8'h10 ;
			data[439] <= 8'h10 ;
			data[440] <= 8'h10 ;
			data[441] <= 8'h10 ;
			data[442] <= 8'h10 ;
			data[443] <= 8'h10 ;
			data[444] <= 8'h10 ;
			data[445] <= 8'h10 ;
			data[446] <= 8'h10 ;
			data[447] <= 8'h10 ;
			data[448] <= 8'h10 ;
			data[449] <= 8'h10 ;
			data[450] <= 8'h10 ;
			data[451] <= 8'h10 ;
			data[452] <= 8'h10 ;
			data[453] <= 8'h10 ;
			data[454] <= 8'h10 ;
			data[455] <= 8'h10 ;
			data[456] <= 8'h10 ;
			data[457] <= 8'h10 ;
			data[458] <= 8'h10 ;
			data[459] <= 8'h10 ;
			data[460] <= 8'h10 ;
			data[461] <= 8'h10 ;
			data[462] <= 8'h10 ;
			data[463] <= 8'h10 ;
			data[464] <= 8'h10 ;
			data[465] <= 8'h10 ;
			data[466] <= 8'h10 ;
			data[467] <= 8'h10 ;
			data[468] <= 8'h10 ;
			data[469] <= 8'h10 ;
			data[470] <= 8'h10 ;
			data[471] <= 8'h10 ;
			data[472] <= 8'h10 ;
			data[473] <= 8'h10 ;
			data[474] <= 8'h10 ;
			data[475] <= 8'h10 ;
			data[476] <= 8'h10 ;
			data[477] <= 8'h10 ;
			data[478] <= 8'h10 ;
			data[479] <= 8'h10 ;
			data[480] <= 8'h10 ;
			data[481] <= 8'h10 ;
			data[482] <= 8'h10 ;
			data[483] <= 8'h10 ;
			data[484] <= 8'h10 ;
			data[485] <= 8'h10 ;
			data[486] <= 8'h10 ;
			data[487] <= 8'h10 ;
			data[488] <= 8'h10 ;
			data[489] <= 8'h10 ;
			data[490] <= 8'h10 ;
			data[491] <= 8'h10 ;
			data[492] <= 8'h10 ;
			data[493] <= 8'h10 ;
			data[494] <= 8'h10 ;
			data[495] <= 8'h10 ;
			data[496] <= 8'h10 ;
			data[497] <= 8'h10 ;
			data[498] <= 8'h10 ;
			data[499] <= 8'h10 ;
			data[500] <= 8'h10 ;
			data[501] <= 8'h10 ;
			data[502] <= 8'h10 ;
			data[503] <= 8'h10 ;
			data[504] <= 8'h10 ;
			data[505] <= 8'h10 ;
			data[506] <= 8'h10 ;
			data[507] <= 8'h10 ;
			data[508] <= 8'h10 ;
			data[509] <= 8'h10 ;
			data[510] <= 8'h10 ;
			data[511] <= 8'h10 ;
			data[512] <= 8'h10 ;
			data[513] <= 8'h10 ;
			data[514] <= 8'h10 ;
			data[515] <= 8'h10 ;
			data[516] <= 8'h10 ;
			data[517] <= 8'h10 ;
			data[518] <= 8'h10 ;
			data[519] <= 8'h10 ;
			data[520] <= 8'h10 ;
			data[521] <= 8'h10 ;
			data[522] <= 8'h10 ;
			data[523] <= 8'h10 ;
			data[524] <= 8'h10 ;
			data[525] <= 8'h10 ;
			data[526] <= 8'h10 ;
			data[527] <= 8'h10 ;
			data[528] <= 8'h10 ;
			data[529] <= 8'h10 ;
			data[530] <= 8'h10 ;
			data[531] <= 8'h10 ;
			data[532] <= 8'h10 ;
			data[533] <= 8'h10 ;
			data[534] <= 8'h10 ;
			data[535] <= 8'h10 ;
			data[536] <= 8'h10 ;
			data[537] <= 8'h10 ;
			data[538] <= 8'h10 ;
			data[539] <= 8'h10 ;
			data[540] <= 8'h10 ;
			data[541] <= 8'h10 ;
			data[542] <= 8'h10 ;
			data[543] <= 8'h10 ;
			data[544] <= 8'h10 ;
			data[545] <= 8'h10 ;
			data[546] <= 8'h10 ;
			data[547] <= 8'h10 ;
			data[548] <= 8'h10 ;
			data[549] <= 8'h10 ;
			data[550] <= 8'h10 ;
			data[551] <= 8'h10 ;
			data[552] <= 8'h10 ;
			data[553] <= 8'h10 ;
			data[554] <= 8'h10 ;
			data[555] <= 8'h10 ;
			data[556] <= 8'h10 ;
			data[557] <= 8'h10 ;
			data[558] <= 8'h10 ;
			data[559] <= 8'h10 ;
			data[560] <= 8'h10 ;
			data[561] <= 8'h10 ;
			data[562] <= 8'h10 ;
			data[563] <= 8'h10 ;
			data[564] <= 8'h10 ;
			data[565] <= 8'h10 ;
			data[566] <= 8'h10 ;
			data[567] <= 8'h10 ;
			data[568] <= 8'h10 ;
			data[569] <= 8'h10 ;
			data[570] <= 8'h10 ;
			data[571] <= 8'h10 ;
			data[572] <= 8'h10 ;
			data[573] <= 8'h10 ;
			data[574] <= 8'h10 ;
			data[575] <= 8'h10 ;
			data[576] <= 8'h10 ;
			data[577] <= 8'h10 ;
			data[578] <= 8'h10 ;
			data[579] <= 8'h10 ;
			data[580] <= 8'h10 ;
			data[581] <= 8'h10 ;
			data[582] <= 8'h10 ;
			data[583] <= 8'h10 ;
			data[584] <= 8'h10 ;
			data[585] <= 8'h10 ;
			data[586] <= 8'h10 ;
			data[587] <= 8'h10 ;
			data[588] <= 8'h10 ;
			data[589] <= 8'h10 ;
			data[590] <= 8'h10 ;
			data[591] <= 8'h10 ;
			data[592] <= 8'h10 ;
			data[593] <= 8'h10 ;
			data[594] <= 8'h10 ;
			data[595] <= 8'h10 ;
			data[596] <= 8'h10 ;
			data[597] <= 8'h10 ;
			data[598] <= 8'h10 ;
			data[599] <= 8'h10 ;
			data[600] <= 8'h10 ;
			data[601] <= 8'h10 ;
			data[602] <= 8'h10 ;
			data[603] <= 8'h10 ;
			data[604] <= 8'h10 ;
			data[605] <= 8'h10 ;
			data[606] <= 8'h10 ;
			data[607] <= 8'h10 ;
			data[608] <= 8'h10 ;
			data[609] <= 8'h10 ;
			data[610] <= 8'h10 ;
			data[611] <= 8'h10 ;
			data[612] <= 8'h10 ;
			data[613] <= 8'h10 ;
			data[614] <= 8'h10 ;
			data[615] <= 8'h10 ;
			data[616] <= 8'h10 ;
			data[617] <= 8'h10 ;
			data[618] <= 8'h10 ;
			data[619] <= 8'h10 ;
			data[620] <= 8'h10 ;
			data[621] <= 8'h10 ;
			data[622] <= 8'h10 ;
			data[623] <= 8'h10 ;
			data[624] <= 8'h10 ;
			data[625] <= 8'h10 ;
			data[626] <= 8'h10 ;
			data[627] <= 8'h10 ;
			data[628] <= 8'h10 ;
			data[629] <= 8'h10 ;
			data[630] <= 8'h10 ;
			data[631] <= 8'h10 ;
			data[632] <= 8'h10 ;
			data[633] <= 8'h10 ;
			data[634] <= 8'h10 ;
			data[635] <= 8'h10 ;
			data[636] <= 8'h10 ;
			data[637] <= 8'h10 ;
			data[638] <= 8'h10 ;
			data[639] <= 8'h10 ;
			data[640] <= 8'h10 ;
			data[641] <= 8'h10 ;
			data[642] <= 8'h10 ;
			data[643] <= 8'h10 ;
			data[644] <= 8'h10 ;
			data[645] <= 8'h10 ;
			data[646] <= 8'h10 ;
			data[647] <= 8'h10 ;
			data[648] <= 8'h10 ;
			data[649] <= 8'h10 ;
			data[650] <= 8'h10 ;
			data[651] <= 8'h10 ;
			data[652] <= 8'h10 ;
			data[653] <= 8'h10 ;
			data[654] <= 8'h10 ;
			data[655] <= 8'h10 ;
			data[656] <= 8'h10 ;
			data[657] <= 8'h10 ;
			data[658] <= 8'h10 ;
			data[659] <= 8'h10 ;
			data[660] <= 8'h10 ;
			data[661] <= 8'h10 ;
			data[662] <= 8'h10 ;
			data[663] <= 8'h10 ;
			data[664] <= 8'h10 ;
			data[665] <= 8'h10 ;
			data[666] <= 8'h10 ;
			data[667] <= 8'h10 ;
			data[668] <= 8'h10 ;
			data[669] <= 8'h10 ;
			data[670] <= 8'h10 ;
			data[671] <= 8'h10 ;
			data[672] <= 8'h10 ;
			data[673] <= 8'h10 ;
			data[674] <= 8'h10 ;
			data[675] <= 8'h10 ;
			data[676] <= 8'h10 ;
			data[677] <= 8'h10 ;
			data[678] <= 8'h10 ;
			data[679] <= 8'h10 ;
			data[680] <= 8'h10 ;
			data[681] <= 8'h10 ;
			data[682] <= 8'h10 ;
			data[683] <= 8'h10 ;
			data[684] <= 8'h10 ;
			data[685] <= 8'h10 ;
			data[686] <= 8'h10 ;
			data[687] <= 8'h10 ;
			data[688] <= 8'h10 ;
			data[689] <= 8'h10 ;
			data[690] <= 8'h10 ;
			data[691] <= 8'h10 ;
			data[692] <= 8'h10 ;
			data[693] <= 8'h10 ;
			data[694] <= 8'h10 ;
			data[695] <= 8'h10 ;
			data[696] <= 8'h10 ;
			data[697] <= 8'h10 ;
			data[698] <= 8'h10 ;
			data[699] <= 8'h10 ;
			data[700] <= 8'h10 ;
			data[701] <= 8'h10 ;
			data[702] <= 8'h10 ;
			data[703] <= 8'h10 ;
			data[704] <= 8'h10 ;
			data[705] <= 8'h10 ;
			data[706] <= 8'h10 ;
			data[707] <= 8'h10 ;
			data[708] <= 8'h10 ;
			data[709] <= 8'h10 ;
			data[710] <= 8'h10 ;
			data[711] <= 8'h10 ;
			data[712] <= 8'h10 ;
			data[713] <= 8'h10 ;
			data[714] <= 8'h10 ;
			data[715] <= 8'h10 ;
			data[716] <= 8'h10 ;
			data[717] <= 8'h10 ;
			data[718] <= 8'h10 ;
			data[719] <= 8'h10 ;
			data[720] <= 8'h10 ;
			data[721] <= 8'h10 ;
			data[722] <= 8'h10 ;
			data[723] <= 8'h10 ;
			data[724] <= 8'h10 ;
			data[725] <= 8'h10 ;
			data[726] <= 8'h10 ;
			data[727] <= 8'h10 ;
			data[728] <= 8'h10 ;
			data[729] <= 8'h10 ;
			data[730] <= 8'h10 ;
			data[731] <= 8'h10 ;
			data[732] <= 8'h10 ;
			data[733] <= 8'h10 ;
			data[734] <= 8'h10 ;
			data[735] <= 8'h10 ;
			data[736] <= 8'h10 ;
			data[737] <= 8'h10 ;
			data[738] <= 8'h10 ;
			data[739] <= 8'h10 ;
			data[740] <= 8'h10 ;
			data[741] <= 8'h10 ;
			data[742] <= 8'h10 ;
			data[743] <= 8'h10 ;
			data[744] <= 8'h10 ;
			data[745] <= 8'h10 ;
			data[746] <= 8'h10 ;
			data[747] <= 8'h10 ;
			data[748] <= 8'h10 ;
			data[749] <= 8'h10 ;
			data[750] <= 8'h10 ;
			data[751] <= 8'h10 ;
			data[752] <= 8'h10 ;
			data[753] <= 8'h10 ;
			data[754] <= 8'h10 ;
			data[755] <= 8'h10 ;
			data[756] <= 8'h10 ;
			data[757] <= 8'h10 ;
			data[758] <= 8'h10 ;
			data[759] <= 8'h10 ;
			data[760] <= 8'h10 ;
			data[761] <= 8'h10 ;
			data[762] <= 8'h10 ;
			data[763] <= 8'h10 ;
			data[764] <= 8'h10 ;
			data[765] <= 8'h10 ;
			data[766] <= 8'h10 ;
			data[767] <= 8'h10 ;
			data[768] <= 8'h10 ;
			data[769] <= 8'h10 ;
			data[770] <= 8'h10 ;
			data[771] <= 8'h10 ;
			data[772] <= 8'h10 ;
			data[773] <= 8'h10 ;
			data[774] <= 8'h10 ;
			data[775] <= 8'h10 ;
			data[776] <= 8'h10 ;
			data[777] <= 8'h10 ;
			data[778] <= 8'h10 ;
			data[779] <= 8'h10 ;
			data[780] <= 8'h10 ;
			data[781] <= 8'h10 ;
			data[782] <= 8'h10 ;
			data[783] <= 8'h10 ;
			data[784] <= 8'h10 ;
			data[785] <= 8'h10 ;
			data[786] <= 8'h10 ;
			data[787] <= 8'h10 ;
			data[788] <= 8'h10 ;
			data[789] <= 8'h10 ;
			data[790] <= 8'h10 ;
			data[791] <= 8'h10 ;
			data[792] <= 8'h10 ;
			data[793] <= 8'h10 ;
			data[794] <= 8'h10 ;
			data[795] <= 8'h10 ;
			data[796] <= 8'h10 ;
			data[797] <= 8'h10 ;
			data[798] <= 8'h10 ;
			data[799] <= 8'h10 ;
			data[800] <= 8'h10 ;
			data[801] <= 8'h10 ;
			data[802] <= 8'h10 ;
			data[803] <= 8'h10 ;
			data[804] <= 8'h10 ;
			data[805] <= 8'h10 ;
			data[806] <= 8'h10 ;
			data[807] <= 8'h10 ;
			data[808] <= 8'h10 ;
			data[809] <= 8'h10 ;
			data[810] <= 8'h10 ;
			data[811] <= 8'h10 ;
			data[812] <= 8'h10 ;
			data[813] <= 8'h10 ;
			data[814] <= 8'h10 ;
			data[815] <= 8'h10 ;
			data[816] <= 8'h10 ;
			data[817] <= 8'h10 ;
			data[818] <= 8'h10 ;
			data[819] <= 8'h10 ;
			data[820] <= 8'h10 ;
			data[821] <= 8'h10 ;
			data[822] <= 8'h10 ;
			data[823] <= 8'h10 ;
			data[824] <= 8'h10 ;
			data[825] <= 8'h10 ;
			data[826] <= 8'h10 ;
			data[827] <= 8'h10 ;
			data[828] <= 8'h10 ;
			data[829] <= 8'h10 ;
			data[830] <= 8'h10 ;
			data[831] <= 8'h10 ;
			data[832] <= 8'h10 ;
			data[833] <= 8'h10 ;
			data[834] <= 8'h10 ;
			data[835] <= 8'h10 ;
			data[836] <= 8'h10 ;
			data[837] <= 8'h10 ;
			data[838] <= 8'h10 ;
			data[839] <= 8'h10 ;
			data[840] <= 8'h10 ;
			data[841] <= 8'h10 ;
			data[842] <= 8'h10 ;
			data[843] <= 8'h10 ;
			data[844] <= 8'h10 ;
			data[845] <= 8'h10 ;
			data[846] <= 8'h10 ;
			data[847] <= 8'h10 ;
			data[848] <= 8'h10 ;
			data[849] <= 8'h10 ;
			data[850] <= 8'h10 ;
			data[851] <= 8'h10 ;
			data[852] <= 8'h10 ;
			data[853] <= 8'h10 ;
			data[854] <= 8'h10 ;
			data[855] <= 8'h10 ;
			data[856] <= 8'h10 ;
			data[857] <= 8'h10 ;
			data[858] <= 8'h10 ;
			data[859] <= 8'h10 ;
			data[860] <= 8'h10 ;
			data[861] <= 8'h10 ;
			data[862] <= 8'h10 ;
			data[863] <= 8'h10 ;
			data[864] <= 8'h10 ;
			data[865] <= 8'h10 ;
			data[866] <= 8'h10 ;
			data[867] <= 8'h10 ;
			data[868] <= 8'h10 ;
			data[869] <= 8'h10 ;
			data[870] <= 8'h10 ;
			data[871] <= 8'h10 ;
			data[872] <= 8'h10 ;
			data[873] <= 8'h10 ;
			data[874] <= 8'h10 ;
			data[875] <= 8'h10 ;
			data[876] <= 8'h10 ;
			data[877] <= 8'h10 ;
			data[878] <= 8'h10 ;
			data[879] <= 8'h10 ;
			data[880] <= 8'h10 ;
			data[881] <= 8'h10 ;
			data[882] <= 8'h10 ;
			data[883] <= 8'h10 ;
			data[884] <= 8'h10 ;
			data[885] <= 8'h10 ;
			data[886] <= 8'h10 ;
			data[887] <= 8'h10 ;
			data[888] <= 8'h10 ;
			data[889] <= 8'h10 ;
			data[890] <= 8'h10 ;
			data[891] <= 8'h10 ;
			data[892] <= 8'h10 ;
			data[893] <= 8'h10 ;
			data[894] <= 8'h10 ;
			data[895] <= 8'h10 ;
			data[896] <= 8'h10 ;
			data[897] <= 8'h10 ;
			data[898] <= 8'h10 ;
			data[899] <= 8'h10 ;
			data[900] <= 8'h10 ;
			data[901] <= 8'h10 ;
			data[902] <= 8'h10 ;
			data[903] <= 8'h10 ;
			data[904] <= 8'h10 ;
			data[905] <= 8'h10 ;
			data[906] <= 8'h10 ;
			data[907] <= 8'h10 ;
			data[908] <= 8'h10 ;
			data[909] <= 8'h10 ;
			data[910] <= 8'h10 ;
			data[911] <= 8'h10 ;
			data[912] <= 8'h10 ;
			data[913] <= 8'h10 ;
			data[914] <= 8'h10 ;
			data[915] <= 8'h10 ;
			data[916] <= 8'h10 ;
			data[917] <= 8'h10 ;
			data[918] <= 8'h10 ;
			data[919] <= 8'h10 ;
			data[920] <= 8'h10 ;
			data[921] <= 8'h10 ;
			data[922] <= 8'h10 ;
			data[923] <= 8'h10 ;
			data[924] <= 8'h10 ;
			data[925] <= 8'h10 ;
			data[926] <= 8'h10 ;
			data[927] <= 8'h10 ;
			data[928] <= 8'h10 ;
			data[929] <= 8'h10 ;
			data[930] <= 8'h10 ;
			data[931] <= 8'h10 ;
			data[932] <= 8'h10 ;
			data[933] <= 8'h10 ;
			data[934] <= 8'h10 ;
			data[935] <= 8'h10 ;
			data[936] <= 8'h10 ;
			data[937] <= 8'h10 ;
			data[938] <= 8'h10 ;
			data[939] <= 8'h10 ;
			data[940] <= 8'h10 ;
			data[941] <= 8'h10 ;
			data[942] <= 8'h10 ;
			data[943] <= 8'h10 ;
			data[944] <= 8'h10 ;
			data[945] <= 8'h10 ;
			data[946] <= 8'h10 ;
			data[947] <= 8'h10 ;
			data[948] <= 8'h10 ;
			data[949] <= 8'h10 ;
			data[950] <= 8'h10 ;
			data[951] <= 8'h10 ;
			data[952] <= 8'h10 ;
			data[953] <= 8'h10 ;
			data[954] <= 8'h10 ;
			data[955] <= 8'h10 ;
			data[956] <= 8'h10 ;
			data[957] <= 8'h10 ;
			data[958] <= 8'h10 ;
			data[959] <= 8'h10 ;
			data[960] <= 8'h10 ;
			data[961] <= 8'h10 ;
			data[962] <= 8'h10 ;
			data[963] <= 8'h10 ;
			data[964] <= 8'h10 ;
			data[965] <= 8'h10 ;
			data[966] <= 8'h10 ;
			data[967] <= 8'h10 ;
			data[968] <= 8'h10 ;
			data[969] <= 8'h10 ;
			data[970] <= 8'h10 ;
			data[971] <= 8'h10 ;
			data[972] <= 8'h10 ;
			data[973] <= 8'h10 ;
			data[974] <= 8'h10 ;
			data[975] <= 8'h10 ;
			data[976] <= 8'h10 ;
			data[977] <= 8'h10 ;
			data[978] <= 8'h10 ;
			data[979] <= 8'h10 ;
			data[980] <= 8'h10 ;
			data[981] <= 8'h10 ;
			data[982] <= 8'h10 ;
			data[983] <= 8'h10 ;
			data[984] <= 8'h10 ;
			data[985] <= 8'h10 ;
			data[986] <= 8'h10 ;
			data[987] <= 8'h10 ;
			data[988] <= 8'h10 ;
			data[989] <= 8'h10 ;
			data[990] <= 8'h10 ;
			data[991] <= 8'h10 ;
			data[992] <= 8'h10 ;
			data[993] <= 8'h10 ;
			data[994] <= 8'h10 ;
			data[995] <= 8'h10 ;
			data[996] <= 8'h10 ;
			data[997] <= 8'h10 ;
			data[998] <= 8'h10 ;
			data[999] <= 8'h10 ;
			data[1000] <= 8'h10 ;
			data[1001] <= 8'h10 ;
			data[1002] <= 8'h10 ;
			data[1003] <= 8'h10 ;
			data[1004] <= 8'h10 ;
			data[1005] <= 8'h10 ;
			data[1006] <= 8'h10 ;
			data[1007] <= 8'h10 ;
			data[1008] <= 8'h10 ;
			data[1009] <= 8'h10 ;
			data[1010] <= 8'h10 ;
			data[1011] <= 8'h10 ;
			data[1012] <= 8'h10 ;
			data[1013] <= 8'h10 ;
			data[1014] <= 8'h10 ;
			data[1015] <= 8'h10 ;
			data[1016] <= 8'h10 ;
			data[1017] <= 8'h10 ;
			data[1018] <= 8'h10 ;
			data[1019] <= 8'h10 ;
			data[1020] <= 8'h10 ;
			data[1021] <= 8'h10 ;
			data[1022] <= 8'h10 ;
			data[1023] <= 8'h10 ;
			data[1024] <= 8'h10 ;
			data[1025] <= 8'h10 ;
			data[1026] <= 8'h10 ;
			data[1027] <= 8'h10 ;
			data[1028] <= 8'h10 ;
			data[1029] <= 8'h10 ;
			data[1030] <= 8'h10 ;
			data[1031] <= 8'h10 ;
			data[1032] <= 8'h10 ;
			data[1033] <= 8'h10 ;
			data[1034] <= 8'h10 ;
			data[1035] <= 8'h10 ;
			data[1036] <= 8'h10 ;
			data[1037] <= 8'h10 ;
			data[1038] <= 8'h10 ;
			data[1039] <= 8'h10 ;
			data[1040] <= 8'h10 ;
			data[1041] <= 8'h10 ;
			data[1042] <= 8'h10 ;
			data[1043] <= 8'h10 ;
			data[1044] <= 8'h10 ;
			data[1045] <= 8'h10 ;
			data[1046] <= 8'h10 ;
			data[1047] <= 8'h10 ;
			data[1048] <= 8'h10 ;
			data[1049] <= 8'h10 ;
			data[1050] <= 8'h10 ;
			data[1051] <= 8'h10 ;
			data[1052] <= 8'h10 ;
			data[1053] <= 8'h10 ;
			data[1054] <= 8'h10 ;
			data[1055] <= 8'h10 ;
			data[1056] <= 8'h10 ;
			data[1057] <= 8'h10 ;
			data[1058] <= 8'h10 ;
			data[1059] <= 8'h10 ;
			data[1060] <= 8'h10 ;
			data[1061] <= 8'h10 ;
			data[1062] <= 8'h10 ;
			data[1063] <= 8'h10 ;
			data[1064] <= 8'h10 ;
			data[1065] <= 8'h10 ;
			data[1066] <= 8'h10 ;
			data[1067] <= 8'h10 ;
			data[1068] <= 8'h10 ;
			data[1069] <= 8'h10 ;
			data[1070] <= 8'h10 ;
			data[1071] <= 8'h10 ;
			data[1072] <= 8'h10 ;
			data[1073] <= 8'h10 ;
			data[1074] <= 8'h10 ;
			data[1075] <= 8'h10 ;
			data[1076] <= 8'h10 ;
			data[1077] <= 8'h10 ;
			data[1078] <= 8'h10 ;
			data[1079] <= 8'h10 ;
			data[1080] <= 8'h10 ;
			data[1081] <= 8'h10 ;
			data[1082] <= 8'h10 ;
			data[1083] <= 8'h10 ;
			data[1084] <= 8'h10 ;
			data[1085] <= 8'h10 ;
			data[1086] <= 8'h10 ;
			data[1087] <= 8'h10 ;
			data[1088] <= 8'h10 ;
			data[1089] <= 8'h10 ;
			data[1090] <= 8'h10 ;
			data[1091] <= 8'h10 ;
			data[1092] <= 8'h10 ;
			data[1093] <= 8'h10 ;
			data[1094] <= 8'h10 ;
			data[1095] <= 8'h10 ;
			data[1096] <= 8'h10 ;
			data[1097] <= 8'h10 ;
			data[1098] <= 8'h10 ;
			data[1099] <= 8'h10 ;
			data[1100] <= 8'h10 ;
			data[1101] <= 8'h10 ;
			data[1102] <= 8'h10 ;
			data[1103] <= 8'h10 ;
			data[1104] <= 8'h10 ;
			data[1105] <= 8'h10 ;
			data[1106] <= 8'h10 ;
			data[1107] <= 8'h10 ;
			data[1108] <= 8'h10 ;
			data[1109] <= 8'h10 ;
			data[1110] <= 8'h10 ;
			data[1111] <= 8'h10 ;
			data[1112] <= 8'h10 ;
			data[1113] <= 8'h10 ;
			data[1114] <= 8'h10 ;
			data[1115] <= 8'h10 ;
			data[1116] <= 8'h10 ;
			data[1117] <= 8'h10 ;
			data[1118] <= 8'h10 ;
			data[1119] <= 8'h10 ;
			data[1120] <= 8'h10 ;
			data[1121] <= 8'h10 ;
			data[1122] <= 8'h10 ;
			data[1123] <= 8'h10 ;
			data[1124] <= 8'h10 ;
			data[1125] <= 8'h10 ;
			data[1126] <= 8'h10 ;
			data[1127] <= 8'h10 ;
			data[1128] <= 8'h10 ;
			data[1129] <= 8'h10 ;
			data[1130] <= 8'h10 ;
			data[1131] <= 8'h10 ;
			data[1132] <= 8'h10 ;
			data[1133] <= 8'h10 ;
			data[1134] <= 8'h10 ;
			data[1135] <= 8'h10 ;
			data[1136] <= 8'h10 ;
			data[1137] <= 8'h10 ;
			data[1138] <= 8'h10 ;
			data[1139] <= 8'h10 ;
			data[1140] <= 8'h10 ;
			data[1141] <= 8'h10 ;
			data[1142] <= 8'h10 ;
			data[1143] <= 8'h10 ;
			data[1144] <= 8'h10 ;
			data[1145] <= 8'h10 ;
			data[1146] <= 8'h10 ;
			data[1147] <= 8'h10 ;
			data[1148] <= 8'h10 ;
			data[1149] <= 8'h10 ;
			data[1150] <= 8'h10 ;
			data[1151] <= 8'h10 ;
			data[1152] <= 8'h10 ;
			data[1153] <= 8'h10 ;
			data[1154] <= 8'h10 ;
			data[1155] <= 8'h10 ;
			data[1156] <= 8'h10 ;
			data[1157] <= 8'h10 ;
			data[1158] <= 8'h10 ;
			data[1159] <= 8'h10 ;
			data[1160] <= 8'h10 ;
			data[1161] <= 8'h10 ;
			data[1162] <= 8'h10 ;
			data[1163] <= 8'h10 ;
			data[1164] <= 8'h10 ;
			data[1165] <= 8'h10 ;
			data[1166] <= 8'h10 ;
			data[1167] <= 8'h10 ;
			data[1168] <= 8'h10 ;
			data[1169] <= 8'h10 ;
			data[1170] <= 8'h10 ;
			data[1171] <= 8'h10 ;
			data[1172] <= 8'h10 ;
			data[1173] <= 8'h10 ;
			data[1174] <= 8'h10 ;
			data[1175] <= 8'h10 ;
			data[1176] <= 8'h10 ;
			data[1177] <= 8'h10 ;
			data[1178] <= 8'h10 ;
			data[1179] <= 8'h10 ;
			data[1180] <= 8'h10 ;
			data[1181] <= 8'h10 ;
			data[1182] <= 8'h10 ;
			data[1183] <= 8'h10 ;
			data[1184] <= 8'h10 ;
			data[1185] <= 8'h10 ;
			data[1186] <= 8'h10 ;
			data[1187] <= 8'h10 ;
			data[1188] <= 8'h10 ;
			data[1189] <= 8'h10 ;
			data[1190] <= 8'h10 ;
			data[1191] <= 8'h10 ;
			data[1192] <= 8'h10 ;
			data[1193] <= 8'h10 ;
			data[1194] <= 8'h10 ;
			data[1195] <= 8'h10 ;
			data[1196] <= 8'h10 ;
			data[1197] <= 8'h10 ;
			data[1198] <= 8'h10 ;
			data[1199] <= 8'h10 ;
			data[1200] <= 8'h10 ;
			data[1201] <= 8'h10 ;
			data[1202] <= 8'h10 ;
			data[1203] <= 8'h10 ;
			data[1204] <= 8'h10 ;
			data[1205] <= 8'h10 ;
			data[1206] <= 8'h10 ;
			data[1207] <= 8'h10 ;
			data[1208] <= 8'h10 ;
			data[1209] <= 8'h10 ;
			data[1210] <= 8'h10 ;
			data[1211] <= 8'h10 ;
			data[1212] <= 8'h10 ;
			data[1213] <= 8'h10 ;
			data[1214] <= 8'h10 ;
			data[1215] <= 8'h10 ;
			data[1216] <= 8'h10 ;
			data[1217] <= 8'h10 ;
			data[1218] <= 8'h10 ;
			data[1219] <= 8'h10 ;
			data[1220] <= 8'h10 ;
			data[1221] <= 8'h10 ;
			data[1222] <= 8'h10 ;
			data[1223] <= 8'h10 ;
			data[1224] <= 8'h10 ;
			data[1225] <= 8'h10 ;
			data[1226] <= 8'h10 ;
			data[1227] <= 8'h10 ;
			data[1228] <= 8'h10 ;
			data[1229] <= 8'h10 ;
			data[1230] <= 8'h10 ;
			data[1231] <= 8'h10 ;
			data[1232] <= 8'h10 ;
			data[1233] <= 8'h10 ;
			data[1234] <= 8'h10 ;
			data[1235] <= 8'h10 ;
			data[1236] <= 8'h10 ;
			data[1237] <= 8'h10 ;
			data[1238] <= 8'h10 ;
			data[1239] <= 8'h10 ;
			data[1240] <= 8'h10 ;
			data[1241] <= 8'h10 ;
			data[1242] <= 8'h10 ;
			data[1243] <= 8'h10 ;
			data[1244] <= 8'h10 ;
			data[1245] <= 8'h10 ;
			data[1246] <= 8'h10 ;
			data[1247] <= 8'h10 ;
			data[1248] <= 8'h10 ;
			data[1249] <= 8'h10 ;
			data[1250] <= 8'h10 ;
			data[1251] <= 8'h10 ;
			data[1252] <= 8'h10 ;
			data[1253] <= 8'h10 ;
			data[1254] <= 8'h10 ;
			data[1255] <= 8'h10 ;
			data[1256] <= 8'h10 ;
			data[1257] <= 8'h10 ;
			data[1258] <= 8'h10 ;
			data[1259] <= 8'h10 ;
			data[1260] <= 8'h10 ;
			data[1261] <= 8'h10 ;
			data[1262] <= 8'h10 ;
			data[1263] <= 8'h10 ;
			data[1264] <= 8'h10 ;
			data[1265] <= 8'h10 ;
			data[1266] <= 8'h10 ;
			data[1267] <= 8'h10 ;
			data[1268] <= 8'h10 ;
			data[1269] <= 8'h10 ;
			data[1270] <= 8'h10 ;
			data[1271] <= 8'h10 ;
			data[1272] <= 8'h10 ;
			data[1273] <= 8'h10 ;
			data[1274] <= 8'h10 ;
			data[1275] <= 8'h10 ;
			data[1276] <= 8'h10 ;
			data[1277] <= 8'h10 ;
			data[1278] <= 8'h10 ;
			data[1279] <= 8'h10 ;
			data[1280] <= 8'h10 ;
			data[1281] <= 8'h10 ;
			data[1282] <= 8'h10 ;
			data[1283] <= 8'h10 ;
			data[1284] <= 8'h10 ;
			data[1285] <= 8'h10 ;
			data[1286] <= 8'h10 ;
			data[1287] <= 8'h10 ;
			data[1288] <= 8'h10 ;
			data[1289] <= 8'h10 ;
			data[1290] <= 8'h10 ;
			data[1291] <= 8'h10 ;
			data[1292] <= 8'h10 ;
			data[1293] <= 8'h10 ;
			data[1294] <= 8'h10 ;
			data[1295] <= 8'h10 ;
			data[1296] <= 8'h10 ;
			data[1297] <= 8'h10 ;
			data[1298] <= 8'h10 ;
			data[1299] <= 8'h10 ;
			data[1300] <= 8'h10 ;
			data[1301] <= 8'h10 ;
			data[1302] <= 8'h10 ;
			data[1303] <= 8'h10 ;
			data[1304] <= 8'h10 ;
			data[1305] <= 8'h10 ;
			data[1306] <= 8'h10 ;
			data[1307] <= 8'h10 ;
			data[1308] <= 8'h10 ;
			data[1309] <= 8'h10 ;
			data[1310] <= 8'h10 ;
			data[1311] <= 8'h10 ;
			data[1312] <= 8'h10 ;
			data[1313] <= 8'h10 ;
			data[1314] <= 8'h10 ;
			data[1315] <= 8'h10 ;
			data[1316] <= 8'h10 ;
			data[1317] <= 8'h10 ;
			data[1318] <= 8'h10 ;
			data[1319] <= 8'h10 ;
			data[1320] <= 8'h10 ;
			data[1321] <= 8'h10 ;
			data[1322] <= 8'h10 ;
			data[1323] <= 8'h10 ;
			data[1324] <= 8'h10 ;
			data[1325] <= 8'h10 ;
			data[1326] <= 8'h10 ;
			data[1327] <= 8'h10 ;
			data[1328] <= 8'h10 ;
			data[1329] <= 8'h10 ;
			data[1330] <= 8'h10 ;
			data[1331] <= 8'h10 ;
			data[1332] <= 8'h10 ;
			data[1333] <= 8'h10 ;
			data[1334] <= 8'h10 ;
			data[1335] <= 8'h10 ;
			data[1336] <= 8'h10 ;
			data[1337] <= 8'h10 ;
			data[1338] <= 8'h10 ;
			data[1339] <= 8'h10 ;
			data[1340] <= 8'h10 ;
			data[1341] <= 8'h10 ;
			data[1342] <= 8'h10 ;
			data[1343] <= 8'h10 ;
			data[1344] <= 8'h10 ;
			data[1345] <= 8'h10 ;
			data[1346] <= 8'h10 ;
			data[1347] <= 8'h10 ;
			data[1348] <= 8'h10 ;
			data[1349] <= 8'h10 ;
			data[1350] <= 8'h10 ;
			data[1351] <= 8'h10 ;
			data[1352] <= 8'h10 ;
			data[1353] <= 8'h10 ;
			data[1354] <= 8'h10 ;
			data[1355] <= 8'h10 ;
			data[1356] <= 8'h10 ;
			data[1357] <= 8'h10 ;
			data[1358] <= 8'h10 ;
			data[1359] <= 8'h10 ;
			data[1360] <= 8'h10 ;
			data[1361] <= 8'h10 ;
			data[1362] <= 8'h10 ;
			data[1363] <= 8'h10 ;
			data[1364] <= 8'h10 ;
			data[1365] <= 8'h10 ;
			data[1366] <= 8'h10 ;
			data[1367] <= 8'h10 ;
			data[1368] <= 8'h10 ;
			data[1369] <= 8'h10 ;
			data[1370] <= 8'h10 ;
			data[1371] <= 8'h10 ;
			data[1372] <= 8'h10 ;
			data[1373] <= 8'h10 ;
			data[1374] <= 8'h10 ;
			data[1375] <= 8'h10 ;
			data[1376] <= 8'h10 ;
			data[1377] <= 8'h10 ;
			data[1378] <= 8'h10 ;
			data[1379] <= 8'h10 ;
			data[1380] <= 8'h10 ;
			data[1381] <= 8'h10 ;
			data[1382] <= 8'h10 ;
			data[1383] <= 8'h10 ;
			data[1384] <= 8'h10 ;
			data[1385] <= 8'h10 ;
			data[1386] <= 8'h10 ;
			data[1387] <= 8'h10 ;
			data[1388] <= 8'h10 ;
			data[1389] <= 8'h10 ;
			data[1390] <= 8'h10 ;
			data[1391] <= 8'h10 ;
			data[1392] <= 8'h10 ;
			data[1393] <= 8'h10 ;
			data[1394] <= 8'h10 ;
			data[1395] <= 8'h10 ;
			data[1396] <= 8'h10 ;
			data[1397] <= 8'h10 ;
			data[1398] <= 8'h10 ;
			data[1399] <= 8'h10 ;
			data[1400] <= 8'h10 ;
			data[1401] <= 8'h10 ;
			data[1402] <= 8'h10 ;
			data[1403] <= 8'h10 ;
			data[1404] <= 8'h10 ;
			data[1405] <= 8'h10 ;
			data[1406] <= 8'h10 ;
			data[1407] <= 8'h10 ;
			data[1408] <= 8'h10 ;
			data[1409] <= 8'h10 ;
			data[1410] <= 8'h10 ;
			data[1411] <= 8'h10 ;
			data[1412] <= 8'h10 ;
			data[1413] <= 8'h10 ;
			data[1414] <= 8'h10 ;
			data[1415] <= 8'h10 ;
			data[1416] <= 8'h10 ;
			data[1417] <= 8'h10 ;
			data[1418] <= 8'h10 ;
			data[1419] <= 8'h10 ;
			data[1420] <= 8'h10 ;
			data[1421] <= 8'h10 ;
			data[1422] <= 8'h10 ;
			data[1423] <= 8'h10 ;
			data[1424] <= 8'h10 ;
			data[1425] <= 8'h10 ;
			data[1426] <= 8'h10 ;
			data[1427] <= 8'h10 ;
			data[1428] <= 8'h10 ;
			data[1429] <= 8'h10 ;
			data[1430] <= 8'h10 ;
			data[1431] <= 8'h10 ;
			data[1432] <= 8'h10 ;
			data[1433] <= 8'h10 ;
			data[1434] <= 8'h10 ;
			data[1435] <= 8'h10 ;
			data[1436] <= 8'h10 ;
			data[1437] <= 8'h10 ;
			data[1438] <= 8'h10 ;
			data[1439] <= 8'h10 ;
			data[1440] <= 8'h10 ;
			data[1441] <= 8'h10 ;
			data[1442] <= 8'h10 ;
			data[1443] <= 8'h10 ;
			data[1444] <= 8'h10 ;
			data[1445] <= 8'h10 ;
			data[1446] <= 8'h10 ;
			data[1447] <= 8'h10 ;
			data[1448] <= 8'h10 ;
			data[1449] <= 8'h10 ;
			data[1450] <= 8'h10 ;
			data[1451] <= 8'h10 ;
			data[1452] <= 8'h10 ;
			data[1453] <= 8'h10 ;
			data[1454] <= 8'h10 ;
			data[1455] <= 8'h10 ;
			data[1456] <= 8'h10 ;
			data[1457] <= 8'h10 ;
			data[1458] <= 8'h10 ;
			data[1459] <= 8'h10 ;
			data[1460] <= 8'h10 ;
			data[1461] <= 8'h10 ;
			data[1462] <= 8'h10 ;
			data[1463] <= 8'h10 ;
			data[1464] <= 8'h10 ;
			data[1465] <= 8'h10 ;
			data[1466] <= 8'h10 ;
			data[1467] <= 8'h10 ;
			data[1468] <= 8'h10 ;
			data[1469] <= 8'h10 ;
			data[1470] <= 8'h10 ;
			data[1471] <= 8'h10 ;
			data[1472] <= 8'h10 ;
			data[1473] <= 8'h10 ;
			data[1474] <= 8'h10 ;
			data[1475] <= 8'h10 ;
			data[1476] <= 8'h10 ;
			data[1477] <= 8'h10 ;
			data[1478] <= 8'h10 ;
			data[1479] <= 8'h10 ;
			data[1480] <= 8'h10 ;
			data[1481] <= 8'h10 ;
			data[1482] <= 8'h10 ;
			data[1483] <= 8'h10 ;
			data[1484] <= 8'h10 ;
			data[1485] <= 8'h10 ;
			data[1486] <= 8'h10 ;
			data[1487] <= 8'h10 ;
			data[1488] <= 8'h10 ;
			data[1489] <= 8'h10 ;
			data[1490] <= 8'h10 ;
			data[1491] <= 8'h10 ;
			data[1492] <= 8'h10 ;
			data[1493] <= 8'h10 ;
			data[1494] <= 8'h10 ;
			data[1495] <= 8'h10 ;
			data[1496] <= 8'h10 ;
			data[1497] <= 8'h10 ;
			data[1498] <= 8'h10 ;
			data[1499] <= 8'h10 ;
			data[1500] <= 8'h10 ;
			data[1501] <= 8'h10 ;
			data[1502] <= 8'h10 ;
			data[1503] <= 8'h10 ;
			data[1504] <= 8'h10 ;
			data[1505] <= 8'h10 ;
			data[1506] <= 8'h10 ;
			data[1507] <= 8'h10 ;
			data[1508] <= 8'h10 ;
			data[1509] <= 8'h10 ;
			data[1510] <= 8'h10 ;
			data[1511] <= 8'h10 ;
			data[1512] <= 8'h10 ;
			data[1513] <= 8'h10 ;
			data[1514] <= 8'h10 ;
			data[1515] <= 8'h10 ;
			data[1516] <= 8'h10 ;
			data[1517] <= 8'h10 ;
			data[1518] <= 8'h10 ;
			data[1519] <= 8'h10 ;
			data[1520] <= 8'h10 ;
			data[1521] <= 8'h10 ;
			data[1522] <= 8'h10 ;
			data[1523] <= 8'h10 ;
			data[1524] <= 8'h10 ;
			data[1525] <= 8'h10 ;
			data[1526] <= 8'h10 ;
			data[1527] <= 8'h10 ;
			data[1528] <= 8'h10 ;
			data[1529] <= 8'h10 ;
			data[1530] <= 8'h10 ;
			data[1531] <= 8'h10 ;
			data[1532] <= 8'h10 ;
			data[1533] <= 8'h10 ;
			data[1534] <= 8'h10 ;
			data[1535] <= 8'h10 ;
			data[1536] <= 8'h10 ;
			data[1537] <= 8'h10 ;
			data[1538] <= 8'h10 ;
			data[1539] <= 8'h10 ;
			data[1540] <= 8'h10 ;
			data[1541] <= 8'h10 ;
			data[1542] <= 8'h10 ;
			data[1543] <= 8'h10 ;
			data[1544] <= 8'h10 ;
			data[1545] <= 8'h10 ;
			data[1546] <= 8'h10 ;
			data[1547] <= 8'h10 ;
			data[1548] <= 8'h10 ;
			data[1549] <= 8'h10 ;
			data[1550] <= 8'h10 ;
			data[1551] <= 8'h10 ;
			data[1552] <= 8'h10 ;
			data[1553] <= 8'h10 ;
			data[1554] <= 8'h10 ;
			data[1555] <= 8'h10 ;
			data[1556] <= 8'h10 ;
			data[1557] <= 8'h10 ;
			data[1558] <= 8'h10 ;
			data[1559] <= 8'h10 ;
			data[1560] <= 8'h10 ;
			data[1561] <= 8'h10 ;
			data[1562] <= 8'h10 ;
			data[1563] <= 8'h10 ;
			data[1564] <= 8'h10 ;
			data[1565] <= 8'h10 ;
			data[1566] <= 8'h10 ;
			data[1567] <= 8'h10 ;
			data[1568] <= 8'h10 ;
			data[1569] <= 8'h10 ;
			data[1570] <= 8'h10 ;
			data[1571] <= 8'h10 ;
			data[1572] <= 8'h10 ;
			data[1573] <= 8'h10 ;
			data[1574] <= 8'h10 ;
			data[1575] <= 8'h10 ;
			data[1576] <= 8'h10 ;
			data[1577] <= 8'h10 ;
			data[1578] <= 8'h10 ;
			data[1579] <= 8'h10 ;
			data[1580] <= 8'h10 ;
			data[1581] <= 8'h10 ;
			data[1582] <= 8'h10 ;
			data[1583] <= 8'h10 ;
			data[1584] <= 8'h10 ;
			data[1585] <= 8'h10 ;
			data[1586] <= 8'h10 ;
			data[1587] <= 8'h10 ;
			data[1588] <= 8'h10 ;
			data[1589] <= 8'h10 ;
			data[1590] <= 8'h10 ;
			data[1591] <= 8'h10 ;
			data[1592] <= 8'h10 ;
			data[1593] <= 8'h10 ;
			data[1594] <= 8'h10 ;
			data[1595] <= 8'h10 ;
			data[1596] <= 8'h10 ;
			data[1597] <= 8'h10 ;
			data[1598] <= 8'h10 ;
			data[1599] <= 8'h10 ;
			data[1600] <= 8'h10 ;
			data[1601] <= 8'h10 ;
			data[1602] <= 8'h10 ;
			data[1603] <= 8'h10 ;
			data[1604] <= 8'h10 ;
			data[1605] <= 8'h10 ;
			data[1606] <= 8'h10 ;
			data[1607] <= 8'h10 ;
			data[1608] <= 8'h10 ;
			data[1609] <= 8'h10 ;
			data[1610] <= 8'h10 ;
			data[1611] <= 8'h10 ;
			data[1612] <= 8'h10 ;
			data[1613] <= 8'h10 ;
			data[1614] <= 8'h10 ;
			data[1615] <= 8'h10 ;
			data[1616] <= 8'h10 ;
			data[1617] <= 8'h10 ;
			data[1618] <= 8'h10 ;
			data[1619] <= 8'h10 ;
			data[1620] <= 8'h10 ;
			data[1621] <= 8'h10 ;
			data[1622] <= 8'h10 ;
			data[1623] <= 8'h10 ;
			data[1624] <= 8'h10 ;
			data[1625] <= 8'h10 ;
			data[1626] <= 8'h10 ;
			data[1627] <= 8'h10 ;
			data[1628] <= 8'h10 ;
			data[1629] <= 8'h10 ;
			data[1630] <= 8'h10 ;
			data[1631] <= 8'h10 ;
			data[1632] <= 8'h10 ;
			data[1633] <= 8'h10 ;
			data[1634] <= 8'h10 ;
			data[1635] <= 8'h10 ;
			data[1636] <= 8'h10 ;
			data[1637] <= 8'h10 ;
			data[1638] <= 8'h10 ;
			data[1639] <= 8'h10 ;
			data[1640] <= 8'h10 ;
			data[1641] <= 8'h10 ;
			data[1642] <= 8'h10 ;
			data[1643] <= 8'h10 ;
			data[1644] <= 8'h10 ;
			data[1645] <= 8'h10 ;
			data[1646] <= 8'h10 ;
			data[1647] <= 8'h10 ;
			data[1648] <= 8'h10 ;
			data[1649] <= 8'h10 ;
			data[1650] <= 8'h10 ;
			data[1651] <= 8'h10 ;
			data[1652] <= 8'h10 ;
			data[1653] <= 8'h10 ;
			data[1654] <= 8'h10 ;
			data[1655] <= 8'h10 ;
			data[1656] <= 8'h10 ;
			data[1657] <= 8'h10 ;
			data[1658] <= 8'h10 ;
			data[1659] <= 8'h10 ;
			data[1660] <= 8'h10 ;
			data[1661] <= 8'h10 ;
			data[1662] <= 8'h10 ;
			data[1663] <= 8'h10 ;
			data[1664] <= 8'h10 ;
			data[1665] <= 8'h10 ;
			data[1666] <= 8'h10 ;
			data[1667] <= 8'h10 ;
			data[1668] <= 8'h10 ;
			data[1669] <= 8'h10 ;
			data[1670] <= 8'h10 ;
			data[1671] <= 8'h10 ;
			data[1672] <= 8'h10 ;
			data[1673] <= 8'h10 ;
			data[1674] <= 8'h10 ;
			data[1675] <= 8'h10 ;
			data[1676] <= 8'h10 ;
			data[1677] <= 8'h10 ;
			data[1678] <= 8'h10 ;
			data[1679] <= 8'h10 ;
			data[1680] <= 8'h10 ;
			data[1681] <= 8'h10 ;
			data[1682] <= 8'h10 ;
			data[1683] <= 8'h10 ;
			data[1684] <= 8'h10 ;
			data[1685] <= 8'h10 ;
			data[1686] <= 8'h10 ;
			data[1687] <= 8'h10 ;
			data[1688] <= 8'h10 ;
			data[1689] <= 8'h10 ;
			data[1690] <= 8'h10 ;
			data[1691] <= 8'h10 ;
			data[1692] <= 8'h10 ;
			data[1693] <= 8'h10 ;
			data[1694] <= 8'h10 ;
			data[1695] <= 8'h10 ;
			data[1696] <= 8'h10 ;
			data[1697] <= 8'h10 ;
			data[1698] <= 8'h10 ;
			data[1699] <= 8'h10 ;
			data[1700] <= 8'h10 ;
			data[1701] <= 8'h10 ;
			data[1702] <= 8'h10 ;
			data[1703] <= 8'h10 ;
			data[1704] <= 8'h10 ;
			data[1705] <= 8'h10 ;
			data[1706] <= 8'h10 ;
			data[1707] <= 8'h10 ;
			data[1708] <= 8'h10 ;
			data[1709] <= 8'h10 ;
			data[1710] <= 8'h10 ;
			data[1711] <= 8'h10 ;
			data[1712] <= 8'h10 ;
			data[1713] <= 8'h10 ;
			data[1714] <= 8'h10 ;
			data[1715] <= 8'h10 ;
			data[1716] <= 8'h10 ;
			data[1717] <= 8'h10 ;
			data[1718] <= 8'h10 ;
			data[1719] <= 8'h10 ;
			data[1720] <= 8'h10 ;
			data[1721] <= 8'h10 ;
			data[1722] <= 8'h10 ;
			data[1723] <= 8'h10 ;
			data[1724] <= 8'h10 ;
			data[1725] <= 8'h10 ;
			data[1726] <= 8'h10 ;
			data[1727] <= 8'h10 ;
			data[1728] <= 8'h10 ;
			data[1729] <= 8'h10 ;
			data[1730] <= 8'h10 ;
			data[1731] <= 8'h10 ;
			data[1732] <= 8'h10 ;
			data[1733] <= 8'h10 ;
			data[1734] <= 8'h10 ;
			data[1735] <= 8'h10 ;
			data[1736] <= 8'h10 ;
			data[1737] <= 8'h10 ;
			data[1738] <= 8'h10 ;
			data[1739] <= 8'h10 ;
			data[1740] <= 8'h10 ;
			data[1741] <= 8'h10 ;
			data[1742] <= 8'h10 ;
			data[1743] <= 8'h10 ;
			data[1744] <= 8'h10 ;
			data[1745] <= 8'h10 ;
			data[1746] <= 8'h10 ;
			data[1747] <= 8'h10 ;
			data[1748] <= 8'h10 ;
			data[1749] <= 8'h10 ;
			data[1750] <= 8'h10 ;
			data[1751] <= 8'h10 ;
			data[1752] <= 8'h10 ;
			data[1753] <= 8'h10 ;
			data[1754] <= 8'h10 ;
			data[1755] <= 8'h10 ;
			data[1756] <= 8'h10 ;
			data[1757] <= 8'h10 ;
			data[1758] <= 8'h10 ;
			data[1759] <= 8'h10 ;
			data[1760] <= 8'h10 ;
			data[1761] <= 8'h10 ;
			data[1762] <= 8'h10 ;
			data[1763] <= 8'h10 ;
			data[1764] <= 8'h10 ;
			data[1765] <= 8'h10 ;
			data[1766] <= 8'h10 ;
			data[1767] <= 8'h10 ;
			data[1768] <= 8'h10 ;
			data[1769] <= 8'h10 ;
			data[1770] <= 8'h10 ;
			data[1771] <= 8'h10 ;
			data[1772] <= 8'h10 ;
			data[1773] <= 8'h10 ;
			data[1774] <= 8'h10 ;
			data[1775] <= 8'h10 ;
			data[1776] <= 8'h10 ;
			data[1777] <= 8'h10 ;
			data[1778] <= 8'h10 ;
			data[1779] <= 8'h10 ;
			data[1780] <= 8'h10 ;
			data[1781] <= 8'h10 ;
			data[1782] <= 8'h10 ;
			data[1783] <= 8'h10 ;
			data[1784] <= 8'h10 ;
			data[1785] <= 8'h10 ;
			data[1786] <= 8'h10 ;
			data[1787] <= 8'h10 ;
			data[1788] <= 8'h10 ;
			data[1789] <= 8'h10 ;
			data[1790] <= 8'h10 ;
			data[1791] <= 8'h10 ;
			data[1792] <= 8'h10 ;
			data[1793] <= 8'h10 ;
			data[1794] <= 8'h10 ;
			data[1795] <= 8'h10 ;
			data[1796] <= 8'h10 ;
			data[1797] <= 8'h10 ;
			data[1798] <= 8'h10 ;
			data[1799] <= 8'h10 ;
			data[1800] <= 8'h10 ;
			data[1801] <= 8'h10 ;
			data[1802] <= 8'h10 ;
			data[1803] <= 8'h10 ;
			data[1804] <= 8'h10 ;
			data[1805] <= 8'h10 ;
			data[1806] <= 8'h10 ;
			data[1807] <= 8'h10 ;
			data[1808] <= 8'h10 ;
			data[1809] <= 8'h10 ;
			data[1810] <= 8'h10 ;
			data[1811] <= 8'h10 ;
			data[1812] <= 8'h10 ;
			data[1813] <= 8'h10 ;
			data[1814] <= 8'h10 ;
			data[1815] <= 8'h10 ;
			data[1816] <= 8'h10 ;
			data[1817] <= 8'h10 ;
			data[1818] <= 8'h10 ;
			data[1819] <= 8'h10 ;
			data[1820] <= 8'h10 ;
			data[1821] <= 8'h10 ;
			data[1822] <= 8'h10 ;
			data[1823] <= 8'h10 ;
			data[1824] <= 8'h10 ;
			data[1825] <= 8'h10 ;
			data[1826] <= 8'h10 ;
			data[1827] <= 8'h10 ;
			data[1828] <= 8'h10 ;
			data[1829] <= 8'h10 ;
			data[1830] <= 8'h10 ;
			data[1831] <= 8'h10 ;
			data[1832] <= 8'h10 ;
			data[1833] <= 8'h10 ;
			data[1834] <= 8'h10 ;
			data[1835] <= 8'h10 ;
			data[1836] <= 8'h10 ;
			data[1837] <= 8'h10 ;
			data[1838] <= 8'h10 ;
			data[1839] <= 8'h10 ;
			data[1840] <= 8'h10 ;
			data[1841] <= 8'h10 ;
			data[1842] <= 8'h10 ;
			data[1843] <= 8'h10 ;
			data[1844] <= 8'h10 ;
			data[1845] <= 8'h10 ;
			data[1846] <= 8'h10 ;
			data[1847] <= 8'h10 ;
			data[1848] <= 8'h10 ;
			data[1849] <= 8'h10 ;
			data[1850] <= 8'h10 ;
			data[1851] <= 8'h10 ;
			data[1852] <= 8'h10 ;
			data[1853] <= 8'h10 ;
			data[1854] <= 8'h10 ;
			data[1855] <= 8'h10 ;
			data[1856] <= 8'h10 ;
			data[1857] <= 8'h10 ;
			data[1858] <= 8'h10 ;
			data[1859] <= 8'h10 ;
			data[1860] <= 8'h10 ;
			data[1861] <= 8'h10 ;
			data[1862] <= 8'h10 ;
			data[1863] <= 8'h10 ;
			data[1864] <= 8'h10 ;
			data[1865] <= 8'h10 ;
			data[1866] <= 8'h10 ;
			data[1867] <= 8'h10 ;
			data[1868] <= 8'h10 ;
			data[1869] <= 8'h10 ;
			data[1870] <= 8'h10 ;
			data[1871] <= 8'h10 ;
			data[1872] <= 8'h10 ;
			data[1873] <= 8'h10 ;
			data[1874] <= 8'h10 ;
			data[1875] <= 8'h10 ;
			data[1876] <= 8'h10 ;
			data[1877] <= 8'h10 ;
			data[1878] <= 8'h10 ;
			data[1879] <= 8'h10 ;
			data[1880] <= 8'h10 ;
			data[1881] <= 8'h10 ;
			data[1882] <= 8'h10 ;
			data[1883] <= 8'h10 ;
			data[1884] <= 8'h10 ;
			data[1885] <= 8'h10 ;
			data[1886] <= 8'h10 ;
			data[1887] <= 8'h10 ;
			data[1888] <= 8'h10 ;
			data[1889] <= 8'h10 ;
			data[1890] <= 8'h10 ;
			data[1891] <= 8'h10 ;
			data[1892] <= 8'h10 ;
			data[1893] <= 8'h10 ;
			data[1894] <= 8'h10 ;
			data[1895] <= 8'h10 ;
			data[1896] <= 8'h10 ;
			data[1897] <= 8'h10 ;
			data[1898] <= 8'h10 ;
			data[1899] <= 8'h10 ;
			data[1900] <= 8'h10 ;
			data[1901] <= 8'h10 ;
			data[1902] <= 8'h10 ;
			data[1903] <= 8'h10 ;
			data[1904] <= 8'h10 ;
			data[1905] <= 8'h10 ;
			data[1906] <= 8'h10 ;
			data[1907] <= 8'h10 ;
			data[1908] <= 8'h10 ;
			data[1909] <= 8'h10 ;
			data[1910] <= 8'h10 ;
			data[1911] <= 8'h10 ;
			data[1912] <= 8'h10 ;
			data[1913] <= 8'h10 ;
			data[1914] <= 8'h10 ;
			data[1915] <= 8'h10 ;
			data[1916] <= 8'h10 ;
			data[1917] <= 8'h10 ;
			data[1918] <= 8'h10 ;
			data[1919] <= 8'h10 ;
			data[1920] <= 8'h10 ;
			data[1921] <= 8'h10 ;
			data[1922] <= 8'h10 ;
			data[1923] <= 8'h10 ;
			data[1924] <= 8'h10 ;
			data[1925] <= 8'h10 ;
			data[1926] <= 8'h10 ;
			data[1927] <= 8'h10 ;
			data[1928] <= 8'h10 ;
			data[1929] <= 8'h10 ;
			data[1930] <= 8'h10 ;
			data[1931] <= 8'h10 ;
			data[1932] <= 8'h10 ;
			data[1933] <= 8'h10 ;
			data[1934] <= 8'h10 ;
			data[1935] <= 8'h10 ;
			data[1936] <= 8'h10 ;
			data[1937] <= 8'h10 ;
			data[1938] <= 8'h10 ;
			data[1939] <= 8'h10 ;
			data[1940] <= 8'h10 ;
			data[1941] <= 8'h10 ;
			data[1942] <= 8'h10 ;
			data[1943] <= 8'h10 ;
			data[1944] <= 8'h10 ;
			data[1945] <= 8'h10 ;
			data[1946] <= 8'h10 ;
			data[1947] <= 8'h10 ;
			data[1948] <= 8'h10 ;
			data[1949] <= 8'h10 ;
			data[1950] <= 8'h10 ;
			data[1951] <= 8'h10 ;
			data[1952] <= 8'h10 ;
			data[1953] <= 8'h10 ;
			data[1954] <= 8'h10 ;
			data[1955] <= 8'h10 ;
			data[1956] <= 8'h10 ;
			data[1957] <= 8'h10 ;
			data[1958] <= 8'h10 ;
			data[1959] <= 8'h10 ;
			data[1960] <= 8'h10 ;
			data[1961] <= 8'h10 ;
			data[1962] <= 8'h10 ;
			data[1963] <= 8'h10 ;
			data[1964] <= 8'h10 ;
			data[1965] <= 8'h10 ;
			data[1966] <= 8'h10 ;
			data[1967] <= 8'h10 ;
			data[1968] <= 8'h10 ;
			data[1969] <= 8'h10 ;
			data[1970] <= 8'h10 ;
			data[1971] <= 8'h10 ;
			data[1972] <= 8'h10 ;
			data[1973] <= 8'h10 ;
			data[1974] <= 8'h10 ;
			data[1975] <= 8'h10 ;
			data[1976] <= 8'h10 ;
			data[1977] <= 8'h10 ;
			data[1978] <= 8'h10 ;
			data[1979] <= 8'h10 ;
			data[1980] <= 8'h10 ;
			data[1981] <= 8'h10 ;
			data[1982] <= 8'h10 ;
			data[1983] <= 8'h10 ;
			data[1984] <= 8'h10 ;
			data[1985] <= 8'h10 ;
			data[1986] <= 8'h10 ;
			data[1987] <= 8'h10 ;
			data[1988] <= 8'h10 ;
			data[1989] <= 8'h10 ;
			data[1990] <= 8'h10 ;
			data[1991] <= 8'h10 ;
			data[1992] <= 8'h10 ;
			data[1993] <= 8'h10 ;
			data[1994] <= 8'h10 ;
			data[1995] <= 8'h10 ;
			data[1996] <= 8'h10 ;
			data[1997] <= 8'h10 ;
			data[1998] <= 8'h10 ;
			data[1999] <= 8'h10 ;
			data[2000] <= 8'h10 ;
			data[2001] <= 8'h10 ;
			data[2002] <= 8'h10 ;
			data[2003] <= 8'h10 ;
			data[2004] <= 8'h10 ;
			data[2005] <= 8'h10 ;
			data[2006] <= 8'h10 ;
			data[2007] <= 8'h10 ;
			data[2008] <= 8'h10 ;
			data[2009] <= 8'h10 ;
			data[2010] <= 8'h10 ;
			data[2011] <= 8'h10 ;
			data[2012] <= 8'h10 ;
			data[2013] <= 8'h10 ;
			data[2014] <= 8'h10 ;
			data[2015] <= 8'h10 ;
			data[2016] <= 8'h10 ;
			data[2017] <= 8'h10 ;
			data[2018] <= 8'h10 ;
			data[2019] <= 8'h10 ;
			data[2020] <= 8'h10 ;
			data[2021] <= 8'h10 ;
			data[2022] <= 8'h10 ;
			data[2023] <= 8'h10 ;
			data[2024] <= 8'h10 ;
			data[2025] <= 8'h10 ;
			data[2026] <= 8'h10 ;
			data[2027] <= 8'h10 ;
			data[2028] <= 8'h10 ;
			data[2029] <= 8'h10 ;
			data[2030] <= 8'h10 ;
			data[2031] <= 8'h10 ;
			data[2032] <= 8'h10 ;
			data[2033] <= 8'h10 ;
			data[2034] <= 8'h10 ;
			data[2035] <= 8'h10 ;
			data[2036] <= 8'h10 ;
			data[2037] <= 8'h10 ;
			data[2038] <= 8'h10 ;
			data[2039] <= 8'h10 ;
			data[2040] <= 8'h10 ;
			data[2041] <= 8'h10 ;
			data[2042] <= 8'h10 ;
			data[2043] <= 8'h10 ;
			data[2044] <= 8'h10 ;
			data[2045] <= 8'h10 ;
			data[2046] <= 8'h10 ;
			data[2047] <= 8'h10 ;
			data[2048] <= 8'h10 ;
			data[2049] <= 8'h10 ;
			data[2050] <= 8'h10 ;
			data[2051] <= 8'h10 ;
			data[2052] <= 8'h10 ;
			data[2053] <= 8'h10 ;
			data[2054] <= 8'h10 ;
			data[2055] <= 8'h10 ;
			data[2056] <= 8'h10 ;
			data[2057] <= 8'h10 ;
			data[2058] <= 8'h10 ;
			data[2059] <= 8'h10 ;
			data[2060] <= 8'h10 ;
			data[2061] <= 8'h10 ;
			data[2062] <= 8'h10 ;
			data[2063] <= 8'h10 ;
			data[2064] <= 8'h10 ;
			data[2065] <= 8'h10 ;
			data[2066] <= 8'h10 ;
			data[2067] <= 8'h10 ;
			data[2068] <= 8'h10 ;
			data[2069] <= 8'h10 ;
			data[2070] <= 8'h10 ;
			data[2071] <= 8'h10 ;
			data[2072] <= 8'h10 ;
			data[2073] <= 8'h10 ;
			data[2074] <= 8'h10 ;
			data[2075] <= 8'h10 ;
			data[2076] <= 8'h10 ;
			data[2077] <= 8'h10 ;
			data[2078] <= 8'h10 ;
			data[2079] <= 8'h10 ;
			data[2080] <= 8'h10 ;
			data[2081] <= 8'h10 ;
			data[2082] <= 8'h10 ;
			data[2083] <= 8'h10 ;
			data[2084] <= 8'h10 ;
			data[2085] <= 8'h10 ;
			data[2086] <= 8'h10 ;
			data[2087] <= 8'h10 ;
			data[2088] <= 8'h10 ;
			data[2089] <= 8'h10 ;
			data[2090] <= 8'h10 ;
			data[2091] <= 8'h10 ;
			data[2092] <= 8'h10 ;
			data[2093] <= 8'h10 ;
			data[2094] <= 8'h10 ;
			data[2095] <= 8'h10 ;
			data[2096] <= 8'h10 ;
			data[2097] <= 8'h10 ;
			data[2098] <= 8'h10 ;
			data[2099] <= 8'h10 ;
			data[2100] <= 8'h10 ;
			data[2101] <= 8'h10 ;
			data[2102] <= 8'h10 ;
			data[2103] <= 8'h10 ;
			data[2104] <= 8'h10 ;
			data[2105] <= 8'h10 ;
			data[2106] <= 8'h10 ;
			data[2107] <= 8'h10 ;
			data[2108] <= 8'h10 ;
			data[2109] <= 8'h10 ;
			data[2110] <= 8'h10 ;
			data[2111] <= 8'h10 ;
			data[2112] <= 8'h10 ;
			data[2113] <= 8'h10 ;
			data[2114] <= 8'h10 ;
			data[2115] <= 8'h10 ;
			data[2116] <= 8'h10 ;
			data[2117] <= 8'h10 ;
			data[2118] <= 8'h10 ;
			data[2119] <= 8'h10 ;
			data[2120] <= 8'h10 ;
			data[2121] <= 8'h10 ;
			data[2122] <= 8'h10 ;
			data[2123] <= 8'h10 ;
			data[2124] <= 8'h10 ;
			data[2125] <= 8'h10 ;
			data[2126] <= 8'h10 ;
			data[2127] <= 8'h10 ;
			data[2128] <= 8'h10 ;
			data[2129] <= 8'h10 ;
			data[2130] <= 8'h10 ;
			data[2131] <= 8'h10 ;
			data[2132] <= 8'h10 ;
			data[2133] <= 8'h10 ;
			data[2134] <= 8'h10 ;
			data[2135] <= 8'h10 ;
			data[2136] <= 8'h10 ;
			data[2137] <= 8'h10 ;
			data[2138] <= 8'h10 ;
			data[2139] <= 8'h10 ;
			data[2140] <= 8'h10 ;
			data[2141] <= 8'h10 ;
			data[2142] <= 8'h10 ;
			data[2143] <= 8'h10 ;
			data[2144] <= 8'h10 ;
			data[2145] <= 8'h10 ;
			data[2146] <= 8'h10 ;
			data[2147] <= 8'h10 ;
			data[2148] <= 8'h10 ;
			data[2149] <= 8'h10 ;
			data[2150] <= 8'h10 ;
			data[2151] <= 8'h10 ;
			data[2152] <= 8'h10 ;
			data[2153] <= 8'h10 ;
			data[2154] <= 8'h10 ;
			data[2155] <= 8'h10 ;
			data[2156] <= 8'h10 ;
			data[2157] <= 8'h10 ;
			data[2158] <= 8'h10 ;
			data[2159] <= 8'h10 ;
			data[2160] <= 8'h10 ;
			data[2161] <= 8'h10 ;
			data[2162] <= 8'h10 ;
			data[2163] <= 8'h10 ;
			data[2164] <= 8'h10 ;
			data[2165] <= 8'h10 ;
			data[2166] <= 8'h10 ;
			data[2167] <= 8'h10 ;
			data[2168] <= 8'h10 ;
			data[2169] <= 8'h10 ;
			data[2170] <= 8'h10 ;
			data[2171] <= 8'h10 ;
			data[2172] <= 8'h10 ;
			data[2173] <= 8'h10 ;
			data[2174] <= 8'h10 ;
			data[2175] <= 8'h10 ;
			data[2176] <= 8'h10 ;
			data[2177] <= 8'h10 ;
			data[2178] <= 8'h10 ;
			data[2179] <= 8'h10 ;
			data[2180] <= 8'h10 ;
			data[2181] <= 8'h10 ;
			data[2182] <= 8'h10 ;
			data[2183] <= 8'h10 ;
			data[2184] <= 8'h10 ;
			data[2185] <= 8'h10 ;
			data[2186] <= 8'h10 ;
			data[2187] <= 8'h10 ;
			data[2188] <= 8'h10 ;
			data[2189] <= 8'h10 ;
			data[2190] <= 8'h10 ;
			data[2191] <= 8'h10 ;
			data[2192] <= 8'h10 ;
			data[2193] <= 8'h10 ;
			data[2194] <= 8'h10 ;
			data[2195] <= 8'h10 ;
			data[2196] <= 8'h10 ;
			data[2197] <= 8'h10 ;
			data[2198] <= 8'h10 ;
			data[2199] <= 8'h10 ;
			data[2200] <= 8'h10 ;
			data[2201] <= 8'h10 ;
			data[2202] <= 8'h10 ;
			data[2203] <= 8'h10 ;
			data[2204] <= 8'h10 ;
			data[2205] <= 8'h10 ;
			data[2206] <= 8'h10 ;
			data[2207] <= 8'h10 ;
			data[2208] <= 8'h10 ;
			data[2209] <= 8'h10 ;
			data[2210] <= 8'h10 ;
			data[2211] <= 8'h10 ;
			data[2212] <= 8'h10 ;
			data[2213] <= 8'h10 ;
			data[2214] <= 8'h10 ;
			data[2215] <= 8'h10 ;
			data[2216] <= 8'h10 ;
			data[2217] <= 8'h10 ;
			data[2218] <= 8'h10 ;
			data[2219] <= 8'h10 ;
			data[2220] <= 8'h10 ;
			data[2221] <= 8'h10 ;
			data[2222] <= 8'h10 ;
			data[2223] <= 8'h10 ;
			data[2224] <= 8'h10 ;
			data[2225] <= 8'h10 ;
			data[2226] <= 8'h10 ;
			data[2227] <= 8'h10 ;
			data[2228] <= 8'h10 ;
			data[2229] <= 8'h10 ;
			data[2230] <= 8'h10 ;
			data[2231] <= 8'h10 ;
			data[2232] <= 8'h10 ;
			data[2233] <= 8'h10 ;
			data[2234] <= 8'h10 ;
			data[2235] <= 8'h10 ;
			data[2236] <= 8'h10 ;
			data[2237] <= 8'h10 ;
			data[2238] <= 8'h10 ;
			data[2239] <= 8'h10 ;
			data[2240] <= 8'h10 ;
			data[2241] <= 8'h10 ;
			data[2242] <= 8'h10 ;
			data[2243] <= 8'h10 ;
			data[2244] <= 8'h10 ;
			data[2245] <= 8'h10 ;
			data[2246] <= 8'h10 ;
			data[2247] <= 8'h10 ;
			data[2248] <= 8'h10 ;
			data[2249] <= 8'h10 ;
			data[2250] <= 8'h10 ;
			data[2251] <= 8'h10 ;
			data[2252] <= 8'h10 ;
			data[2253] <= 8'h10 ;
			data[2254] <= 8'h10 ;
			data[2255] <= 8'h10 ;
			data[2256] <= 8'h10 ;
			data[2257] <= 8'h10 ;
			data[2258] <= 8'h10 ;
			data[2259] <= 8'h10 ;
			data[2260] <= 8'h10 ;
			data[2261] <= 8'h10 ;
			data[2262] <= 8'h10 ;
			data[2263] <= 8'h10 ;
			data[2264] <= 8'h10 ;
			data[2265] <= 8'h10 ;
			data[2266] <= 8'h10 ;
			data[2267] <= 8'h10 ;
			data[2268] <= 8'h10 ;
			data[2269] <= 8'h10 ;
			data[2270] <= 8'h10 ;
			data[2271] <= 8'h10 ;
			data[2272] <= 8'h10 ;
			data[2273] <= 8'h10 ;
			data[2274] <= 8'h10 ;
			data[2275] <= 8'h10 ;
			data[2276] <= 8'h10 ;
			data[2277] <= 8'h10 ;
			data[2278] <= 8'h10 ;
			data[2279] <= 8'h10 ;
			data[2280] <= 8'h10 ;
			data[2281] <= 8'h10 ;
			data[2282] <= 8'h10 ;
			data[2283] <= 8'h10 ;
			data[2284] <= 8'h10 ;
			data[2285] <= 8'h10 ;
			data[2286] <= 8'h10 ;
			data[2287] <= 8'h10 ;
			data[2288] <= 8'h10 ;
			data[2289] <= 8'h10 ;
			data[2290] <= 8'h10 ;
			data[2291] <= 8'h10 ;
			data[2292] <= 8'h10 ;
			data[2293] <= 8'h10 ;
			data[2294] <= 8'h10 ;
			data[2295] <= 8'h10 ;
			data[2296] <= 8'h10 ;
			data[2297] <= 8'h10 ;
			data[2298] <= 8'h10 ;
			data[2299] <= 8'h10 ;
			data[2300] <= 8'h10 ;
			data[2301] <= 8'h10 ;
			data[2302] <= 8'h10 ;
			data[2303] <= 8'h10 ;
			data[2304] <= 8'h10 ;
			data[2305] <= 8'h10 ;
			data[2306] <= 8'h10 ;
			data[2307] <= 8'h10 ;
			data[2308] <= 8'h10 ;
			data[2309] <= 8'h10 ;
			data[2310] <= 8'h10 ;
			data[2311] <= 8'h10 ;
			data[2312] <= 8'h10 ;
			data[2313] <= 8'h10 ;
			data[2314] <= 8'h10 ;
			data[2315] <= 8'h10 ;
			data[2316] <= 8'h10 ;
			data[2317] <= 8'h10 ;
			data[2318] <= 8'h10 ;
			data[2319] <= 8'h10 ;
			data[2320] <= 8'h10 ;
			data[2321] <= 8'h10 ;
			data[2322] <= 8'h10 ;
			data[2323] <= 8'h10 ;
			data[2324] <= 8'h10 ;
			data[2325] <= 8'h10 ;
			data[2326] <= 8'h10 ;
			data[2327] <= 8'h10 ;
			data[2328] <= 8'h10 ;
			data[2329] <= 8'h10 ;
			data[2330] <= 8'h10 ;
			data[2331] <= 8'h10 ;
			data[2332] <= 8'h10 ;
			data[2333] <= 8'h10 ;
			data[2334] <= 8'h10 ;
			data[2335] <= 8'h10 ;
			data[2336] <= 8'h10 ;
			data[2337] <= 8'h10 ;
			data[2338] <= 8'h10 ;
			data[2339] <= 8'h10 ;
			data[2340] <= 8'h10 ;
			data[2341] <= 8'h10 ;
			data[2342] <= 8'h10 ;
			data[2343] <= 8'h10 ;
			data[2344] <= 8'h10 ;
			data[2345] <= 8'h10 ;
			data[2346] <= 8'h10 ;
			data[2347] <= 8'h10 ;
			data[2348] <= 8'h10 ;
			data[2349] <= 8'h10 ;
			data[2350] <= 8'h10 ;
			data[2351] <= 8'h10 ;
			data[2352] <= 8'h10 ;
			data[2353] <= 8'h10 ;
			data[2354] <= 8'h10 ;
			data[2355] <= 8'h10 ;
			data[2356] <= 8'h10 ;
			data[2357] <= 8'h10 ;
			data[2358] <= 8'h10 ;
			data[2359] <= 8'h10 ;
			data[2360] <= 8'h10 ;
			data[2361] <= 8'h10 ;
			data[2362] <= 8'h10 ;
			data[2363] <= 8'h10 ;
			data[2364] <= 8'h10 ;
			data[2365] <= 8'h10 ;
			data[2366] <= 8'h10 ;
			data[2367] <= 8'h10 ;
			data[2368] <= 8'h10 ;
			data[2369] <= 8'h10 ;
			data[2370] <= 8'h10 ;
			data[2371] <= 8'h10 ;
			data[2372] <= 8'h10 ;
			data[2373] <= 8'h10 ;
			data[2374] <= 8'h10 ;
			data[2375] <= 8'h10 ;
			data[2376] <= 8'h10 ;
			data[2377] <= 8'h10 ;
			data[2378] <= 8'h10 ;
			data[2379] <= 8'h10 ;
			data[2380] <= 8'h10 ;
			data[2381] <= 8'h10 ;
			data[2382] <= 8'h10 ;
			data[2383] <= 8'h10 ;
			data[2384] <= 8'h10 ;
			data[2385] <= 8'h10 ;
			data[2386] <= 8'h10 ;
			data[2387] <= 8'h10 ;
			data[2388] <= 8'h10 ;
			data[2389] <= 8'h10 ;
			data[2390] <= 8'h10 ;
			data[2391] <= 8'h10 ;
			data[2392] <= 8'h10 ;
			data[2393] <= 8'h10 ;
			data[2394] <= 8'h10 ;
			data[2395] <= 8'h10 ;
			data[2396] <= 8'h10 ;
			data[2397] <= 8'h10 ;
			data[2398] <= 8'h10 ;
			data[2399] <= 8'h10 ;
			data[2400] <= 8'h10 ;
			data[2401] <= 8'h10 ;
			data[2402] <= 8'h10 ;
			data[2403] <= 8'h10 ;
			data[2404] <= 8'h10 ;
			data[2405] <= 8'h10 ;
			data[2406] <= 8'h10 ;
			data[2407] <= 8'h10 ;
			data[2408] <= 8'h10 ;
			data[2409] <= 8'h10 ;
			data[2410] <= 8'h10 ;
			data[2411] <= 8'h10 ;
			data[2412] <= 8'h10 ;
			data[2413] <= 8'h10 ;
			data[2414] <= 8'h10 ;
			data[2415] <= 8'h10 ;
			data[2416] <= 8'h10 ;
			data[2417] <= 8'h10 ;
			data[2418] <= 8'h10 ;
			data[2419] <= 8'h10 ;
			data[2420] <= 8'h10 ;
			data[2421] <= 8'h10 ;
			data[2422] <= 8'h10 ;
			data[2423] <= 8'h10 ;
			data[2424] <= 8'h10 ;
			data[2425] <= 8'h10 ;
			data[2426] <= 8'h10 ;
			data[2427] <= 8'h10 ;
			data[2428] <= 8'h10 ;
			data[2429] <= 8'h10 ;
			data[2430] <= 8'h10 ;
			data[2431] <= 8'h10 ;
			data[2432] <= 8'h10 ;
			data[2433] <= 8'h10 ;
			data[2434] <= 8'h10 ;
			data[2435] <= 8'h10 ;
			data[2436] <= 8'h10 ;
			data[2437] <= 8'h10 ;
			data[2438] <= 8'h10 ;
			data[2439] <= 8'h10 ;
			data[2440] <= 8'h10 ;
			data[2441] <= 8'h10 ;
			data[2442] <= 8'h10 ;
			data[2443] <= 8'h10 ;
			data[2444] <= 8'h10 ;
			data[2445] <= 8'h10 ;
			data[2446] <= 8'h10 ;
			data[2447] <= 8'h10 ;
			data[2448] <= 8'h10 ;
			data[2449] <= 8'h10 ;
			data[2450] <= 8'h10 ;
			data[2451] <= 8'h10 ;
			data[2452] <= 8'h10 ;
			data[2453] <= 8'h10 ;
			data[2454] <= 8'h10 ;
			data[2455] <= 8'h10 ;
			data[2456] <= 8'h10 ;
			data[2457] <= 8'h10 ;
			data[2458] <= 8'h10 ;
			data[2459] <= 8'h10 ;
			data[2460] <= 8'h10 ;
			data[2461] <= 8'h10 ;
			data[2462] <= 8'h10 ;
			data[2463] <= 8'h10 ;
			data[2464] <= 8'h10 ;
			data[2465] <= 8'h10 ;
			data[2466] <= 8'h10 ;
			data[2467] <= 8'h10 ;
			data[2468] <= 8'h10 ;
			data[2469] <= 8'h10 ;
			data[2470] <= 8'h10 ;
			data[2471] <= 8'h10 ;
			data[2472] <= 8'h10 ;
			data[2473] <= 8'h10 ;
			data[2474] <= 8'h10 ;
			data[2475] <= 8'h10 ;
			data[2476] <= 8'h10 ;
			data[2477] <= 8'h10 ;
			data[2478] <= 8'h10 ;
			data[2479] <= 8'h10 ;
			data[2480] <= 8'h10 ;
			data[2481] <= 8'h10 ;
			data[2482] <= 8'h10 ;
			data[2483] <= 8'h10 ;
			data[2484] <= 8'h10 ;
			data[2485] <= 8'h10 ;
			data[2486] <= 8'h10 ;
			data[2487] <= 8'h10 ;
			data[2488] <= 8'h10 ;
			data[2489] <= 8'h10 ;
			data[2490] <= 8'h10 ;
			data[2491] <= 8'h10 ;
			data[2492] <= 8'h10 ;
			data[2493] <= 8'h10 ;
			data[2494] <= 8'h10 ;
			data[2495] <= 8'h10 ;
			data[2496] <= 8'h10 ;
			data[2497] <= 8'h10 ;
			data[2498] <= 8'h10 ;
			data[2499] <= 8'h10 ;
			data[2500] <= 8'h10 ;
			data[2501] <= 8'h10 ;
			data[2502] <= 8'h10 ;
			data[2503] <= 8'h10 ;
			data[2504] <= 8'h10 ;
			data[2505] <= 8'h10 ;
			data[2506] <= 8'h10 ;
			data[2507] <= 8'h10 ;
			data[2508] <= 8'h10 ;
			data[2509] <= 8'h10 ;
			data[2510] <= 8'h10 ;
			data[2511] <= 8'h10 ;
			data[2512] <= 8'h10 ;
			data[2513] <= 8'h10 ;
			data[2514] <= 8'h10 ;
			data[2515] <= 8'h10 ;
			data[2516] <= 8'h10 ;
			data[2517] <= 8'h10 ;
			data[2518] <= 8'h10 ;
			data[2519] <= 8'h10 ;
			data[2520] <= 8'h10 ;
			data[2521] <= 8'h10 ;
			data[2522] <= 8'h10 ;
			data[2523] <= 8'h10 ;
			data[2524] <= 8'h10 ;
			data[2525] <= 8'h10 ;
			data[2526] <= 8'h10 ;
			data[2527] <= 8'h10 ;
			data[2528] <= 8'h10 ;
			data[2529] <= 8'h10 ;
			data[2530] <= 8'h10 ;
			data[2531] <= 8'h10 ;
			data[2532] <= 8'h10 ;
			data[2533] <= 8'h10 ;
			data[2534] <= 8'h10 ;
			data[2535] <= 8'h10 ;
			data[2536] <= 8'h10 ;
			data[2537] <= 8'h10 ;
			data[2538] <= 8'h10 ;
			data[2539] <= 8'h10 ;
			data[2540] <= 8'h10 ;
			data[2541] <= 8'h10 ;
			data[2542] <= 8'h10 ;
			data[2543] <= 8'h10 ;
			data[2544] <= 8'h10 ;
			data[2545] <= 8'h10 ;
			data[2546] <= 8'h10 ;
			data[2547] <= 8'h10 ;
			data[2548] <= 8'h10 ;
			data[2549] <= 8'h10 ;
			data[2550] <= 8'h10 ;
			data[2551] <= 8'h10 ;
			data[2552] <= 8'h10 ;
			data[2553] <= 8'h10 ;
			data[2554] <= 8'h10 ;
			data[2555] <= 8'h10 ;
			data[2556] <= 8'h10 ;
			data[2557] <= 8'h10 ;
			data[2558] <= 8'h10 ;
			data[2559] <= 8'h10 ;
			data[2560] <= 8'h10 ;
			data[2561] <= 8'h10 ;
			data[2562] <= 8'h10 ;
			data[2563] <= 8'h10 ;
			data[2564] <= 8'h10 ;
			data[2565] <= 8'h10 ;
			data[2566] <= 8'h10 ;
			data[2567] <= 8'h10 ;
			data[2568] <= 8'h10 ;
			data[2569] <= 8'h10 ;
			data[2570] <= 8'h10 ;
			data[2571] <= 8'h10 ;
			data[2572] <= 8'h10 ;
			data[2573] <= 8'h10 ;
			data[2574] <= 8'h10 ;
			data[2575] <= 8'h10 ;
			data[2576] <= 8'h10 ;
			data[2577] <= 8'h10 ;
			data[2578] <= 8'h10 ;
			data[2579] <= 8'h10 ;
			data[2580] <= 8'h10 ;
			data[2581] <= 8'h10 ;
			data[2582] <= 8'h10 ;
			data[2583] <= 8'h10 ;
			data[2584] <= 8'h10 ;
			data[2585] <= 8'h10 ;
			data[2586] <= 8'h10 ;
			data[2587] <= 8'h10 ;
			data[2588] <= 8'h10 ;
			data[2589] <= 8'h10 ;
			data[2590] <= 8'h10 ;
			data[2591] <= 8'h10 ;
			data[2592] <= 8'h10 ;
			data[2593] <= 8'h10 ;
			data[2594] <= 8'h10 ;
			data[2595] <= 8'h10 ;
			data[2596] <= 8'h10 ;
			data[2597] <= 8'h10 ;
			data[2598] <= 8'h10 ;
			data[2599] <= 8'h10 ;
			data[2600] <= 8'h10 ;
			data[2601] <= 8'h10 ;
			data[2602] <= 8'h10 ;
			data[2603] <= 8'h10 ;
			data[2604] <= 8'h10 ;
			data[2605] <= 8'h10 ;
			data[2606] <= 8'h10 ;
			data[2607] <= 8'h10 ;
			data[2608] <= 8'h10 ;
			data[2609] <= 8'h10 ;
			data[2610] <= 8'h10 ;
			data[2611] <= 8'h10 ;
			data[2612] <= 8'h10 ;
			data[2613] <= 8'h10 ;
			data[2614] <= 8'h10 ;
			data[2615] <= 8'h10 ;
			data[2616] <= 8'h10 ;
			data[2617] <= 8'h10 ;
			data[2618] <= 8'h10 ;
			data[2619] <= 8'h10 ;
			data[2620] <= 8'h10 ;
			data[2621] <= 8'h10 ;
			data[2622] <= 8'h10 ;
			data[2623] <= 8'h10 ;
			data[2624] <= 8'h10 ;
			data[2625] <= 8'h10 ;
			data[2626] <= 8'h10 ;
			data[2627] <= 8'h10 ;
			data[2628] <= 8'h10 ;
			data[2629] <= 8'h10 ;
			data[2630] <= 8'h10 ;
			data[2631] <= 8'h10 ;
			data[2632] <= 8'h10 ;
			data[2633] <= 8'h10 ;
			data[2634] <= 8'h10 ;
			data[2635] <= 8'h10 ;
			data[2636] <= 8'h10 ;
			data[2637] <= 8'h10 ;
			data[2638] <= 8'h10 ;
			data[2639] <= 8'h10 ;
			data[2640] <= 8'h10 ;
			data[2641] <= 8'h10 ;
			data[2642] <= 8'h10 ;
			data[2643] <= 8'h10 ;
			data[2644] <= 8'h10 ;
			data[2645] <= 8'h10 ;
			data[2646] <= 8'h10 ;
			data[2647] <= 8'h10 ;
			data[2648] <= 8'h10 ;
			data[2649] <= 8'h10 ;
			data[2650] <= 8'h10 ;
			data[2651] <= 8'h10 ;
			data[2652] <= 8'h10 ;
			data[2653] <= 8'h10 ;
			data[2654] <= 8'h10 ;
			data[2655] <= 8'h10 ;
			data[2656] <= 8'h10 ;
			data[2657] <= 8'h10 ;
			data[2658] <= 8'h10 ;
			data[2659] <= 8'h10 ;
			data[2660] <= 8'h10 ;
			data[2661] <= 8'h10 ;
			data[2662] <= 8'h10 ;
			data[2663] <= 8'h10 ;
			data[2664] <= 8'h10 ;
			data[2665] <= 8'h10 ;
			data[2666] <= 8'h10 ;
			data[2667] <= 8'h10 ;
			data[2668] <= 8'h10 ;
			data[2669] <= 8'h10 ;
			data[2670] <= 8'h10 ;
			data[2671] <= 8'h10 ;
			data[2672] <= 8'h10 ;
			data[2673] <= 8'h10 ;
			data[2674] <= 8'h10 ;
			data[2675] <= 8'h10 ;
			data[2676] <= 8'h10 ;
			data[2677] <= 8'h10 ;
			data[2678] <= 8'h10 ;
			data[2679] <= 8'h10 ;
			data[2680] <= 8'h10 ;
			data[2681] <= 8'h10 ;
			data[2682] <= 8'h10 ;
			data[2683] <= 8'h10 ;
			data[2684] <= 8'h10 ;
			data[2685] <= 8'h10 ;
			data[2686] <= 8'h10 ;
			data[2687] <= 8'h10 ;
			data[2688] <= 8'h10 ;
			data[2689] <= 8'h10 ;
			data[2690] <= 8'h10 ;
			data[2691] <= 8'h10 ;
			data[2692] <= 8'h10 ;
			data[2693] <= 8'h10 ;
			data[2694] <= 8'h10 ;
			data[2695] <= 8'h10 ;
			data[2696] <= 8'h10 ;
			data[2697] <= 8'h10 ;
			data[2698] <= 8'h10 ;
			data[2699] <= 8'h10 ;
			data[2700] <= 8'h10 ;
			data[2701] <= 8'h10 ;
			data[2702] <= 8'h10 ;
			data[2703] <= 8'h10 ;
			data[2704] <= 8'h10 ;
			data[2705] <= 8'h10 ;
			data[2706] <= 8'h10 ;
			data[2707] <= 8'h10 ;
			data[2708] <= 8'h10 ;
			data[2709] <= 8'h10 ;
			data[2710] <= 8'h10 ;
			data[2711] <= 8'h10 ;
			data[2712] <= 8'h10 ;
			data[2713] <= 8'h10 ;
			data[2714] <= 8'h10 ;
			data[2715] <= 8'h10 ;
			data[2716] <= 8'h10 ;
			data[2717] <= 8'h10 ;
			data[2718] <= 8'h10 ;
			data[2719] <= 8'h10 ;
			data[2720] <= 8'h10 ;
			data[2721] <= 8'h10 ;
			data[2722] <= 8'h10 ;
			data[2723] <= 8'h10 ;
			data[2724] <= 8'h10 ;
			data[2725] <= 8'h10 ;
			data[2726] <= 8'h10 ;
			data[2727] <= 8'h10 ;
			data[2728] <= 8'h10 ;
			data[2729] <= 8'h10 ;
			data[2730] <= 8'h10 ;
			data[2731] <= 8'h10 ;
			data[2732] <= 8'h10 ;
			data[2733] <= 8'h10 ;
			data[2734] <= 8'h10 ;
			data[2735] <= 8'h10 ;
			data[2736] <= 8'h10 ;
			data[2737] <= 8'h10 ;
			data[2738] <= 8'h10 ;
			data[2739] <= 8'h10 ;
			data[2740] <= 8'h10 ;
			data[2741] <= 8'h10 ;
			data[2742] <= 8'h10 ;
			data[2743] <= 8'h10 ;
			data[2744] <= 8'h10 ;
			data[2745] <= 8'h10 ;
			data[2746] <= 8'h10 ;
			data[2747] <= 8'h10 ;
			data[2748] <= 8'h10 ;
			data[2749] <= 8'h10 ;
			data[2750] <= 8'h10 ;
			data[2751] <= 8'h10 ;
			data[2752] <= 8'h10 ;
			data[2753] <= 8'h10 ;
			data[2754] <= 8'h10 ;
			data[2755] <= 8'h10 ;
			data[2756] <= 8'h10 ;
			data[2757] <= 8'h10 ;
			data[2758] <= 8'h10 ;
			data[2759] <= 8'h10 ;
			data[2760] <= 8'h10 ;
			data[2761] <= 8'h10 ;
			data[2762] <= 8'h10 ;
			data[2763] <= 8'h10 ;
			data[2764] <= 8'h10 ;
			data[2765] <= 8'h10 ;
			data[2766] <= 8'h10 ;
			data[2767] <= 8'h10 ;
			data[2768] <= 8'h10 ;
			data[2769] <= 8'h10 ;
			data[2770] <= 8'h10 ;
			data[2771] <= 8'h10 ;
			data[2772] <= 8'h10 ;
			data[2773] <= 8'h10 ;
			data[2774] <= 8'h10 ;
			data[2775] <= 8'h10 ;
			data[2776] <= 8'h10 ;
			data[2777] <= 8'h10 ;
			data[2778] <= 8'h10 ;
			data[2779] <= 8'h10 ;
			data[2780] <= 8'h10 ;
			data[2781] <= 8'h10 ;
			data[2782] <= 8'h10 ;
			data[2783] <= 8'h10 ;
			data[2784] <= 8'h10 ;
			data[2785] <= 8'h10 ;
			data[2786] <= 8'h10 ;
			data[2787] <= 8'h10 ;
			data[2788] <= 8'h10 ;
			data[2789] <= 8'h10 ;
			data[2790] <= 8'h10 ;
			data[2791] <= 8'h10 ;
			data[2792] <= 8'h10 ;
			data[2793] <= 8'h10 ;
			data[2794] <= 8'h10 ;
			data[2795] <= 8'h10 ;
			data[2796] <= 8'h10 ;
			data[2797] <= 8'h10 ;
			data[2798] <= 8'h10 ;
			data[2799] <= 8'h10 ;
			data[2800] <= 8'h10 ;
			data[2801] <= 8'h10 ;
			data[2802] <= 8'h10 ;
			data[2803] <= 8'h10 ;
			data[2804] <= 8'h10 ;
			data[2805] <= 8'h10 ;
			data[2806] <= 8'h10 ;
			data[2807] <= 8'h10 ;
			data[2808] <= 8'h10 ;
			data[2809] <= 8'h10 ;
			data[2810] <= 8'h10 ;
			data[2811] <= 8'h10 ;
			data[2812] <= 8'h10 ;
			data[2813] <= 8'h10 ;
			data[2814] <= 8'h10 ;
			data[2815] <= 8'h10 ;
			data[2816] <= 8'h10 ;
			data[2817] <= 8'h10 ;
			data[2818] <= 8'h10 ;
			data[2819] <= 8'h10 ;
			data[2820] <= 8'h10 ;
			data[2821] <= 8'h10 ;
			data[2822] <= 8'h10 ;
			data[2823] <= 8'h10 ;
			data[2824] <= 8'h10 ;
			data[2825] <= 8'h10 ;
			data[2826] <= 8'h10 ;
			data[2827] <= 8'h10 ;
			data[2828] <= 8'h10 ;
			data[2829] <= 8'h10 ;
			data[2830] <= 8'h10 ;
			data[2831] <= 8'h10 ;
			data[2832] <= 8'h10 ;
			data[2833] <= 8'h10 ;
			data[2834] <= 8'h10 ;
			data[2835] <= 8'h10 ;
			data[2836] <= 8'h10 ;
			data[2837] <= 8'h10 ;
			data[2838] <= 8'h10 ;
			data[2839] <= 8'h10 ;
			data[2840] <= 8'h10 ;
			data[2841] <= 8'h10 ;
			data[2842] <= 8'h10 ;
			data[2843] <= 8'h10 ;
			data[2844] <= 8'h10 ;
			data[2845] <= 8'h10 ;
			data[2846] <= 8'h10 ;
			data[2847] <= 8'h10 ;
			data[2848] <= 8'h10 ;
			data[2849] <= 8'h10 ;
			data[2850] <= 8'h10 ;
			data[2851] <= 8'h10 ;
			data[2852] <= 8'h10 ;
			data[2853] <= 8'h10 ;
			data[2854] <= 8'h10 ;
			data[2855] <= 8'h10 ;
			data[2856] <= 8'h10 ;
			data[2857] <= 8'h10 ;
			data[2858] <= 8'h10 ;
			data[2859] <= 8'h10 ;
			data[2860] <= 8'h10 ;
			data[2861] <= 8'h10 ;
			data[2862] <= 8'h10 ;
			data[2863] <= 8'h10 ;
			data[2864] <= 8'h10 ;
			data[2865] <= 8'h10 ;
			data[2866] <= 8'h10 ;
			data[2867] <= 8'h10 ;
			data[2868] <= 8'h10 ;
			data[2869] <= 8'h10 ;
			data[2870] <= 8'h10 ;
			data[2871] <= 8'h10 ;
			data[2872] <= 8'h10 ;
			data[2873] <= 8'h10 ;
			data[2874] <= 8'h10 ;
			data[2875] <= 8'h10 ;
			data[2876] <= 8'h10 ;
			data[2877] <= 8'h10 ;
			data[2878] <= 8'h10 ;
			data[2879] <= 8'h10 ;
			data[2880] <= 8'h10 ;
			data[2881] <= 8'h10 ;
			data[2882] <= 8'h10 ;
			data[2883] <= 8'h10 ;
			data[2884] <= 8'h10 ;
			data[2885] <= 8'h10 ;
			data[2886] <= 8'h10 ;
			data[2887] <= 8'h10 ;
			data[2888] <= 8'h10 ;
			data[2889] <= 8'h10 ;
			data[2890] <= 8'h10 ;
			data[2891] <= 8'h10 ;
			data[2892] <= 8'h10 ;
			data[2893] <= 8'h10 ;
			data[2894] <= 8'h10 ;
			data[2895] <= 8'h10 ;
			data[2896] <= 8'h10 ;
			data[2897] <= 8'h10 ;
			data[2898] <= 8'h10 ;
			data[2899] <= 8'h10 ;
			data[2900] <= 8'h10 ;
			data[2901] <= 8'h10 ;
			data[2902] <= 8'h10 ;
			data[2903] <= 8'h10 ;
			data[2904] <= 8'h10 ;
			data[2905] <= 8'h10 ;
			data[2906] <= 8'h10 ;
			data[2907] <= 8'h10 ;
			data[2908] <= 8'h10 ;
			data[2909] <= 8'h10 ;
			data[2910] <= 8'h10 ;
			data[2911] <= 8'h10 ;
			data[2912] <= 8'h10 ;
			data[2913] <= 8'h10 ;
			data[2914] <= 8'h10 ;
			data[2915] <= 8'h10 ;
			data[2916] <= 8'h10 ;
			data[2917] <= 8'h10 ;
			data[2918] <= 8'h10 ;
			data[2919] <= 8'h10 ;
			data[2920] <= 8'h10 ;
			data[2921] <= 8'h10 ;
			data[2922] <= 8'h10 ;
			data[2923] <= 8'h10 ;
			data[2924] <= 8'h10 ;
			data[2925] <= 8'h10 ;
			data[2926] <= 8'h10 ;
			data[2927] <= 8'h10 ;
			data[2928] <= 8'h10 ;
			data[2929] <= 8'h10 ;
			data[2930] <= 8'h10 ;
			data[2931] <= 8'h10 ;
			data[2932] <= 8'h10 ;
			data[2933] <= 8'h10 ;
			data[2934] <= 8'h10 ;
			data[2935] <= 8'h10 ;
			data[2936] <= 8'h10 ;
			data[2937] <= 8'h10 ;
			data[2938] <= 8'h10 ;
			data[2939] <= 8'h10 ;
			data[2940] <= 8'h10 ;
			data[2941] <= 8'h10 ;
			data[2942] <= 8'h10 ;
			data[2943] <= 8'h10 ;
			data[2944] <= 8'h10 ;
			data[2945] <= 8'h10 ;
			data[2946] <= 8'h10 ;
			data[2947] <= 8'h10 ;
			data[2948] <= 8'h10 ;
			data[2949] <= 8'h10 ;
			data[2950] <= 8'h10 ;
			data[2951] <= 8'h10 ;
			data[2952] <= 8'h10 ;
			data[2953] <= 8'h10 ;
			data[2954] <= 8'h10 ;
			data[2955] <= 8'h10 ;
			data[2956] <= 8'h10 ;
			data[2957] <= 8'h10 ;
			data[2958] <= 8'h10 ;
			data[2959] <= 8'h10 ;
			data[2960] <= 8'h10 ;
			data[2961] <= 8'h10 ;
			data[2962] <= 8'h10 ;
			data[2963] <= 8'h10 ;
			data[2964] <= 8'h10 ;
			data[2965] <= 8'h10 ;
			data[2966] <= 8'h10 ;
			data[2967] <= 8'h10 ;
			data[2968] <= 8'h10 ;
			data[2969] <= 8'h10 ;
			data[2970] <= 8'h10 ;
			data[2971] <= 8'h10 ;
			data[2972] <= 8'h10 ;
			data[2973] <= 8'h10 ;
			data[2974] <= 8'h10 ;
			data[2975] <= 8'h10 ;
			data[2976] <= 8'h10 ;
			data[2977] <= 8'h10 ;
			data[2978] <= 8'h10 ;
			data[2979] <= 8'h10 ;
			data[2980] <= 8'h10 ;
			data[2981] <= 8'h10 ;
			data[2982] <= 8'h10 ;
			data[2983] <= 8'h10 ;
			data[2984] <= 8'h10 ;
			data[2985] <= 8'h10 ;
			data[2986] <= 8'h10 ;
			data[2987] <= 8'h10 ;
			data[2988] <= 8'h10 ;
			data[2989] <= 8'h10 ;
			data[2990] <= 8'h10 ;
			data[2991] <= 8'h10 ;
			data[2992] <= 8'h10 ;
			data[2993] <= 8'h10 ;
			data[2994] <= 8'h10 ;
			data[2995] <= 8'h10 ;
			data[2996] <= 8'h10 ;
			data[2997] <= 8'h10 ;
			data[2998] <= 8'h10 ;
			data[2999] <= 8'h10 ;
			data[3000] <= 8'h10 ;
			data[3001] <= 8'h10 ;
			data[3002] <= 8'h10 ;
			data[3003] <= 8'h10 ;
			data[3004] <= 8'h10 ;
			data[3005] <= 8'h10 ;
			data[3006] <= 8'h10 ;
			data[3007] <= 8'h10 ;
			data[3008] <= 8'h10 ;
			data[3009] <= 8'h10 ;
			data[3010] <= 8'h10 ;
			data[3011] <= 8'h10 ;
			data[3012] <= 8'h10 ;
			data[3013] <= 8'h10 ;
			data[3014] <= 8'h10 ;
			data[3015] <= 8'h10 ;
			data[3016] <= 8'h10 ;
			data[3017] <= 8'h10 ;
			data[3018] <= 8'h10 ;
			data[3019] <= 8'h10 ;
			data[3020] <= 8'h10 ;
			data[3021] <= 8'h10 ;
			data[3022] <= 8'h10 ;
			data[3023] <= 8'h10 ;
			data[3024] <= 8'h10 ;
			data[3025] <= 8'h10 ;
			data[3026] <= 8'h10 ;
			data[3027] <= 8'h10 ;
			data[3028] <= 8'h10 ;
			data[3029] <= 8'h10 ;
			data[3030] <= 8'h10 ;
			data[3031] <= 8'h10 ;
			data[3032] <= 8'h10 ;
			data[3033] <= 8'h10 ;
			data[3034] <= 8'h10 ;
			data[3035] <= 8'h10 ;
			data[3036] <= 8'h10 ;
			data[3037] <= 8'h10 ;
			data[3038] <= 8'h10 ;
			data[3039] <= 8'h10 ;
			data[3040] <= 8'h10 ;
			data[3041] <= 8'h10 ;
			data[3042] <= 8'h10 ;
			data[3043] <= 8'h10 ;
			data[3044] <= 8'h10 ;
			data[3045] <= 8'h10 ;
			data[3046] <= 8'h10 ;
			data[3047] <= 8'h10 ;
			data[3048] <= 8'h10 ;
			data[3049] <= 8'h10 ;
			data[3050] <= 8'h10 ;
			data[3051] <= 8'h10 ;
			data[3052] <= 8'h10 ;
			data[3053] <= 8'h10 ;
			data[3054] <= 8'h10 ;
			data[3055] <= 8'h10 ;
			data[3056] <= 8'h10 ;
			data[3057] <= 8'h10 ;
			data[3058] <= 8'h10 ;
			data[3059] <= 8'h10 ;
			data[3060] <= 8'h10 ;
			data[3061] <= 8'h10 ;
			data[3062] <= 8'h10 ;
			data[3063] <= 8'h10 ;
			data[3064] <= 8'h10 ;
			data[3065] <= 8'h10 ;
			data[3066] <= 8'h10 ;
			data[3067] <= 8'h10 ;
			data[3068] <= 8'h10 ;
			data[3069] <= 8'h10 ;
			data[3070] <= 8'h10 ;
			data[3071] <= 8'h10 ;
			data[3072] <= 8'h10 ;
			data[3073] <= 8'h10 ;
			data[3074] <= 8'h10 ;
			data[3075] <= 8'h10 ;
			data[3076] <= 8'h10 ;
			data[3077] <= 8'h10 ;
			data[3078] <= 8'h10 ;
			data[3079] <= 8'h10 ;
			data[3080] <= 8'h10 ;
			data[3081] <= 8'h10 ;
			data[3082] <= 8'h10 ;
			data[3083] <= 8'h10 ;
			data[3084] <= 8'h10 ;
			data[3085] <= 8'h10 ;
			data[3086] <= 8'h10 ;
			data[3087] <= 8'h10 ;
			data[3088] <= 8'h10 ;
			data[3089] <= 8'h10 ;
			data[3090] <= 8'h10 ;
			data[3091] <= 8'h10 ;
			data[3092] <= 8'h10 ;
			data[3093] <= 8'h10 ;
			data[3094] <= 8'h10 ;
			data[3095] <= 8'h10 ;
			data[3096] <= 8'h10 ;
			data[3097] <= 8'h10 ;
			data[3098] <= 8'h10 ;
			data[3099] <= 8'h10 ;
			data[3100] <= 8'h10 ;
			data[3101] <= 8'h10 ;
			data[3102] <= 8'h10 ;
			data[3103] <= 8'h10 ;
			data[3104] <= 8'h10 ;
			data[3105] <= 8'h10 ;
			data[3106] <= 8'h10 ;
			data[3107] <= 8'h10 ;
			data[3108] <= 8'h10 ;
			data[3109] <= 8'h10 ;
			data[3110] <= 8'h10 ;
			data[3111] <= 8'h10 ;
			data[3112] <= 8'h10 ;
			data[3113] <= 8'h10 ;
			data[3114] <= 8'h10 ;
			data[3115] <= 8'h10 ;
			data[3116] <= 8'h10 ;
			data[3117] <= 8'h10 ;
			data[3118] <= 8'h10 ;
			data[3119] <= 8'h10 ;
			data[3120] <= 8'h10 ;
			data[3121] <= 8'h10 ;
			data[3122] <= 8'h10 ;
			data[3123] <= 8'h10 ;
			data[3124] <= 8'h10 ;
			data[3125] <= 8'h10 ;
			data[3126] <= 8'h10 ;
			data[3127] <= 8'h10 ;
			data[3128] <= 8'h10 ;
			data[3129] <= 8'h10 ;
			data[3130] <= 8'h10 ;
			data[3131] <= 8'h10 ;
			data[3132] <= 8'h10 ;
			data[3133] <= 8'h10 ;
			data[3134] <= 8'h10 ;
			data[3135] <= 8'h10 ;
			data[3136] <= 8'h10 ;
			data[3137] <= 8'h10 ;
			data[3138] <= 8'h10 ;
			data[3139] <= 8'h10 ;
			data[3140] <= 8'h10 ;
			data[3141] <= 8'h10 ;
			data[3142] <= 8'h10 ;
			data[3143] <= 8'h10 ;
			data[3144] <= 8'h10 ;
			data[3145] <= 8'h10 ;
			data[3146] <= 8'h10 ;
			data[3147] <= 8'h10 ;
			data[3148] <= 8'h10 ;
			data[3149] <= 8'h10 ;
			data[3150] <= 8'h10 ;
			data[3151] <= 8'h10 ;
			data[3152] <= 8'h10 ;
			data[3153] <= 8'h10 ;
			data[3154] <= 8'h10 ;
			data[3155] <= 8'h10 ;
			data[3156] <= 8'h10 ;
			data[3157] <= 8'h10 ;
			data[3158] <= 8'h10 ;
			data[3159] <= 8'h10 ;
			data[3160] <= 8'h10 ;
			data[3161] <= 8'h10 ;
			data[3162] <= 8'h10 ;
			data[3163] <= 8'h10 ;
			data[3164] <= 8'h10 ;
			data[3165] <= 8'h10 ;
			data[3166] <= 8'h10 ;
			data[3167] <= 8'h10 ;
			data[3168] <= 8'h10 ;
			data[3169] <= 8'h10 ;
			data[3170] <= 8'h10 ;
			data[3171] <= 8'h10 ;
			data[3172] <= 8'h10 ;
			data[3173] <= 8'h10 ;
			data[3174] <= 8'h10 ;
			data[3175] <= 8'h10 ;
			data[3176] <= 8'h10 ;
			data[3177] <= 8'h10 ;
			data[3178] <= 8'h10 ;
			data[3179] <= 8'h10 ;
			data[3180] <= 8'h10 ;
			data[3181] <= 8'h10 ;
			data[3182] <= 8'h10 ;
			data[3183] <= 8'h10 ;
			data[3184] <= 8'h10 ;
			data[3185] <= 8'h10 ;
			data[3186] <= 8'h10 ;
			data[3187] <= 8'h10 ;
			data[3188] <= 8'h10 ;
			data[3189] <= 8'h10 ;
			data[3190] <= 8'h10 ;
			data[3191] <= 8'h10 ;
			data[3192] <= 8'h10 ;
			data[3193] <= 8'h10 ;
			data[3194] <= 8'h10 ;
			data[3195] <= 8'h10 ;
			data[3196] <= 8'h10 ;
			data[3197] <= 8'h10 ;
			data[3198] <= 8'h10 ;
			data[3199] <= 8'h10 ;
			data[3200] <= 8'h10 ;
			data[3201] <= 8'h10 ;
			data[3202] <= 8'h10 ;
			data[3203] <= 8'h10 ;
			data[3204] <= 8'h10 ;
			data[3205] <= 8'h10 ;
			data[3206] <= 8'h10 ;
			data[3207] <= 8'h10 ;
			data[3208] <= 8'h10 ;
			data[3209] <= 8'h10 ;
			data[3210] <= 8'h10 ;
			data[3211] <= 8'h10 ;
			data[3212] <= 8'h10 ;
			data[3213] <= 8'h10 ;
			data[3214] <= 8'h10 ;
			data[3215] <= 8'h10 ;
			data[3216] <= 8'h10 ;
			data[3217] <= 8'h10 ;
			data[3218] <= 8'h10 ;
			data[3219] <= 8'h10 ;
			data[3220] <= 8'h10 ;
			data[3221] <= 8'h10 ;
			data[3222] <= 8'h10 ;
			data[3223] <= 8'h10 ;
			data[3224] <= 8'h10 ;
			data[3225] <= 8'h10 ;
			data[3226] <= 8'h10 ;
			data[3227] <= 8'h10 ;
			data[3228] <= 8'h10 ;
			data[3229] <= 8'h10 ;
			data[3230] <= 8'h10 ;
			data[3231] <= 8'h10 ;
			data[3232] <= 8'h10 ;
			data[3233] <= 8'h10 ;
			data[3234] <= 8'h10 ;
			data[3235] <= 8'h10 ;
			data[3236] <= 8'h10 ;
			data[3237] <= 8'h10 ;
			data[3238] <= 8'h10 ;
			data[3239] <= 8'h10 ;
			data[3240] <= 8'h10 ;
			data[3241] <= 8'h10 ;
			data[3242] <= 8'h10 ;
			data[3243] <= 8'h10 ;
			data[3244] <= 8'h10 ;
			data[3245] <= 8'h10 ;
			data[3246] <= 8'h10 ;
			data[3247] <= 8'h10 ;
			data[3248] <= 8'h10 ;
			data[3249] <= 8'h10 ;
			data[3250] <= 8'h10 ;
			data[3251] <= 8'h10 ;
			data[3252] <= 8'h10 ;
			data[3253] <= 8'h10 ;
			data[3254] <= 8'h10 ;
			data[3255] <= 8'h10 ;
			data[3256] <= 8'h10 ;
			data[3257] <= 8'h10 ;
			data[3258] <= 8'h10 ;
			data[3259] <= 8'h10 ;
			data[3260] <= 8'h10 ;
			data[3261] <= 8'h10 ;
			data[3262] <= 8'h10 ;
			data[3263] <= 8'h10 ;
			data[3264] <= 8'h10 ;
			data[3265] <= 8'h10 ;
			data[3266] <= 8'h10 ;
			data[3267] <= 8'h10 ;
			data[3268] <= 8'h10 ;
			data[3269] <= 8'h10 ;
			data[3270] <= 8'h10 ;
			data[3271] <= 8'h10 ;
			data[3272] <= 8'h10 ;
			data[3273] <= 8'h10 ;
			data[3274] <= 8'h10 ;
			data[3275] <= 8'h10 ;
			data[3276] <= 8'h10 ;
			data[3277] <= 8'h10 ;
			data[3278] <= 8'h10 ;
			data[3279] <= 8'h10 ;
			data[3280] <= 8'h10 ;
			data[3281] <= 8'h10 ;
			data[3282] <= 8'h10 ;
			data[3283] <= 8'h10 ;
			data[3284] <= 8'h10 ;
			data[3285] <= 8'h10 ;
			data[3286] <= 8'h10 ;
			data[3287] <= 8'h10 ;
			data[3288] <= 8'h10 ;
			data[3289] <= 8'h10 ;
			data[3290] <= 8'h10 ;
			data[3291] <= 8'h10 ;
			data[3292] <= 8'h10 ;
			data[3293] <= 8'h10 ;
			data[3294] <= 8'h10 ;
			data[3295] <= 8'h10 ;
			data[3296] <= 8'h10 ;
			data[3297] <= 8'h10 ;
			data[3298] <= 8'h10 ;
			data[3299] <= 8'h10 ;
			data[3300] <= 8'h10 ;
			data[3301] <= 8'h10 ;
			data[3302] <= 8'h10 ;
			data[3303] <= 8'h10 ;
			data[3304] <= 8'h10 ;
			data[3305] <= 8'h10 ;
			data[3306] <= 8'h10 ;
			data[3307] <= 8'h10 ;
			data[3308] <= 8'h10 ;
			data[3309] <= 8'h10 ;
			data[3310] <= 8'h10 ;
			data[3311] <= 8'h10 ;
			data[3312] <= 8'h10 ;
			data[3313] <= 8'h10 ;
			data[3314] <= 8'h10 ;
			data[3315] <= 8'h10 ;
			data[3316] <= 8'h10 ;
			data[3317] <= 8'h10 ;
			data[3318] <= 8'h10 ;
			data[3319] <= 8'h10 ;
			data[3320] <= 8'h10 ;
			data[3321] <= 8'h10 ;
			data[3322] <= 8'h10 ;
			data[3323] <= 8'h10 ;
			data[3324] <= 8'h10 ;
			data[3325] <= 8'h10 ;
			data[3326] <= 8'h10 ;
			data[3327] <= 8'h10 ;
			data[3328] <= 8'h10 ;
			data[3329] <= 8'h10 ;
			data[3330] <= 8'h10 ;
			data[3331] <= 8'h10 ;
			data[3332] <= 8'h10 ;
			data[3333] <= 8'h10 ;
			data[3334] <= 8'h10 ;
			data[3335] <= 8'h10 ;
			data[3336] <= 8'h10 ;
			data[3337] <= 8'h10 ;
			data[3338] <= 8'h10 ;
			data[3339] <= 8'h10 ;
			data[3340] <= 8'h10 ;
			data[3341] <= 8'h10 ;
			data[3342] <= 8'h10 ;
			data[3343] <= 8'h10 ;
			data[3344] <= 8'h10 ;
			data[3345] <= 8'h10 ;
			data[3346] <= 8'h10 ;
			data[3347] <= 8'h10 ;
			data[3348] <= 8'h10 ;
			data[3349] <= 8'h10 ;
			data[3350] <= 8'h10 ;
			data[3351] <= 8'h10 ;
			data[3352] <= 8'h10 ;
			data[3353] <= 8'h10 ;
			data[3354] <= 8'h10 ;
			data[3355] <= 8'h10 ;
			data[3356] <= 8'h10 ;
			data[3357] <= 8'h10 ;
			data[3358] <= 8'h10 ;
			data[3359] <= 8'h10 ;
			data[3360] <= 8'h10 ;
			data[3361] <= 8'h10 ;
			data[3362] <= 8'h10 ;
			data[3363] <= 8'h10 ;
			data[3364] <= 8'h10 ;
			data[3365] <= 8'h10 ;
			data[3366] <= 8'h10 ;
			data[3367] <= 8'h10 ;
			data[3368] <= 8'h10 ;
			data[3369] <= 8'h10 ;
			data[3370] <= 8'h10 ;
			data[3371] <= 8'h10 ;
			data[3372] <= 8'h10 ;
			data[3373] <= 8'h10 ;
			data[3374] <= 8'h10 ;
			data[3375] <= 8'h10 ;
			data[3376] <= 8'h10 ;
			data[3377] <= 8'h10 ;
			data[3378] <= 8'h10 ;
			data[3379] <= 8'h10 ;
			data[3380] <= 8'h10 ;
			data[3381] <= 8'h10 ;
			data[3382] <= 8'h10 ;
			data[3383] <= 8'h10 ;
			data[3384] <= 8'h10 ;
			data[3385] <= 8'h10 ;
			data[3386] <= 8'h10 ;
			data[3387] <= 8'h10 ;
			data[3388] <= 8'h10 ;
			data[3389] <= 8'h10 ;
			data[3390] <= 8'h10 ;
			data[3391] <= 8'h10 ;
			data[3392] <= 8'h10 ;
			data[3393] <= 8'h10 ;
			data[3394] <= 8'h10 ;
			data[3395] <= 8'h10 ;
			data[3396] <= 8'h10 ;
			data[3397] <= 8'h10 ;
			data[3398] <= 8'h10 ;
			data[3399] <= 8'h10 ;
			data[3400] <= 8'h10 ;
			data[3401] <= 8'h10 ;
			data[3402] <= 8'h10 ;
			data[3403] <= 8'h10 ;
			data[3404] <= 8'h10 ;
			data[3405] <= 8'h10 ;
			data[3406] <= 8'h10 ;
			data[3407] <= 8'h10 ;
			data[3408] <= 8'h10 ;
			data[3409] <= 8'h10 ;
			data[3410] <= 8'h10 ;
			data[3411] <= 8'h10 ;
			data[3412] <= 8'h10 ;
			data[3413] <= 8'h10 ;
			data[3414] <= 8'h10 ;
			data[3415] <= 8'h10 ;
			data[3416] <= 8'h10 ;
			data[3417] <= 8'h10 ;
			data[3418] <= 8'h10 ;
			data[3419] <= 8'h10 ;
			data[3420] <= 8'h10 ;
			data[3421] <= 8'h10 ;
			data[3422] <= 8'h10 ;
			data[3423] <= 8'h10 ;
			data[3424] <= 8'h10 ;
			data[3425] <= 8'h10 ;
			data[3426] <= 8'h10 ;
			data[3427] <= 8'h10 ;
			data[3428] <= 8'h10 ;
			data[3429] <= 8'h10 ;
			data[3430] <= 8'h10 ;
			data[3431] <= 8'h10 ;
			data[3432] <= 8'h10 ;
			data[3433] <= 8'h10 ;
			data[3434] <= 8'h10 ;
			data[3435] <= 8'h10 ;
			data[3436] <= 8'h10 ;
			data[3437] <= 8'h10 ;
			data[3438] <= 8'h10 ;
			data[3439] <= 8'h10 ;
			data[3440] <= 8'h10 ;
			data[3441] <= 8'h10 ;
			data[3442] <= 8'h10 ;
			data[3443] <= 8'h10 ;
			data[3444] <= 8'h10 ;
			data[3445] <= 8'h10 ;
			data[3446] <= 8'h10 ;
			data[3447] <= 8'h10 ;
			data[3448] <= 8'h10 ;
			data[3449] <= 8'h10 ;
			data[3450] <= 8'h10 ;
			data[3451] <= 8'h10 ;
			data[3452] <= 8'h10 ;
			data[3453] <= 8'h10 ;
			data[3454] <= 8'h10 ;
			data[3455] <= 8'h10 ;
			data[3456] <= 8'h10 ;
			data[3457] <= 8'h10 ;
			data[3458] <= 8'h10 ;
			data[3459] <= 8'h10 ;
			data[3460] <= 8'h10 ;
			data[3461] <= 8'h10 ;
			data[3462] <= 8'h10 ;
			data[3463] <= 8'h10 ;
			data[3464] <= 8'h10 ;
			data[3465] <= 8'h10 ;
			data[3466] <= 8'h10 ;
			data[3467] <= 8'h10 ;
			data[3468] <= 8'h10 ;
			data[3469] <= 8'h10 ;
			data[3470] <= 8'h10 ;
			data[3471] <= 8'h10 ;
			data[3472] <= 8'h10 ;
			data[3473] <= 8'h10 ;
			data[3474] <= 8'h10 ;
			data[3475] <= 8'h10 ;
			data[3476] <= 8'h10 ;
			data[3477] <= 8'h10 ;
			data[3478] <= 8'h10 ;
			data[3479] <= 8'h10 ;
			data[3480] <= 8'h10 ;
			data[3481] <= 8'h10 ;
			data[3482] <= 8'h10 ;
			data[3483] <= 8'h10 ;
			data[3484] <= 8'h10 ;
			data[3485] <= 8'h10 ;
			data[3486] <= 8'h10 ;
			data[3487] <= 8'h10 ;
			data[3488] <= 8'h10 ;
			data[3489] <= 8'h10 ;
			data[3490] <= 8'h10 ;
			data[3491] <= 8'h10 ;
			data[3492] <= 8'h10 ;
			data[3493] <= 8'h10 ;
			data[3494] <= 8'h10 ;
			data[3495] <= 8'h10 ;
			data[3496] <= 8'h10 ;
			data[3497] <= 8'h10 ;
			data[3498] <= 8'h10 ;
			data[3499] <= 8'h10 ;
			data[3500] <= 8'h10 ;
			data[3501] <= 8'h10 ;
			data[3502] <= 8'h10 ;
			data[3503] <= 8'h10 ;
			data[3504] <= 8'h10 ;
			data[3505] <= 8'h10 ;
			data[3506] <= 8'h10 ;
			data[3507] <= 8'h10 ;
			data[3508] <= 8'h10 ;
			data[3509] <= 8'h10 ;
			data[3510] <= 8'h10 ;
			data[3511] <= 8'h10 ;
			data[3512] <= 8'h10 ;
			data[3513] <= 8'h10 ;
			data[3514] <= 8'h10 ;
			data[3515] <= 8'h10 ;
			data[3516] <= 8'h10 ;
			data[3517] <= 8'h10 ;
			data[3518] <= 8'h10 ;
			data[3519] <= 8'h10 ;
			data[3520] <= 8'h10 ;
			data[3521] <= 8'h10 ;
			data[3522] <= 8'h10 ;
			data[3523] <= 8'h10 ;
			data[3524] <= 8'h10 ;
			data[3525] <= 8'h10 ;
			data[3526] <= 8'h10 ;
			data[3527] <= 8'h10 ;
			data[3528] <= 8'h10 ;
			data[3529] <= 8'h10 ;
			data[3530] <= 8'h10 ;
			data[3531] <= 8'h10 ;
			data[3532] <= 8'h10 ;
			data[3533] <= 8'h10 ;
			data[3534] <= 8'h10 ;
			data[3535] <= 8'h10 ;
			data[3536] <= 8'h10 ;
			data[3537] <= 8'h10 ;
			data[3538] <= 8'h10 ;
			data[3539] <= 8'h10 ;
			data[3540] <= 8'h10 ;
			data[3541] <= 8'h10 ;
			data[3542] <= 8'h10 ;
			data[3543] <= 8'h10 ;
			data[3544] <= 8'h10 ;
			data[3545] <= 8'h10 ;
			data[3546] <= 8'h10 ;
			data[3547] <= 8'h10 ;
			data[3548] <= 8'h10 ;
			data[3549] <= 8'h10 ;
			data[3550] <= 8'h10 ;
			data[3551] <= 8'h10 ;
			data[3552] <= 8'h10 ;
			data[3553] <= 8'h10 ;
			data[3554] <= 8'h10 ;
			data[3555] <= 8'h10 ;
			data[3556] <= 8'h10 ;
			data[3557] <= 8'h10 ;
			data[3558] <= 8'h10 ;
			data[3559] <= 8'h10 ;
			data[3560] <= 8'h10 ;
			data[3561] <= 8'h10 ;
			data[3562] <= 8'h10 ;
			data[3563] <= 8'h10 ;
			data[3564] <= 8'h10 ;
			data[3565] <= 8'h10 ;
			data[3566] <= 8'h10 ;
			data[3567] <= 8'h10 ;
			data[3568] <= 8'h10 ;
			data[3569] <= 8'h10 ;
			data[3570] <= 8'h10 ;
			data[3571] <= 8'h10 ;
			data[3572] <= 8'h10 ;
			data[3573] <= 8'h10 ;
			data[3574] <= 8'h10 ;
			data[3575] <= 8'h10 ;
			data[3576] <= 8'h10 ;
			data[3577] <= 8'h10 ;
			data[3578] <= 8'h10 ;
			data[3579] <= 8'h10 ;
			data[3580] <= 8'h10 ;
			data[3581] <= 8'h10 ;
			data[3582] <= 8'h10 ;
			data[3583] <= 8'h10 ;
			data[3584] <= 8'h10 ;
			data[3585] <= 8'h10 ;
			data[3586] <= 8'h10 ;
			data[3587] <= 8'h10 ;
			data[3588] <= 8'h10 ;
			data[3589] <= 8'h10 ;
			data[3590] <= 8'h10 ;
			data[3591] <= 8'h10 ;
			data[3592] <= 8'h10 ;
			data[3593] <= 8'h10 ;
			data[3594] <= 8'h10 ;
			data[3595] <= 8'h10 ;
			data[3596] <= 8'h10 ;
			data[3597] <= 8'h10 ;
			data[3598] <= 8'h10 ;
			data[3599] <= 8'h10 ;
			data[3600] <= 8'h10 ;
			data[3601] <= 8'h10 ;
			data[3602] <= 8'h10 ;
			data[3603] <= 8'h10 ;
			data[3604] <= 8'h10 ;
			data[3605] <= 8'h10 ;
			data[3606] <= 8'h10 ;
			data[3607] <= 8'h10 ;
			data[3608] <= 8'h10 ;
			data[3609] <= 8'h10 ;
			data[3610] <= 8'h10 ;
			data[3611] <= 8'h10 ;
			data[3612] <= 8'h10 ;
			data[3613] <= 8'h10 ;
			data[3614] <= 8'h10 ;
			data[3615] <= 8'h10 ;
			data[3616] <= 8'h10 ;
			data[3617] <= 8'h10 ;
			data[3618] <= 8'h10 ;
			data[3619] <= 8'h10 ;
			data[3620] <= 8'h10 ;
			data[3621] <= 8'h10 ;
			data[3622] <= 8'h10 ;
			data[3623] <= 8'h10 ;
			data[3624] <= 8'h10 ;
			data[3625] <= 8'h10 ;
			data[3626] <= 8'h10 ;
			data[3627] <= 8'h10 ;
			data[3628] <= 8'h10 ;
			data[3629] <= 8'h10 ;
			data[3630] <= 8'h10 ;
			data[3631] <= 8'h10 ;
			data[3632] <= 8'h10 ;
			data[3633] <= 8'h10 ;
			data[3634] <= 8'h10 ;
			data[3635] <= 8'h10 ;
			data[3636] <= 8'h10 ;
			data[3637] <= 8'h10 ;
			data[3638] <= 8'h10 ;
			data[3639] <= 8'h10 ;
			data[3640] <= 8'h10 ;
			data[3641] <= 8'h10 ;
			data[3642] <= 8'h10 ;
			data[3643] <= 8'h10 ;
			data[3644] <= 8'h10 ;
			data[3645] <= 8'h10 ;
			data[3646] <= 8'h10 ;
			data[3647] <= 8'h10 ;
			data[3648] <= 8'h10 ;
			data[3649] <= 8'h10 ;
			data[3650] <= 8'h10 ;
			data[3651] <= 8'h10 ;
			data[3652] <= 8'h10 ;
			data[3653] <= 8'h10 ;
			data[3654] <= 8'h10 ;
			data[3655] <= 8'h10 ;
			data[3656] <= 8'h10 ;
			data[3657] <= 8'h10 ;
			data[3658] <= 8'h10 ;
			data[3659] <= 8'h10 ;
			data[3660] <= 8'h10 ;
			data[3661] <= 8'h10 ;
			data[3662] <= 8'h10 ;
			data[3663] <= 8'h10 ;
			data[3664] <= 8'h10 ;
			data[3665] <= 8'h10 ;
			data[3666] <= 8'h10 ;
			data[3667] <= 8'h10 ;
			data[3668] <= 8'h10 ;
			data[3669] <= 8'h10 ;
			data[3670] <= 8'h10 ;
			data[3671] <= 8'h10 ;
			data[3672] <= 8'h10 ;
			data[3673] <= 8'h10 ;
			data[3674] <= 8'h10 ;
			data[3675] <= 8'h10 ;
			data[3676] <= 8'h10 ;
			data[3677] <= 8'h10 ;
			data[3678] <= 8'h10 ;
			data[3679] <= 8'h10 ;
			data[3680] <= 8'h10 ;
			data[3681] <= 8'h10 ;
			data[3682] <= 8'h10 ;
			data[3683] <= 8'h10 ;
			data[3684] <= 8'h10 ;
			data[3685] <= 8'h10 ;
			data[3686] <= 8'h10 ;
			data[3687] <= 8'h10 ;
			data[3688] <= 8'h10 ;
			data[3689] <= 8'h10 ;
			data[3690] <= 8'h10 ;
			data[3691] <= 8'h10 ;
			data[3692] <= 8'h10 ;
			data[3693] <= 8'h10 ;
			data[3694] <= 8'h10 ;
			data[3695] <= 8'h10 ;
			data[3696] <= 8'h10 ;
			data[3697] <= 8'h10 ;
			data[3698] <= 8'h10 ;
			data[3699] <= 8'h10 ;
			data[3700] <= 8'h10 ;
			data[3701] <= 8'h10 ;
			data[3702] <= 8'h10 ;
			data[3703] <= 8'h10 ;
			data[3704] <= 8'h10 ;
			data[3705] <= 8'h10 ;
			data[3706] <= 8'h10 ;
			data[3707] <= 8'h10 ;
			data[3708] <= 8'h10 ;
			data[3709] <= 8'h10 ;
			data[3710] <= 8'h10 ;
			data[3711] <= 8'h10 ;
			data[3712] <= 8'h10 ;
			data[3713] <= 8'h10 ;
			data[3714] <= 8'h10 ;
			data[3715] <= 8'h10 ;
			data[3716] <= 8'h10 ;
			data[3717] <= 8'h10 ;
			data[3718] <= 8'h10 ;
			data[3719] <= 8'h10 ;
			data[3720] <= 8'h10 ;
			data[3721] <= 8'h10 ;
			data[3722] <= 8'h10 ;
			data[3723] <= 8'h10 ;
			data[3724] <= 8'h10 ;
			data[3725] <= 8'h10 ;
			data[3726] <= 8'h10 ;
			data[3727] <= 8'h10 ;
			data[3728] <= 8'h10 ;
			data[3729] <= 8'h10 ;
			data[3730] <= 8'h10 ;
			data[3731] <= 8'h10 ;
			data[3732] <= 8'h10 ;
			data[3733] <= 8'h10 ;
			data[3734] <= 8'h10 ;
			data[3735] <= 8'h10 ;
			data[3736] <= 8'h10 ;
			data[3737] <= 8'h10 ;
			data[3738] <= 8'h10 ;
			data[3739] <= 8'h10 ;
			data[3740] <= 8'h10 ;
			data[3741] <= 8'h10 ;
			data[3742] <= 8'h10 ;
			data[3743] <= 8'h10 ;
			data[3744] <= 8'h10 ;
			data[3745] <= 8'h10 ;
			data[3746] <= 8'h10 ;
			data[3747] <= 8'h10 ;
			data[3748] <= 8'h10 ;
			data[3749] <= 8'h10 ;
			data[3750] <= 8'h10 ;
			data[3751] <= 8'h10 ;
			data[3752] <= 8'h10 ;
			data[3753] <= 8'h10 ;
			data[3754] <= 8'h10 ;
			data[3755] <= 8'h10 ;
			data[3756] <= 8'h10 ;
			data[3757] <= 8'h10 ;
			data[3758] <= 8'h10 ;
			data[3759] <= 8'h10 ;
			data[3760] <= 8'h10 ;
			data[3761] <= 8'h10 ;
			data[3762] <= 8'h10 ;
			data[3763] <= 8'h10 ;
			data[3764] <= 8'h10 ;
			data[3765] <= 8'h10 ;
			data[3766] <= 8'h10 ;
			data[3767] <= 8'h10 ;
			data[3768] <= 8'h10 ;
			data[3769] <= 8'h10 ;
			data[3770] <= 8'h10 ;
			data[3771] <= 8'h10 ;
			data[3772] <= 8'h10 ;
			data[3773] <= 8'h10 ;
			data[3774] <= 8'h10 ;
			data[3775] <= 8'h10 ;
			data[3776] <= 8'h10 ;
			data[3777] <= 8'h10 ;
			data[3778] <= 8'h10 ;
			data[3779] <= 8'h10 ;
			data[3780] <= 8'h10 ;
			data[3781] <= 8'h10 ;
			data[3782] <= 8'h10 ;
			data[3783] <= 8'h10 ;
			data[3784] <= 8'h10 ;
			data[3785] <= 8'h10 ;
			data[3786] <= 8'h10 ;
			data[3787] <= 8'h10 ;
			data[3788] <= 8'h10 ;
			data[3789] <= 8'h10 ;
			data[3790] <= 8'h10 ;
			data[3791] <= 8'h10 ;
			data[3792] <= 8'h10 ;
			data[3793] <= 8'h10 ;
			data[3794] <= 8'h10 ;
			data[3795] <= 8'h10 ;
			data[3796] <= 8'h10 ;
			data[3797] <= 8'h10 ;
			data[3798] <= 8'h10 ;
			data[3799] <= 8'h10 ;
			data[3800] <= 8'h10 ;
			data[3801] <= 8'h10 ;
			data[3802] <= 8'h10 ;
			data[3803] <= 8'h10 ;
			data[3804] <= 8'h10 ;
			data[3805] <= 8'h10 ;
			data[3806] <= 8'h10 ;
			data[3807] <= 8'h10 ;
			data[3808] <= 8'h10 ;
			data[3809] <= 8'h10 ;
			data[3810] <= 8'h10 ;
			data[3811] <= 8'h10 ;
			data[3812] <= 8'h10 ;
			data[3813] <= 8'h10 ;
			data[3814] <= 8'h10 ;
			data[3815] <= 8'h10 ;
			data[3816] <= 8'h10 ;
			data[3817] <= 8'h10 ;
			data[3818] <= 8'h10 ;
			data[3819] <= 8'h10 ;
			data[3820] <= 8'h10 ;
			data[3821] <= 8'h10 ;
			data[3822] <= 8'h10 ;
			data[3823] <= 8'h10 ;
			data[3824] <= 8'h10 ;
			data[3825] <= 8'h10 ;
			data[3826] <= 8'h10 ;
			data[3827] <= 8'h10 ;
			data[3828] <= 8'h10 ;
			data[3829] <= 8'h10 ;
			data[3830] <= 8'h10 ;
			data[3831] <= 8'h10 ;
			data[3832] <= 8'h10 ;
			data[3833] <= 8'h10 ;
			data[3834] <= 8'h10 ;
			data[3835] <= 8'h10 ;
			data[3836] <= 8'h10 ;
			data[3837] <= 8'h10 ;
			data[3838] <= 8'h10 ;
			data[3839] <= 8'h10 ;
			data[3840] <= 8'h10 ;
			data[3841] <= 8'h10 ;
			data[3842] <= 8'h10 ;
			data[3843] <= 8'h10 ;
			data[3844] <= 8'h10 ;
			data[3845] <= 8'h10 ;
			data[3846] <= 8'h10 ;
			data[3847] <= 8'h10 ;
			data[3848] <= 8'h10 ;
			data[3849] <= 8'h10 ;
			data[3850] <= 8'h10 ;
			data[3851] <= 8'h10 ;
			data[3852] <= 8'h10 ;
			data[3853] <= 8'h10 ;
			data[3854] <= 8'h10 ;
			data[3855] <= 8'h10 ;
			data[3856] <= 8'h10 ;
			data[3857] <= 8'h10 ;
			data[3858] <= 8'h10 ;
			data[3859] <= 8'h10 ;
			data[3860] <= 8'h10 ;
			data[3861] <= 8'h10 ;
			data[3862] <= 8'h10 ;
			data[3863] <= 8'h10 ;
			data[3864] <= 8'h10 ;
			data[3865] <= 8'h10 ;
			data[3866] <= 8'h10 ;
			data[3867] <= 8'h10 ;
			data[3868] <= 8'h10 ;
			data[3869] <= 8'h10 ;
			data[3870] <= 8'h10 ;
			data[3871] <= 8'h10 ;
			data[3872] <= 8'h10 ;
			data[3873] <= 8'h10 ;
			data[3874] <= 8'h10 ;
			data[3875] <= 8'h10 ;
			data[3876] <= 8'h10 ;
			data[3877] <= 8'h10 ;
			data[3878] <= 8'h10 ;
			data[3879] <= 8'h10 ;
			data[3880] <= 8'h10 ;
			data[3881] <= 8'h10 ;
			data[3882] <= 8'h10 ;
			data[3883] <= 8'h10 ;
			data[3884] <= 8'h10 ;
			data[3885] <= 8'h10 ;
			data[3886] <= 8'h10 ;
			data[3887] <= 8'h10 ;
			data[3888] <= 8'h10 ;
			data[3889] <= 8'h10 ;
			data[3890] <= 8'h10 ;
			data[3891] <= 8'h10 ;
			data[3892] <= 8'h10 ;
			data[3893] <= 8'h10 ;
			data[3894] <= 8'h10 ;
			data[3895] <= 8'h10 ;
			data[3896] <= 8'h10 ;
			data[3897] <= 8'h10 ;
			data[3898] <= 8'h10 ;
			data[3899] <= 8'h10 ;
			data[3900] <= 8'h10 ;
			data[3901] <= 8'h10 ;
			data[3902] <= 8'h10 ;
			data[3903] <= 8'h10 ;
			data[3904] <= 8'h10 ;
			data[3905] <= 8'h10 ;
			data[3906] <= 8'h10 ;
			data[3907] <= 8'h10 ;
			data[3908] <= 8'h10 ;
			data[3909] <= 8'h10 ;
			data[3910] <= 8'h10 ;
			data[3911] <= 8'h10 ;
			data[3912] <= 8'h10 ;
			data[3913] <= 8'h10 ;
			data[3914] <= 8'h10 ;
			data[3915] <= 8'h10 ;
			data[3916] <= 8'h10 ;
			data[3917] <= 8'h10 ;
			data[3918] <= 8'h10 ;
			data[3919] <= 8'h10 ;
			data[3920] <= 8'h10 ;
			data[3921] <= 8'h10 ;
			data[3922] <= 8'h10 ;
			data[3923] <= 8'h10 ;
			data[3924] <= 8'h10 ;
			data[3925] <= 8'h10 ;
			data[3926] <= 8'h10 ;
			data[3927] <= 8'h10 ;
			data[3928] <= 8'h10 ;
			data[3929] <= 8'h10 ;
			data[3930] <= 8'h10 ;
			data[3931] <= 8'h10 ;
			data[3932] <= 8'h10 ;
			data[3933] <= 8'h10 ;
			data[3934] <= 8'h10 ;
			data[3935] <= 8'h10 ;
			data[3936] <= 8'h10 ;
			data[3937] <= 8'h10 ;
			data[3938] <= 8'h10 ;
			data[3939] <= 8'h10 ;
			data[3940] <= 8'h10 ;
			data[3941] <= 8'h10 ;
			data[3942] <= 8'h10 ;
			data[3943] <= 8'h10 ;
			data[3944] <= 8'h10 ;
			data[3945] <= 8'h10 ;
			data[3946] <= 8'h10 ;
			data[3947] <= 8'h10 ;
			data[3948] <= 8'h10 ;
			data[3949] <= 8'h10 ;
			data[3950] <= 8'h10 ;
			data[3951] <= 8'h10 ;
			data[3952] <= 8'h10 ;
			data[3953] <= 8'h10 ;
			data[3954] <= 8'h10 ;
			data[3955] <= 8'h10 ;
			data[3956] <= 8'h10 ;
			data[3957] <= 8'h10 ;
			data[3958] <= 8'h10 ;
			data[3959] <= 8'h10 ;
			data[3960] <= 8'h10 ;
			data[3961] <= 8'h10 ;
			data[3962] <= 8'h10 ;
			data[3963] <= 8'h10 ;
			data[3964] <= 8'h10 ;
			data[3965] <= 8'h10 ;
			data[3966] <= 8'h10 ;
			data[3967] <= 8'h10 ;
			data[3968] <= 8'h10 ;
			data[3969] <= 8'h10 ;
			data[3970] <= 8'h10 ;
			data[3971] <= 8'h10 ;
			data[3972] <= 8'h10 ;
			data[3973] <= 8'h10 ;
			data[3974] <= 8'h10 ;
			data[3975] <= 8'h10 ;
			data[3976] <= 8'h10 ;
			data[3977] <= 8'h10 ;
			data[3978] <= 8'h10 ;
			data[3979] <= 8'h10 ;
			data[3980] <= 8'h10 ;
			data[3981] <= 8'h10 ;
			data[3982] <= 8'h10 ;
			data[3983] <= 8'h10 ;
			data[3984] <= 8'h10 ;
			data[3985] <= 8'h10 ;
			data[3986] <= 8'h10 ;
			data[3987] <= 8'h10 ;
			data[3988] <= 8'h10 ;
			data[3989] <= 8'h10 ;
			data[3990] <= 8'h10 ;
			data[3991] <= 8'h10 ;
			data[3992] <= 8'h10 ;
			data[3993] <= 8'h10 ;
			data[3994] <= 8'h10 ;
			data[3995] <= 8'h10 ;
			data[3996] <= 8'h10 ;
			data[3997] <= 8'h10 ;
			data[3998] <= 8'h10 ;
			data[3999] <= 8'h10 ;
			data[4000] <= 8'h10 ;
			data[4001] <= 8'h10 ;
			data[4002] <= 8'h10 ;
			data[4003] <= 8'h10 ;
			data[4004] <= 8'h10 ;
			data[4005] <= 8'h10 ;
			data[4006] <= 8'h10 ;
			data[4007] <= 8'h10 ;
			data[4008] <= 8'h10 ;
			data[4009] <= 8'h10 ;
			data[4010] <= 8'h10 ;
			data[4011] <= 8'h10 ;
			data[4012] <= 8'h10 ;
			data[4013] <= 8'h10 ;
			data[4014] <= 8'h10 ;
			data[4015] <= 8'h10 ;
			data[4016] <= 8'h10 ;
			data[4017] <= 8'h10 ;
			data[4018] <= 8'h10 ;
			data[4019] <= 8'h10 ;
			data[4020] <= 8'h10 ;
			data[4021] <= 8'h10 ;
			data[4022] <= 8'h10 ;
			data[4023] <= 8'h10 ;
			data[4024] <= 8'h10 ;
			data[4025] <= 8'h10 ;
			data[4026] <= 8'h10 ;
			data[4027] <= 8'h10 ;
			data[4028] <= 8'h10 ;
			data[4029] <= 8'h10 ;
			data[4030] <= 8'h10 ;
			data[4031] <= 8'h10 ;
			data[4032] <= 8'h10 ;
			data[4033] <= 8'h10 ;
			data[4034] <= 8'h10 ;
			data[4035] <= 8'h10 ;
			data[4036] <= 8'h10 ;
			data[4037] <= 8'h10 ;
			data[4038] <= 8'h10 ;
			data[4039] <= 8'h10 ;
			data[4040] <= 8'h10 ;
			data[4041] <= 8'h10 ;
			data[4042] <= 8'h10 ;
			data[4043] <= 8'h10 ;
			data[4044] <= 8'h10 ;
			data[4045] <= 8'h10 ;
			data[4046] <= 8'h10 ;
			data[4047] <= 8'h10 ;
			data[4048] <= 8'h10 ;
			data[4049] <= 8'h10 ;
			data[4050] <= 8'h10 ;
			data[4051] <= 8'h10 ;
			data[4052] <= 8'h10 ;
			data[4053] <= 8'h10 ;
			data[4054] <= 8'h10 ;
			data[4055] <= 8'h10 ;
			data[4056] <= 8'h10 ;
			data[4057] <= 8'h10 ;
			data[4058] <= 8'h10 ;
			data[4059] <= 8'h10 ;
			data[4060] <= 8'h10 ;
			data[4061] <= 8'h10 ;
			data[4062] <= 8'h10 ;
			data[4063] <= 8'h10 ;
			data[4064] <= 8'h10 ;
			data[4065] <= 8'h10 ;
			data[4066] <= 8'h10 ;
			data[4067] <= 8'h10 ;
			data[4068] <= 8'h10 ;
			data[4069] <= 8'h10 ;
			data[4070] <= 8'h10 ;
			data[4071] <= 8'h10 ;
			data[4072] <= 8'h10 ;
			data[4073] <= 8'h10 ;
			data[4074] <= 8'h10 ;
			data[4075] <= 8'h10 ;
			data[4076] <= 8'h10 ;
			data[4077] <= 8'h10 ;
			data[4078] <= 8'h10 ;
			data[4079] <= 8'h10 ;
			data[4080] <= 8'h10 ;
			data[4081] <= 8'h10 ;
			data[4082] <= 8'h10 ;
			data[4083] <= 8'h10 ;
			data[4084] <= 8'h10 ;
			data[4085] <= 8'h10 ;
			data[4086] <= 8'h10 ;
			data[4087] <= 8'h10 ;
			data[4088] <= 8'h10 ;
			data[4089] <= 8'h10 ;
			data[4090] <= 8'h10 ;
			data[4091] <= 8'h10 ;
			data[4092] <= 8'h10 ;
			data[4093] <= 8'h10 ;
			data[4094] <= 8'h10 ;
			data[4095] <= 8'h10 ;
			data[4096] <= 8'h10 ;
			data[4097] <= 8'h10 ;
			data[4098] <= 8'h10 ;
			data[4099] <= 8'h10 ;
			data[4100] <= 8'h10 ;
			data[4101] <= 8'h10 ;
			data[4102] <= 8'h10 ;
			data[4103] <= 8'h10 ;
			data[4104] <= 8'h10 ;
			data[4105] <= 8'h10 ;
			data[4106] <= 8'h10 ;
			data[4107] <= 8'h10 ;
			data[4108] <= 8'h10 ;
			data[4109] <= 8'h10 ;
			data[4110] <= 8'h10 ;
			data[4111] <= 8'h10 ;
			data[4112] <= 8'h10 ;
			data[4113] <= 8'h10 ;
			data[4114] <= 8'h10 ;
			data[4115] <= 8'h10 ;
			data[4116] <= 8'h10 ;
			data[4117] <= 8'h10 ;
			data[4118] <= 8'h10 ;
			data[4119] <= 8'h10 ;
			data[4120] <= 8'h10 ;
			data[4121] <= 8'h10 ;
			data[4122] <= 8'h10 ;
			data[4123] <= 8'h10 ;
			data[4124] <= 8'h10 ;
			data[4125] <= 8'h10 ;
			data[4126] <= 8'h10 ;
			data[4127] <= 8'h10 ;
			data[4128] <= 8'h10 ;
			data[4129] <= 8'h10 ;
			data[4130] <= 8'h10 ;
			data[4131] <= 8'h10 ;
			data[4132] <= 8'h10 ;
			data[4133] <= 8'h10 ;
			data[4134] <= 8'h10 ;
			data[4135] <= 8'h10 ;
			data[4136] <= 8'h10 ;
			data[4137] <= 8'h10 ;
			data[4138] <= 8'h10 ;
			data[4139] <= 8'h10 ;
			data[4140] <= 8'h10 ;
			data[4141] <= 8'h10 ;
			data[4142] <= 8'h10 ;
			data[4143] <= 8'h10 ;
			data[4144] <= 8'h10 ;
			data[4145] <= 8'h10 ;
			data[4146] <= 8'h10 ;
			data[4147] <= 8'h10 ;
			data[4148] <= 8'h10 ;
			data[4149] <= 8'h10 ;
			data[4150] <= 8'h10 ;
			data[4151] <= 8'h10 ;
			data[4152] <= 8'h10 ;
			data[4153] <= 8'h10 ;
			data[4154] <= 8'h10 ;
			data[4155] <= 8'h10 ;
			data[4156] <= 8'h10 ;
			data[4157] <= 8'h10 ;
			data[4158] <= 8'h10 ;
			data[4159] <= 8'h10 ;
			data[4160] <= 8'h10 ;
			data[4161] <= 8'h10 ;
			data[4162] <= 8'h10 ;
			data[4163] <= 8'h10 ;
			data[4164] <= 8'h10 ;
			data[4165] <= 8'h10 ;
			data[4166] <= 8'h10 ;
			data[4167] <= 8'h10 ;
			data[4168] <= 8'h10 ;
			data[4169] <= 8'h10 ;
			data[4170] <= 8'h10 ;
			data[4171] <= 8'h10 ;
			data[4172] <= 8'h10 ;
			data[4173] <= 8'h10 ;
			data[4174] <= 8'h10 ;
			data[4175] <= 8'h10 ;
			data[4176] <= 8'h10 ;
			data[4177] <= 8'h10 ;
			data[4178] <= 8'h10 ;
			data[4179] <= 8'h10 ;
			data[4180] <= 8'h10 ;
			data[4181] <= 8'h10 ;
			data[4182] <= 8'h10 ;
			data[4183] <= 8'h10 ;
			data[4184] <= 8'h10 ;
			data[4185] <= 8'h10 ;
			data[4186] <= 8'h10 ;
			data[4187] <= 8'h10 ;
			data[4188] <= 8'h10 ;
			data[4189] <= 8'h10 ;
			data[4190] <= 8'h10 ;
			data[4191] <= 8'h10 ;
			data[4192] <= 8'h10 ;
			data[4193] <= 8'h10 ;
			data[4194] <= 8'h10 ;
			data[4195] <= 8'h10 ;
			data[4196] <= 8'h10 ;
			data[4197] <= 8'h10 ;
			data[4198] <= 8'h10 ;
			data[4199] <= 8'h10 ;
			data[4200] <= 8'h10 ;
			data[4201] <= 8'h10 ;
			data[4202] <= 8'h10 ;
			data[4203] <= 8'h10 ;
			data[4204] <= 8'h10 ;
			data[4205] <= 8'h10 ;
			data[4206] <= 8'h10 ;
			data[4207] <= 8'h10 ;
			data[4208] <= 8'h10 ;
			data[4209] <= 8'h10 ;
			data[4210] <= 8'h10 ;
			data[4211] <= 8'h10 ;
			data[4212] <= 8'h10 ;
			data[4213] <= 8'h10 ;
			data[4214] <= 8'h10 ;
			data[4215] <= 8'h10 ;
			data[4216] <= 8'h10 ;
			data[4217] <= 8'h10 ;
			data[4218] <= 8'h10 ;
			data[4219] <= 8'h10 ;
			data[4220] <= 8'h10 ;
			data[4221] <= 8'h10 ;
			data[4222] <= 8'h10 ;
			data[4223] <= 8'h10 ;
			data[4224] <= 8'h10 ;
			data[4225] <= 8'h10 ;
			data[4226] <= 8'h10 ;
			data[4227] <= 8'h10 ;
			data[4228] <= 8'h10 ;
			data[4229] <= 8'h10 ;
			data[4230] <= 8'h10 ;
			data[4231] <= 8'h10 ;
			data[4232] <= 8'h10 ;
			data[4233] <= 8'h10 ;
			data[4234] <= 8'h10 ;
			data[4235] <= 8'h10 ;
			data[4236] <= 8'h10 ;
			data[4237] <= 8'h10 ;
			data[4238] <= 8'h10 ;
			data[4239] <= 8'h10 ;
			data[4240] <= 8'h10 ;
			data[4241] <= 8'h10 ;
			data[4242] <= 8'h10 ;
			data[4243] <= 8'h10 ;
			data[4244] <= 8'h10 ;
			data[4245] <= 8'h10 ;
			data[4246] <= 8'h10 ;
			data[4247] <= 8'h10 ;
			data[4248] <= 8'h10 ;
			data[4249] <= 8'h10 ;
			data[4250] <= 8'h10 ;
			data[4251] <= 8'h10 ;
			data[4252] <= 8'h10 ;
			data[4253] <= 8'h10 ;
			data[4254] <= 8'h10 ;
			data[4255] <= 8'h10 ;
			data[4256] <= 8'h10 ;
			data[4257] <= 8'h10 ;
			data[4258] <= 8'h10 ;
			data[4259] <= 8'h10 ;
			data[4260] <= 8'h10 ;
			data[4261] <= 8'h10 ;
			data[4262] <= 8'h10 ;
			data[4263] <= 8'h10 ;
			data[4264] <= 8'h10 ;
			data[4265] <= 8'h10 ;
			data[4266] <= 8'h10 ;
			data[4267] <= 8'h10 ;
			data[4268] <= 8'h10 ;
			data[4269] <= 8'h10 ;
			data[4270] <= 8'h10 ;
			data[4271] <= 8'h10 ;
			data[4272] <= 8'h10 ;
			data[4273] <= 8'h10 ;
			data[4274] <= 8'h10 ;
			data[4275] <= 8'h10 ;
			data[4276] <= 8'h10 ;
			data[4277] <= 8'h10 ;
			data[4278] <= 8'h10 ;
			data[4279] <= 8'h10 ;
			data[4280] <= 8'h10 ;
			data[4281] <= 8'h10 ;
			data[4282] <= 8'h10 ;
			data[4283] <= 8'h10 ;
			data[4284] <= 8'h10 ;
			data[4285] <= 8'h10 ;
			data[4286] <= 8'h10 ;
			data[4287] <= 8'h10 ;
			data[4288] <= 8'h10 ;
			data[4289] <= 8'h10 ;
			data[4290] <= 8'h10 ;
			data[4291] <= 8'h10 ;
			data[4292] <= 8'h10 ;
			data[4293] <= 8'h10 ;
			data[4294] <= 8'h10 ;
			data[4295] <= 8'h10 ;
			data[4296] <= 8'h10 ;
			data[4297] <= 8'h10 ;
			data[4298] <= 8'h10 ;
			data[4299] <= 8'h10 ;
			data[4300] <= 8'h10 ;
			data[4301] <= 8'h10 ;
			data[4302] <= 8'h10 ;
			data[4303] <= 8'h10 ;
			data[4304] <= 8'h10 ;
			data[4305] <= 8'h10 ;
			data[4306] <= 8'h10 ;
			data[4307] <= 8'h10 ;
			data[4308] <= 8'h10 ;
			data[4309] <= 8'h10 ;
			data[4310] <= 8'h10 ;
			data[4311] <= 8'h10 ;
			data[4312] <= 8'h10 ;
			data[4313] <= 8'h10 ;
			data[4314] <= 8'h10 ;
			data[4315] <= 8'h10 ;
			data[4316] <= 8'h10 ;
			data[4317] <= 8'h10 ;
			data[4318] <= 8'h10 ;
			data[4319] <= 8'h10 ;
			data[4320] <= 8'h10 ;
			data[4321] <= 8'h10 ;
			data[4322] <= 8'h10 ;
			data[4323] <= 8'h10 ;
			data[4324] <= 8'h10 ;
			data[4325] <= 8'h10 ;
			data[4326] <= 8'h10 ;
			data[4327] <= 8'h10 ;
			data[4328] <= 8'h10 ;
			data[4329] <= 8'h10 ;
			data[4330] <= 8'h10 ;
			data[4331] <= 8'h10 ;
			data[4332] <= 8'h10 ;
			data[4333] <= 8'h10 ;
			data[4334] <= 8'h10 ;
			data[4335] <= 8'h10 ;
			data[4336] <= 8'h10 ;
			data[4337] <= 8'h10 ;
			data[4338] <= 8'h10 ;
			data[4339] <= 8'h10 ;
			data[4340] <= 8'h10 ;
			data[4341] <= 8'h10 ;
			data[4342] <= 8'h10 ;
			data[4343] <= 8'h10 ;
			data[4344] <= 8'h10 ;
			data[4345] <= 8'h10 ;
			data[4346] <= 8'h10 ;
			data[4347] <= 8'h10 ;
			data[4348] <= 8'h10 ;
			data[4349] <= 8'h10 ;
			data[4350] <= 8'h10 ;
			data[4351] <= 8'h10 ;
			data[4352] <= 8'h10 ;
			data[4353] <= 8'h10 ;
			data[4354] <= 8'h10 ;
			data[4355] <= 8'h10 ;
			data[4356] <= 8'h10 ;
			data[4357] <= 8'h10 ;
			data[4358] <= 8'h10 ;
			data[4359] <= 8'h10 ;
			data[4360] <= 8'h10 ;
			data[4361] <= 8'h10 ;
			data[4362] <= 8'h10 ;
			data[4363] <= 8'h10 ;
			data[4364] <= 8'h10 ;
			data[4365] <= 8'h10 ;
			data[4366] <= 8'h10 ;
			data[4367] <= 8'h10 ;
			data[4368] <= 8'h10 ;
			data[4369] <= 8'h10 ;
			data[4370] <= 8'h10 ;
			data[4371] <= 8'h10 ;
			data[4372] <= 8'h10 ;
			data[4373] <= 8'h10 ;
			data[4374] <= 8'h10 ;
			data[4375] <= 8'h10 ;
			data[4376] <= 8'h10 ;
			data[4377] <= 8'h10 ;
			data[4378] <= 8'h10 ;
			data[4379] <= 8'h10 ;
			data[4380] <= 8'h10 ;
			data[4381] <= 8'h10 ;
			data[4382] <= 8'h10 ;
			data[4383] <= 8'h10 ;
			data[4384] <= 8'h10 ;
			data[4385] <= 8'h10 ;
			data[4386] <= 8'h10 ;
			data[4387] <= 8'h10 ;
			data[4388] <= 8'h10 ;
			data[4389] <= 8'h10 ;
			data[4390] <= 8'h10 ;
			data[4391] <= 8'h10 ;
			data[4392] <= 8'h10 ;
			data[4393] <= 8'h10 ;
			data[4394] <= 8'h10 ;
			data[4395] <= 8'h10 ;
			data[4396] <= 8'h10 ;
			data[4397] <= 8'h10 ;
			data[4398] <= 8'h10 ;
			data[4399] <= 8'h10 ;
			data[4400] <= 8'h10 ;
			data[4401] <= 8'h10 ;
			data[4402] <= 8'h10 ;
			data[4403] <= 8'h10 ;
			data[4404] <= 8'h10 ;
			data[4405] <= 8'h10 ;
			data[4406] <= 8'h10 ;
			data[4407] <= 8'h10 ;
			data[4408] <= 8'h10 ;
			data[4409] <= 8'h10 ;
			data[4410] <= 8'h10 ;
			data[4411] <= 8'h10 ;
			data[4412] <= 8'h10 ;
			data[4413] <= 8'h10 ;
			data[4414] <= 8'h10 ;
			data[4415] <= 8'h10 ;
			data[4416] <= 8'h10 ;
			data[4417] <= 8'h10 ;
			data[4418] <= 8'h10 ;
			data[4419] <= 8'h10 ;
			data[4420] <= 8'h10 ;
			data[4421] <= 8'h10 ;
			data[4422] <= 8'h10 ;
			data[4423] <= 8'h10 ;
			data[4424] <= 8'h10 ;
			data[4425] <= 8'h10 ;
			data[4426] <= 8'h10 ;
			data[4427] <= 8'h10 ;
			data[4428] <= 8'h10 ;
			data[4429] <= 8'h10 ;
			data[4430] <= 8'h10 ;
			data[4431] <= 8'h10 ;
			data[4432] <= 8'h10 ;
			data[4433] <= 8'h10 ;
			data[4434] <= 8'h10 ;
			data[4435] <= 8'h10 ;
			data[4436] <= 8'h10 ;
			data[4437] <= 8'h10 ;
			data[4438] <= 8'h10 ;
			data[4439] <= 8'h10 ;
			data[4440] <= 8'h10 ;
			data[4441] <= 8'h10 ;
			data[4442] <= 8'h10 ;
			data[4443] <= 8'h10 ;
			data[4444] <= 8'h10 ;
			data[4445] <= 8'h10 ;
			data[4446] <= 8'h10 ;
			data[4447] <= 8'h10 ;
			data[4448] <= 8'h10 ;
			data[4449] <= 8'h10 ;
			data[4450] <= 8'h10 ;
			data[4451] <= 8'h10 ;
			data[4452] <= 8'h10 ;
			data[4453] <= 8'h10 ;
			data[4454] <= 8'h10 ;
			data[4455] <= 8'h10 ;
			data[4456] <= 8'h10 ;
			data[4457] <= 8'h10 ;
			data[4458] <= 8'h10 ;
			data[4459] <= 8'h10 ;
			data[4460] <= 8'h10 ;
			data[4461] <= 8'h10 ;
			data[4462] <= 8'h10 ;
			data[4463] <= 8'h10 ;
			data[4464] <= 8'h10 ;
			data[4465] <= 8'h10 ;
			data[4466] <= 8'h10 ;
			data[4467] <= 8'h10 ;
			data[4468] <= 8'h10 ;
			data[4469] <= 8'h10 ;
			data[4470] <= 8'h10 ;
			data[4471] <= 8'h10 ;
			data[4472] <= 8'h10 ;
			data[4473] <= 8'h10 ;
			data[4474] <= 8'h10 ;
			data[4475] <= 8'h10 ;
			data[4476] <= 8'h10 ;
			data[4477] <= 8'h10 ;
			data[4478] <= 8'h10 ;
			data[4479] <= 8'h10 ;
			data[4480] <= 8'h10 ;
			data[4481] <= 8'h10 ;
			data[4482] <= 8'h10 ;
			data[4483] <= 8'h10 ;
			data[4484] <= 8'h10 ;
			data[4485] <= 8'h10 ;
			data[4486] <= 8'h10 ;
			data[4487] <= 8'h10 ;
			data[4488] <= 8'h10 ;
			data[4489] <= 8'h10 ;
			data[4490] <= 8'h10 ;
			data[4491] <= 8'h10 ;
			data[4492] <= 8'h10 ;
			data[4493] <= 8'h10 ;
			data[4494] <= 8'h10 ;
			data[4495] <= 8'h10 ;
			data[4496] <= 8'h10 ;
			data[4497] <= 8'h10 ;
			data[4498] <= 8'h10 ;
			data[4499] <= 8'h10 ;
			data[4500] <= 8'h10 ;
			data[4501] <= 8'h10 ;
			data[4502] <= 8'h10 ;
			data[4503] <= 8'h10 ;
			data[4504] <= 8'h10 ;
			data[4505] <= 8'h10 ;
			data[4506] <= 8'h10 ;
			data[4507] <= 8'h10 ;
			data[4508] <= 8'h10 ;
			data[4509] <= 8'h10 ;
			data[4510] <= 8'h10 ;
			data[4511] <= 8'h10 ;
			data[4512] <= 8'h10 ;
			data[4513] <= 8'h10 ;
			data[4514] <= 8'h10 ;
			data[4515] <= 8'h10 ;
			data[4516] <= 8'h10 ;
			data[4517] <= 8'h10 ;
			data[4518] <= 8'h10 ;
			data[4519] <= 8'h10 ;
			data[4520] <= 8'h10 ;
			data[4521] <= 8'h10 ;
			data[4522] <= 8'h10 ;
			data[4523] <= 8'h10 ;
			data[4524] <= 8'h10 ;
			data[4525] <= 8'h10 ;
			data[4526] <= 8'h10 ;
			data[4527] <= 8'h10 ;
			data[4528] <= 8'h10 ;
			data[4529] <= 8'h10 ;
			data[4530] <= 8'h10 ;
			data[4531] <= 8'h10 ;
			data[4532] <= 8'h10 ;
			data[4533] <= 8'h10 ;
			data[4534] <= 8'h10 ;
			data[4535] <= 8'h10 ;
			data[4536] <= 8'h10 ;
			data[4537] <= 8'h10 ;
			data[4538] <= 8'h10 ;
			data[4539] <= 8'h10 ;
			data[4540] <= 8'h10 ;
			data[4541] <= 8'h10 ;
			data[4542] <= 8'h10 ;
			data[4543] <= 8'h10 ;
			data[4544] <= 8'h10 ;
			data[4545] <= 8'h10 ;
			data[4546] <= 8'h10 ;
			data[4547] <= 8'h10 ;
			data[4548] <= 8'h10 ;
			data[4549] <= 8'h10 ;
			data[4550] <= 8'h10 ;
			data[4551] <= 8'h10 ;
			data[4552] <= 8'h10 ;
			data[4553] <= 8'h10 ;
			data[4554] <= 8'h10 ;
			data[4555] <= 8'h10 ;
			data[4556] <= 8'h10 ;
			data[4557] <= 8'h10 ;
			data[4558] <= 8'h10 ;
			data[4559] <= 8'h10 ;
			data[4560] <= 8'h10 ;
			data[4561] <= 8'h10 ;
			data[4562] <= 8'h10 ;
			data[4563] <= 8'h10 ;
			data[4564] <= 8'h10 ;
			data[4565] <= 8'h10 ;
			data[4566] <= 8'h10 ;
			data[4567] <= 8'h10 ;
			data[4568] <= 8'h10 ;
			data[4569] <= 8'h10 ;
			data[4570] <= 8'h10 ;
			data[4571] <= 8'h10 ;
			data[4572] <= 8'h10 ;
			data[4573] <= 8'h10 ;
			data[4574] <= 8'h10 ;
			data[4575] <= 8'h10 ;
			data[4576] <= 8'h10 ;
			data[4577] <= 8'h10 ;
			data[4578] <= 8'h10 ;
			data[4579] <= 8'h10 ;
			data[4580] <= 8'h10 ;
			data[4581] <= 8'h10 ;
			data[4582] <= 8'h10 ;
			data[4583] <= 8'h10 ;
			data[4584] <= 8'h10 ;
			data[4585] <= 8'h10 ;
			data[4586] <= 8'h10 ;
			data[4587] <= 8'h10 ;
			data[4588] <= 8'h10 ;
			data[4589] <= 8'h10 ;
			data[4590] <= 8'h10 ;
			data[4591] <= 8'h10 ;
			data[4592] <= 8'h10 ;
			data[4593] <= 8'h10 ;
			data[4594] <= 8'h10 ;
			data[4595] <= 8'h10 ;
			data[4596] <= 8'h10 ;
			data[4597] <= 8'h10 ;
			data[4598] <= 8'h10 ;
			data[4599] <= 8'h10 ;
			data[4600] <= 8'h10 ;
			data[4601] <= 8'h10 ;
			data[4602] <= 8'h10 ;
			data[4603] <= 8'h10 ;
			data[4604] <= 8'h10 ;
			data[4605] <= 8'h10 ;
			data[4606] <= 8'h10 ;
			data[4607] <= 8'h10 ;
			data[4608] <= 8'h10 ;
			data[4609] <= 8'h10 ;
			data[4610] <= 8'h10 ;
			data[4611] <= 8'h10 ;
			data[4612] <= 8'h10 ;
			data[4613] <= 8'h10 ;
			data[4614] <= 8'h10 ;
			data[4615] <= 8'h10 ;
			data[4616] <= 8'h10 ;
			data[4617] <= 8'h10 ;
			data[4618] <= 8'h10 ;
			data[4619] <= 8'h10 ;
			data[4620] <= 8'h10 ;
			data[4621] <= 8'h10 ;
			data[4622] <= 8'h10 ;
			data[4623] <= 8'h10 ;
			data[4624] <= 8'h10 ;
			data[4625] <= 8'h10 ;
			data[4626] <= 8'h10 ;
			data[4627] <= 8'h10 ;
			data[4628] <= 8'h10 ;
			data[4629] <= 8'h10 ;
			data[4630] <= 8'h10 ;
			data[4631] <= 8'h10 ;
			data[4632] <= 8'h10 ;
			data[4633] <= 8'h10 ;
			data[4634] <= 8'h10 ;
			data[4635] <= 8'h10 ;
			data[4636] <= 8'h10 ;
			data[4637] <= 8'h10 ;
			data[4638] <= 8'h10 ;
			data[4639] <= 8'h10 ;
			data[4640] <= 8'h10 ;
			data[4641] <= 8'h10 ;
			data[4642] <= 8'h10 ;
			data[4643] <= 8'h10 ;
			data[4644] <= 8'h10 ;
			data[4645] <= 8'h10 ;
			data[4646] <= 8'h10 ;
			data[4647] <= 8'h10 ;
			data[4648] <= 8'h10 ;
			data[4649] <= 8'h10 ;
			data[4650] <= 8'h10 ;
			data[4651] <= 8'h10 ;
			data[4652] <= 8'h10 ;
			data[4653] <= 8'h10 ;
			data[4654] <= 8'h10 ;
			data[4655] <= 8'h10 ;
			data[4656] <= 8'h10 ;
			data[4657] <= 8'h10 ;
			data[4658] <= 8'h10 ;
			data[4659] <= 8'h10 ;
			data[4660] <= 8'h10 ;
			data[4661] <= 8'h10 ;
			data[4662] <= 8'h10 ;
			data[4663] <= 8'h10 ;
			data[4664] <= 8'h10 ;
			data[4665] <= 8'h10 ;
			data[4666] <= 8'h10 ;
			data[4667] <= 8'h10 ;
			data[4668] <= 8'h10 ;
			data[4669] <= 8'h10 ;
			data[4670] <= 8'h10 ;
			data[4671] <= 8'h10 ;
			data[4672] <= 8'h10 ;
			data[4673] <= 8'h10 ;
			data[4674] <= 8'h10 ;
			data[4675] <= 8'h10 ;
			data[4676] <= 8'h10 ;
			data[4677] <= 8'h10 ;
			data[4678] <= 8'h10 ;
			data[4679] <= 8'h10 ;
			data[4680] <= 8'h10 ;
			data[4681] <= 8'h10 ;
			data[4682] <= 8'h10 ;
			data[4683] <= 8'h10 ;
			data[4684] <= 8'h10 ;
			data[4685] <= 8'h10 ;
			data[4686] <= 8'h10 ;
			data[4687] <= 8'h10 ;
			data[4688] <= 8'h10 ;
			data[4689] <= 8'h10 ;
			data[4690] <= 8'h10 ;
			data[4691] <= 8'h10 ;
			data[4692] <= 8'h10 ;
			data[4693] <= 8'h10 ;
			data[4694] <= 8'h10 ;
			data[4695] <= 8'h10 ;
			data[4696] <= 8'h10 ;
			data[4697] <= 8'h10 ;
			data[4698] <= 8'h10 ;
			data[4699] <= 8'h10 ;
			data[4700] <= 8'h10 ;
			data[4701] <= 8'h10 ;
			data[4702] <= 8'h10 ;
			data[4703] <= 8'h10 ;
			data[4704] <= 8'h10 ;
			data[4705] <= 8'h10 ;
			data[4706] <= 8'h10 ;
			data[4707] <= 8'h10 ;
			data[4708] <= 8'h10 ;
			data[4709] <= 8'h10 ;
			data[4710] <= 8'h10 ;
			data[4711] <= 8'h10 ;
			data[4712] <= 8'h10 ;
			data[4713] <= 8'h10 ;
			data[4714] <= 8'h10 ;
			data[4715] <= 8'h10 ;
			data[4716] <= 8'h10 ;
			data[4717] <= 8'h10 ;
			data[4718] <= 8'h10 ;
			data[4719] <= 8'h10 ;
			data[4720] <= 8'h10 ;
			data[4721] <= 8'h10 ;
			data[4722] <= 8'h10 ;
			data[4723] <= 8'h10 ;
			data[4724] <= 8'h10 ;
			data[4725] <= 8'h10 ;
			data[4726] <= 8'h10 ;
			data[4727] <= 8'h10 ;
			data[4728] <= 8'h10 ;
			data[4729] <= 8'h10 ;
			data[4730] <= 8'h10 ;
			data[4731] <= 8'h10 ;
			data[4732] <= 8'h10 ;
			data[4733] <= 8'h10 ;
			data[4734] <= 8'h10 ;
			data[4735] <= 8'h10 ;
			data[4736] <= 8'h10 ;
			data[4737] <= 8'h10 ;
			data[4738] <= 8'h10 ;
			data[4739] <= 8'h10 ;
			data[4740] <= 8'h10 ;
			data[4741] <= 8'h10 ;
			data[4742] <= 8'h10 ;
			data[4743] <= 8'h10 ;
			data[4744] <= 8'h10 ;
			data[4745] <= 8'h10 ;
			data[4746] <= 8'h10 ;
			data[4747] <= 8'h10 ;
			data[4748] <= 8'h10 ;
			data[4749] <= 8'h10 ;
			data[4750] <= 8'h10 ;
			data[4751] <= 8'h10 ;
			data[4752] <= 8'h10 ;
			data[4753] <= 8'h10 ;
			data[4754] <= 8'h10 ;
			data[4755] <= 8'h10 ;
			data[4756] <= 8'h10 ;
			data[4757] <= 8'h10 ;
			data[4758] <= 8'h10 ;
			data[4759] <= 8'h10 ;
			data[4760] <= 8'h10 ;
			data[4761] <= 8'h10 ;
			data[4762] <= 8'h10 ;
			data[4763] <= 8'h10 ;
			data[4764] <= 8'h10 ;
			data[4765] <= 8'h10 ;
			data[4766] <= 8'h10 ;
			data[4767] <= 8'h10 ;
			data[4768] <= 8'h10 ;
			data[4769] <= 8'h10 ;
			data[4770] <= 8'h10 ;
			data[4771] <= 8'h10 ;
			data[4772] <= 8'h10 ;
			data[4773] <= 8'h10 ;
			data[4774] <= 8'h10 ;
			data[4775] <= 8'h10 ;
			data[4776] <= 8'h10 ;
			data[4777] <= 8'h10 ;
			data[4778] <= 8'h10 ;
			data[4779] <= 8'h10 ;
			data[4780] <= 8'h10 ;
			data[4781] <= 8'h10 ;
			data[4782] <= 8'h10 ;
			data[4783] <= 8'h10 ;
			data[4784] <= 8'h10 ;
			data[4785] <= 8'h10 ;
			data[4786] <= 8'h10 ;
			data[4787] <= 8'h10 ;
			data[4788] <= 8'h10 ;
			data[4789] <= 8'h10 ;
			data[4790] <= 8'h10 ;
			data[4791] <= 8'h10 ;
			data[4792] <= 8'h10 ;
			data[4793] <= 8'h10 ;
			data[4794] <= 8'h10 ;
			data[4795] <= 8'h10 ;
			data[4796] <= 8'h10 ;
			data[4797] <= 8'h10 ;
			data[4798] <= 8'h10 ;
			data[4799] <= 8'h10 ;
			data[4800] <= 8'h10 ;
			data[4801] <= 8'h10 ;
			data[4802] <= 8'h10 ;
			data[4803] <= 8'h10 ;
			data[4804] <= 8'h10 ;
			data[4805] <= 8'h10 ;
			data[4806] <= 8'h10 ;
			data[4807] <= 8'h10 ;
			data[4808] <= 8'h10 ;
			data[4809] <= 8'h10 ;
			data[4810] <= 8'h10 ;
			data[4811] <= 8'h10 ;
			data[4812] <= 8'h10 ;
			data[4813] <= 8'h10 ;
			data[4814] <= 8'h10 ;
			data[4815] <= 8'h10 ;
			data[4816] <= 8'h10 ;
			data[4817] <= 8'h10 ;
			data[4818] <= 8'h10 ;
			data[4819] <= 8'h10 ;
			data[4820] <= 8'h10 ;
			data[4821] <= 8'h10 ;
			data[4822] <= 8'h10 ;
			data[4823] <= 8'h10 ;
			data[4824] <= 8'h10 ;
			data[4825] <= 8'h10 ;
			data[4826] <= 8'h10 ;
			data[4827] <= 8'h10 ;
			data[4828] <= 8'h10 ;
			data[4829] <= 8'h10 ;
			data[4830] <= 8'h10 ;
			data[4831] <= 8'h10 ;
			data[4832] <= 8'h10 ;
			data[4833] <= 8'h10 ;
			data[4834] <= 8'h10 ;
			data[4835] <= 8'h10 ;
			data[4836] <= 8'h10 ;
			data[4837] <= 8'h10 ;
			data[4838] <= 8'h10 ;
			data[4839] <= 8'h10 ;
			data[4840] <= 8'h10 ;
			data[4841] <= 8'h10 ;
			data[4842] <= 8'h10 ;
			data[4843] <= 8'h10 ;
			data[4844] <= 8'h10 ;
			data[4845] <= 8'h10 ;
			data[4846] <= 8'h10 ;
			data[4847] <= 8'h10 ;
			data[4848] <= 8'h10 ;
			data[4849] <= 8'h10 ;
			data[4850] <= 8'h10 ;
			data[4851] <= 8'h10 ;
			data[4852] <= 8'h10 ;
			data[4853] <= 8'h10 ;
			data[4854] <= 8'h10 ;
			data[4855] <= 8'h10 ;
			data[4856] <= 8'h10 ;
			data[4857] <= 8'h10 ;
			data[4858] <= 8'h10 ;
			data[4859] <= 8'h10 ;
			data[4860] <= 8'h10 ;
			data[4861] <= 8'h10 ;
			data[4862] <= 8'h10 ;
			data[4863] <= 8'h10 ;
			data[4864] <= 8'h10 ;
			data[4865] <= 8'h10 ;
			data[4866] <= 8'h10 ;
			data[4867] <= 8'h10 ;
			data[4868] <= 8'h10 ;
			data[4869] <= 8'h10 ;
			data[4870] <= 8'h10 ;
			data[4871] <= 8'h10 ;
			data[4872] <= 8'h10 ;
			data[4873] <= 8'h10 ;
			data[4874] <= 8'h10 ;
			data[4875] <= 8'h10 ;
			data[4876] <= 8'h10 ;
			data[4877] <= 8'h10 ;
			data[4878] <= 8'h10 ;
			data[4879] <= 8'h10 ;
			data[4880] <= 8'h10 ;
			data[4881] <= 8'h10 ;
			data[4882] <= 8'h10 ;
			data[4883] <= 8'h10 ;
			data[4884] <= 8'h10 ;
			data[4885] <= 8'h10 ;
			data[4886] <= 8'h10 ;
			data[4887] <= 8'h10 ;
			data[4888] <= 8'h10 ;
			data[4889] <= 8'h10 ;
			data[4890] <= 8'h10 ;
			data[4891] <= 8'h10 ;
			data[4892] <= 8'h10 ;
			data[4893] <= 8'h10 ;
			data[4894] <= 8'h10 ;
			data[4895] <= 8'h10 ;
			data[4896] <= 8'h10 ;
			data[4897] <= 8'h10 ;
			data[4898] <= 8'h10 ;
			data[4899] <= 8'h10 ;
			data[4900] <= 8'h10 ;
			data[4901] <= 8'h10 ;
			data[4902] <= 8'h10 ;
			data[4903] <= 8'h10 ;
			data[4904] <= 8'h10 ;
			data[4905] <= 8'h10 ;
			data[4906] <= 8'h10 ;
			data[4907] <= 8'h10 ;
			data[4908] <= 8'h10 ;
			data[4909] <= 8'h10 ;
			data[4910] <= 8'h10 ;
			data[4911] <= 8'h10 ;
			data[4912] <= 8'h10 ;
			data[4913] <= 8'h10 ;
			data[4914] <= 8'h10 ;
			data[4915] <= 8'h10 ;
			data[4916] <= 8'h10 ;
			data[4917] <= 8'h10 ;
			data[4918] <= 8'h10 ;
			data[4919] <= 8'h10 ;
			data[4920] <= 8'h10 ;
			data[4921] <= 8'h10 ;
			data[4922] <= 8'h10 ;
			data[4923] <= 8'h10 ;
			data[4924] <= 8'h10 ;
			data[4925] <= 8'h10 ;
			data[4926] <= 8'h10 ;
			data[4927] <= 8'h10 ;
			data[4928] <= 8'h10 ;
			data[4929] <= 8'h10 ;
			data[4930] <= 8'h10 ;
			data[4931] <= 8'h10 ;
			data[4932] <= 8'h10 ;
			data[4933] <= 8'h10 ;
			data[4934] <= 8'h10 ;
			data[4935] <= 8'h10 ;
			data[4936] <= 8'h10 ;
			data[4937] <= 8'h10 ;
			data[4938] <= 8'h10 ;
			data[4939] <= 8'h10 ;
			data[4940] <= 8'h10 ;
			data[4941] <= 8'h10 ;
			data[4942] <= 8'h10 ;
			data[4943] <= 8'h10 ;
			data[4944] <= 8'h10 ;
			data[4945] <= 8'h10 ;
			data[4946] <= 8'h10 ;
			data[4947] <= 8'h10 ;
			data[4948] <= 8'h10 ;
			data[4949] <= 8'h10 ;
			data[4950] <= 8'h10 ;
			data[4951] <= 8'h10 ;
			data[4952] <= 8'h10 ;
			data[4953] <= 8'h10 ;
			data[4954] <= 8'h10 ;
			data[4955] <= 8'h10 ;
			data[4956] <= 8'h10 ;
			data[4957] <= 8'h10 ;
			data[4958] <= 8'h10 ;
			data[4959] <= 8'h10 ;
			data[4960] <= 8'h10 ;
			data[4961] <= 8'h10 ;
			data[4962] <= 8'h10 ;
			data[4963] <= 8'h10 ;
			data[4964] <= 8'h10 ;
			data[4965] <= 8'h10 ;
			data[4966] <= 8'h10 ;
			data[4967] <= 8'h10 ;
			data[4968] <= 8'h10 ;
			data[4969] <= 8'h10 ;
			data[4970] <= 8'h10 ;
			data[4971] <= 8'h10 ;
			data[4972] <= 8'h10 ;
			data[4973] <= 8'h10 ;
			data[4974] <= 8'h10 ;
			data[4975] <= 8'h10 ;
			data[4976] <= 8'h10 ;
			data[4977] <= 8'h10 ;
			data[4978] <= 8'h10 ;
			data[4979] <= 8'h10 ;
			data[4980] <= 8'h10 ;
			data[4981] <= 8'h10 ;
			data[4982] <= 8'h10 ;
			data[4983] <= 8'h10 ;
			data[4984] <= 8'h10 ;
			data[4985] <= 8'h10 ;
			data[4986] <= 8'h10 ;
			data[4987] <= 8'h10 ;
			data[4988] <= 8'h10 ;
			data[4989] <= 8'h10 ;
			data[4990] <= 8'h10 ;
			data[4991] <= 8'h10 ;
			data[4992] <= 8'h10 ;
			data[4993] <= 8'h10 ;
			data[4994] <= 8'h10 ;
			data[4995] <= 8'h10 ;
			data[4996] <= 8'h10 ;
			data[4997] <= 8'h10 ;
			data[4998] <= 8'h10 ;
			data[4999] <= 8'h10 ;
			data[5000] <= 8'h10 ;
			data[5001] <= 8'h10 ;
			data[5002] <= 8'h10 ;
			data[5003] <= 8'h10 ;
			data[5004] <= 8'h10 ;
			data[5005] <= 8'h10 ;
			data[5006] <= 8'h10 ;
			data[5007] <= 8'h10 ;
			data[5008] <= 8'h10 ;
			data[5009] <= 8'h10 ;
			data[5010] <= 8'h10 ;
			data[5011] <= 8'h10 ;
			data[5012] <= 8'h10 ;
			data[5013] <= 8'h10 ;
			data[5014] <= 8'h10 ;
			data[5015] <= 8'h10 ;
			data[5016] <= 8'h10 ;
			data[5017] <= 8'h10 ;
			data[5018] <= 8'h10 ;
			data[5019] <= 8'h10 ;
			data[5020] <= 8'h10 ;
			data[5021] <= 8'h10 ;
			data[5022] <= 8'h10 ;
			data[5023] <= 8'h10 ;
			data[5024] <= 8'h10 ;
			data[5025] <= 8'h10 ;
			data[5026] <= 8'h10 ;
			data[5027] <= 8'h10 ;
			data[5028] <= 8'h10 ;
			data[5029] <= 8'h10 ;
			data[5030] <= 8'h10 ;
			data[5031] <= 8'h10 ;
			data[5032] <= 8'h10 ;
			data[5033] <= 8'h10 ;
			data[5034] <= 8'h10 ;
			data[5035] <= 8'h10 ;
			data[5036] <= 8'h10 ;
			data[5037] <= 8'h10 ;
			data[5038] <= 8'h10 ;
			data[5039] <= 8'h10 ;
			data[5040] <= 8'h10 ;
			data[5041] <= 8'h10 ;
			data[5042] <= 8'h10 ;
			data[5043] <= 8'h10 ;
			data[5044] <= 8'h10 ;
			data[5045] <= 8'h10 ;
			data[5046] <= 8'h10 ;
			data[5047] <= 8'h10 ;
			data[5048] <= 8'h10 ;
			data[5049] <= 8'h10 ;
			data[5050] <= 8'h10 ;
			data[5051] <= 8'h10 ;
			data[5052] <= 8'h10 ;
			data[5053] <= 8'h10 ;
			data[5054] <= 8'h10 ;
			data[5055] <= 8'h10 ;
			data[5056] <= 8'h10 ;
			data[5057] <= 8'h10 ;
			data[5058] <= 8'h10 ;
			data[5059] <= 8'h10 ;
			data[5060] <= 8'h10 ;
			data[5061] <= 8'h10 ;
			data[5062] <= 8'h10 ;
			data[5063] <= 8'h10 ;
			data[5064] <= 8'h10 ;
			data[5065] <= 8'h10 ;
			data[5066] <= 8'h10 ;
			data[5067] <= 8'h10 ;
			data[5068] <= 8'h10 ;
			data[5069] <= 8'h10 ;
			data[5070] <= 8'h10 ;
			data[5071] <= 8'h10 ;
			data[5072] <= 8'h10 ;
			data[5073] <= 8'h10 ;
			data[5074] <= 8'h10 ;
			data[5075] <= 8'h10 ;
			data[5076] <= 8'h10 ;
			data[5077] <= 8'h10 ;
			data[5078] <= 8'h10 ;
			data[5079] <= 8'h10 ;
			data[5080] <= 8'h10 ;
			data[5081] <= 8'h10 ;
			data[5082] <= 8'h10 ;
			data[5083] <= 8'h10 ;
			data[5084] <= 8'h10 ;
			data[5085] <= 8'h10 ;
			data[5086] <= 8'h10 ;
			data[5087] <= 8'h10 ;
			data[5088] <= 8'h10 ;
			data[5089] <= 8'h10 ;
			data[5090] <= 8'h10 ;
			data[5091] <= 8'h10 ;
			data[5092] <= 8'h10 ;
			data[5093] <= 8'h10 ;
			data[5094] <= 8'h10 ;
			data[5095] <= 8'h10 ;
			data[5096] <= 8'h10 ;
			data[5097] <= 8'h10 ;
			data[5098] <= 8'h10 ;
			data[5099] <= 8'h10 ;
			data[5100] <= 8'h10 ;
			data[5101] <= 8'h10 ;
			data[5102] <= 8'h10 ;
			data[5103] <= 8'h10 ;
			data[5104] <= 8'h10 ;
			data[5105] <= 8'h10 ;
			data[5106] <= 8'h10 ;
			data[5107] <= 8'h10 ;
			data[5108] <= 8'h10 ;
			data[5109] <= 8'h10 ;
			data[5110] <= 8'h10 ;
			data[5111] <= 8'h10 ;
			data[5112] <= 8'h10 ;
			data[5113] <= 8'h10 ;
			data[5114] <= 8'h10 ;
			data[5115] <= 8'h10 ;
			data[5116] <= 8'h10 ;
			data[5117] <= 8'h10 ;
			data[5118] <= 8'h10 ;
			data[5119] <= 8'h10 ;
			data[5120] <= 8'h10 ;
			data[5121] <= 8'h10 ;
			data[5122] <= 8'h10 ;
			data[5123] <= 8'h10 ;
			data[5124] <= 8'h10 ;
			data[5125] <= 8'h10 ;
			data[5126] <= 8'h10 ;
			data[5127] <= 8'h10 ;
			data[5128] <= 8'h10 ;
			data[5129] <= 8'h10 ;
			data[5130] <= 8'h10 ;
			data[5131] <= 8'h10 ;
			data[5132] <= 8'h10 ;
			data[5133] <= 8'h10 ;
			data[5134] <= 8'h10 ;
			data[5135] <= 8'h10 ;
			data[5136] <= 8'h10 ;
			data[5137] <= 8'h10 ;
			data[5138] <= 8'h10 ;
			data[5139] <= 8'h10 ;
			data[5140] <= 8'h10 ;
			data[5141] <= 8'h10 ;
			data[5142] <= 8'h10 ;
			data[5143] <= 8'h10 ;
			data[5144] <= 8'h10 ;
			data[5145] <= 8'h10 ;
			data[5146] <= 8'h10 ;
			data[5147] <= 8'h10 ;
			data[5148] <= 8'h10 ;
			data[5149] <= 8'h10 ;
			data[5150] <= 8'h10 ;
			data[5151] <= 8'h10 ;
			data[5152] <= 8'h10 ;
			data[5153] <= 8'h10 ;
			data[5154] <= 8'h10 ;
			data[5155] <= 8'h10 ;
			data[5156] <= 8'h10 ;
			data[5157] <= 8'h10 ;
			data[5158] <= 8'h10 ;
			data[5159] <= 8'h10 ;
			data[5160] <= 8'h10 ;
			data[5161] <= 8'h10 ;
			data[5162] <= 8'h10 ;
			data[5163] <= 8'h10 ;
			data[5164] <= 8'h10 ;
			data[5165] <= 8'h10 ;
			data[5166] <= 8'h10 ;
			data[5167] <= 8'h10 ;
			data[5168] <= 8'h10 ;
			data[5169] <= 8'h10 ;
			data[5170] <= 8'h10 ;
			data[5171] <= 8'h10 ;
			data[5172] <= 8'h10 ;
			data[5173] <= 8'h10 ;
			data[5174] <= 8'h10 ;
			data[5175] <= 8'h10 ;
			data[5176] <= 8'h10 ;
			data[5177] <= 8'h10 ;
			data[5178] <= 8'h10 ;
			data[5179] <= 8'h10 ;
			data[5180] <= 8'h10 ;
			data[5181] <= 8'h10 ;
			data[5182] <= 8'h10 ;
			data[5183] <= 8'h10 ;
			data[5184] <= 8'h10 ;
			data[5185] <= 8'h10 ;
			data[5186] <= 8'h10 ;
			data[5187] <= 8'h10 ;
			data[5188] <= 8'h10 ;
			data[5189] <= 8'h10 ;
			data[5190] <= 8'h10 ;
			data[5191] <= 8'h10 ;
			data[5192] <= 8'h10 ;
			data[5193] <= 8'h10 ;
			data[5194] <= 8'h10 ;
			data[5195] <= 8'h10 ;
			data[5196] <= 8'h10 ;
			data[5197] <= 8'h10 ;
			data[5198] <= 8'h10 ;
			data[5199] <= 8'h10 ;
			data[5200] <= 8'h10 ;
			data[5201] <= 8'h10 ;
			data[5202] <= 8'h10 ;
			data[5203] <= 8'h10 ;
			data[5204] <= 8'h10 ;
			data[5205] <= 8'h10 ;
			data[5206] <= 8'h10 ;
			data[5207] <= 8'h10 ;
			data[5208] <= 8'h10 ;
			data[5209] <= 8'h10 ;
			data[5210] <= 8'h10 ;
			data[5211] <= 8'h10 ;
			data[5212] <= 8'h10 ;
			data[5213] <= 8'h10 ;
			data[5214] <= 8'h10 ;
			data[5215] <= 8'h10 ;
			data[5216] <= 8'h10 ;
			data[5217] <= 8'h10 ;
			data[5218] <= 8'h10 ;
			data[5219] <= 8'h10 ;
			data[5220] <= 8'h10 ;
			data[5221] <= 8'h10 ;
			data[5222] <= 8'h10 ;
			data[5223] <= 8'h10 ;
			data[5224] <= 8'h10 ;
			data[5225] <= 8'h10 ;
			data[5226] <= 8'h10 ;
			data[5227] <= 8'h10 ;
			data[5228] <= 8'h10 ;
			data[5229] <= 8'h10 ;
			data[5230] <= 8'h10 ;
			data[5231] <= 8'h10 ;
			data[5232] <= 8'h10 ;
			data[5233] <= 8'h10 ;
			data[5234] <= 8'h10 ;
			data[5235] <= 8'h10 ;
			data[5236] <= 8'h10 ;
			data[5237] <= 8'h10 ;
			data[5238] <= 8'h10 ;
			data[5239] <= 8'h10 ;
			data[5240] <= 8'h10 ;
			data[5241] <= 8'h10 ;
			data[5242] <= 8'h10 ;
			data[5243] <= 8'h10 ;
			data[5244] <= 8'h10 ;
			data[5245] <= 8'h10 ;
			data[5246] <= 8'h10 ;
			data[5247] <= 8'h10 ;
			data[5248] <= 8'h10 ;
			data[5249] <= 8'h10 ;
			data[5250] <= 8'h10 ;
			data[5251] <= 8'h10 ;
			data[5252] <= 8'h10 ;
			data[5253] <= 8'h10 ;
			data[5254] <= 8'h10 ;
			data[5255] <= 8'h10 ;
			data[5256] <= 8'h10 ;
			data[5257] <= 8'h10 ;
			data[5258] <= 8'h10 ;
			data[5259] <= 8'h10 ;
			data[5260] <= 8'h10 ;
			data[5261] <= 8'h10 ;
			data[5262] <= 8'h10 ;
			data[5263] <= 8'h10 ;
			data[5264] <= 8'h10 ;
			data[5265] <= 8'h10 ;
			data[5266] <= 8'h10 ;
			data[5267] <= 8'h10 ;
			data[5268] <= 8'h10 ;
			data[5269] <= 8'h10 ;
			data[5270] <= 8'h10 ;
			data[5271] <= 8'h10 ;
			data[5272] <= 8'h10 ;
			data[5273] <= 8'h10 ;
			data[5274] <= 8'h10 ;
			data[5275] <= 8'h10 ;
			data[5276] <= 8'h10 ;
			data[5277] <= 8'h10 ;
			data[5278] <= 8'h10 ;
			data[5279] <= 8'h10 ;
			data[5280] <= 8'h10 ;
			data[5281] <= 8'h10 ;
			data[5282] <= 8'h10 ;
			data[5283] <= 8'h10 ;
			data[5284] <= 8'h10 ;
			data[5285] <= 8'h10 ;
			data[5286] <= 8'h10 ;
			data[5287] <= 8'h10 ;
			data[5288] <= 8'h10 ;
			data[5289] <= 8'h10 ;
			data[5290] <= 8'h10 ;
			data[5291] <= 8'h10 ;
			data[5292] <= 8'h10 ;
			data[5293] <= 8'h10 ;
			data[5294] <= 8'h10 ;
			data[5295] <= 8'h10 ;
			data[5296] <= 8'h10 ;
			data[5297] <= 8'h10 ;
			data[5298] <= 8'h10 ;
			data[5299] <= 8'h10 ;
			data[5300] <= 8'h10 ;
			data[5301] <= 8'h10 ;
			data[5302] <= 8'h10 ;
			data[5303] <= 8'h10 ;
			data[5304] <= 8'h10 ;
			data[5305] <= 8'h10 ;
			data[5306] <= 8'h10 ;
			data[5307] <= 8'h10 ;
			data[5308] <= 8'h10 ;
			data[5309] <= 8'h10 ;
			data[5310] <= 8'h10 ;
			data[5311] <= 8'h10 ;
			data[5312] <= 8'h10 ;
			data[5313] <= 8'h10 ;
			data[5314] <= 8'h10 ;
			data[5315] <= 8'h10 ;
			data[5316] <= 8'h10 ;
			data[5317] <= 8'h10 ;
			data[5318] <= 8'h10 ;
			data[5319] <= 8'h10 ;
			data[5320] <= 8'h10 ;
			data[5321] <= 8'h10 ;
			data[5322] <= 8'h10 ;
			data[5323] <= 8'h10 ;
			data[5324] <= 8'h10 ;
			data[5325] <= 8'h10 ;
			data[5326] <= 8'h10 ;
			data[5327] <= 8'h10 ;
			data[5328] <= 8'h10 ;
			data[5329] <= 8'h10 ;
			data[5330] <= 8'h10 ;
			data[5331] <= 8'h10 ;
			data[5332] <= 8'h10 ;
			data[5333] <= 8'h10 ;
			data[5334] <= 8'h10 ;
			data[5335] <= 8'h10 ;
			data[5336] <= 8'h10 ;
			data[5337] <= 8'h10 ;
			data[5338] <= 8'h10 ;
			data[5339] <= 8'h10 ;
			data[5340] <= 8'h10 ;
			data[5341] <= 8'h10 ;
			data[5342] <= 8'h10 ;
			data[5343] <= 8'h10 ;
			data[5344] <= 8'h10 ;
			data[5345] <= 8'h10 ;
			data[5346] <= 8'h10 ;
			data[5347] <= 8'h10 ;
			data[5348] <= 8'h10 ;
			data[5349] <= 8'h10 ;
			data[5350] <= 8'h10 ;
			data[5351] <= 8'h10 ;
			data[5352] <= 8'h10 ;
			data[5353] <= 8'h10 ;
			data[5354] <= 8'h10 ;
			data[5355] <= 8'h10 ;
			data[5356] <= 8'h10 ;
			data[5357] <= 8'h10 ;
			data[5358] <= 8'h10 ;
			data[5359] <= 8'h10 ;
			data[5360] <= 8'h10 ;
			data[5361] <= 8'h10 ;
			data[5362] <= 8'h10 ;
			data[5363] <= 8'h10 ;
			data[5364] <= 8'h10 ;
			data[5365] <= 8'h10 ;
			data[5366] <= 8'h10 ;
			data[5367] <= 8'h10 ;
			data[5368] <= 8'h10 ;
			data[5369] <= 8'h10 ;
			data[5370] <= 8'h10 ;
			data[5371] <= 8'h10 ;
			data[5372] <= 8'h10 ;
			data[5373] <= 8'h10 ;
			data[5374] <= 8'h10 ;
			data[5375] <= 8'h10 ;
			data[5376] <= 8'h10 ;
			data[5377] <= 8'h10 ;
			data[5378] <= 8'h10 ;
			data[5379] <= 8'h10 ;
			data[5380] <= 8'h10 ;
			data[5381] <= 8'h10 ;
			data[5382] <= 8'h10 ;
			data[5383] <= 8'h10 ;
			data[5384] <= 8'h10 ;
			data[5385] <= 8'h10 ;
			data[5386] <= 8'h10 ;
			data[5387] <= 8'h10 ;
			data[5388] <= 8'h10 ;
			data[5389] <= 8'h10 ;
			data[5390] <= 8'h10 ;
			data[5391] <= 8'h10 ;
			data[5392] <= 8'h10 ;
			data[5393] <= 8'h10 ;
			data[5394] <= 8'h10 ;
			data[5395] <= 8'h10 ;
			data[5396] <= 8'h10 ;
			data[5397] <= 8'h10 ;
			data[5398] <= 8'h10 ;
			data[5399] <= 8'h10 ;
			data[5400] <= 8'h10 ;
			data[5401] <= 8'h10 ;
			data[5402] <= 8'h10 ;
			data[5403] <= 8'h10 ;
			data[5404] <= 8'h10 ;
			data[5405] <= 8'h10 ;
			data[5406] <= 8'h10 ;
			data[5407] <= 8'h10 ;
			data[5408] <= 8'h10 ;
			data[5409] <= 8'h10 ;
			data[5410] <= 8'h10 ;
			data[5411] <= 8'h10 ;
			data[5412] <= 8'h10 ;
			data[5413] <= 8'h10 ;
			data[5414] <= 8'h10 ;
			data[5415] <= 8'h10 ;
			data[5416] <= 8'h10 ;
			data[5417] <= 8'h10 ;
			data[5418] <= 8'h10 ;
			data[5419] <= 8'h10 ;
			data[5420] <= 8'h10 ;
			data[5421] <= 8'h10 ;
			data[5422] <= 8'h10 ;
			data[5423] <= 8'h10 ;
			data[5424] <= 8'h10 ;
			data[5425] <= 8'h10 ;
			data[5426] <= 8'h10 ;
			data[5427] <= 8'h10 ;
			data[5428] <= 8'h10 ;
			data[5429] <= 8'h10 ;
			data[5430] <= 8'h10 ;
			data[5431] <= 8'h10 ;
			data[5432] <= 8'h10 ;
			data[5433] <= 8'h10 ;
			data[5434] <= 8'h10 ;
			data[5435] <= 8'h10 ;
			data[5436] <= 8'h10 ;
			data[5437] <= 8'h10 ;
			data[5438] <= 8'h10 ;
			data[5439] <= 8'h10 ;
			data[5440] <= 8'h10 ;
			data[5441] <= 8'h10 ;
			data[5442] <= 8'h10 ;
			data[5443] <= 8'h10 ;
			data[5444] <= 8'h10 ;
			data[5445] <= 8'h10 ;
			data[5446] <= 8'h10 ;
			data[5447] <= 8'h10 ;
			data[5448] <= 8'h10 ;
			data[5449] <= 8'h10 ;
			data[5450] <= 8'h10 ;
			data[5451] <= 8'h10 ;
			data[5452] <= 8'h10 ;
			data[5453] <= 8'h10 ;
			data[5454] <= 8'h10 ;
			data[5455] <= 8'h10 ;
			data[5456] <= 8'h10 ;
			data[5457] <= 8'h10 ;
			data[5458] <= 8'h10 ;
			data[5459] <= 8'h10 ;
			data[5460] <= 8'h10 ;
			data[5461] <= 8'h10 ;
			data[5462] <= 8'h10 ;
			data[5463] <= 8'h10 ;
			data[5464] <= 8'h10 ;
			data[5465] <= 8'h10 ;
			data[5466] <= 8'h10 ;
			data[5467] <= 8'h10 ;
			data[5468] <= 8'h10 ;
			data[5469] <= 8'h10 ;
			data[5470] <= 8'h10 ;
			data[5471] <= 8'h10 ;
			data[5472] <= 8'h10 ;
			data[5473] <= 8'h10 ;
			data[5474] <= 8'h10 ;
			data[5475] <= 8'h10 ;
			data[5476] <= 8'h10 ;
			data[5477] <= 8'h10 ;
			data[5478] <= 8'h10 ;
			data[5479] <= 8'h10 ;
			data[5480] <= 8'h10 ;
			data[5481] <= 8'h10 ;
			data[5482] <= 8'h10 ;
			data[5483] <= 8'h10 ;
			data[5484] <= 8'h10 ;
			data[5485] <= 8'h10 ;
			data[5486] <= 8'h10 ;
			data[5487] <= 8'h10 ;
			data[5488] <= 8'h10 ;
			data[5489] <= 8'h10 ;
			data[5490] <= 8'h10 ;
			data[5491] <= 8'h10 ;
			data[5492] <= 8'h10 ;
			data[5493] <= 8'h10 ;
			data[5494] <= 8'h10 ;
			data[5495] <= 8'h10 ;
			data[5496] <= 8'h10 ;
			data[5497] <= 8'h10 ;
			data[5498] <= 8'h10 ;
			data[5499] <= 8'h10 ;
			data[5500] <= 8'h10 ;
			data[5501] <= 8'h10 ;
			data[5502] <= 8'h10 ;
			data[5503] <= 8'h10 ;
			data[5504] <= 8'h10 ;
			data[5505] <= 8'h10 ;
			data[5506] <= 8'h10 ;
			data[5507] <= 8'h10 ;
			data[5508] <= 8'h10 ;
			data[5509] <= 8'h10 ;
			data[5510] <= 8'h10 ;
			data[5511] <= 8'h10 ;
			data[5512] <= 8'h10 ;
			data[5513] <= 8'h10 ;
			data[5514] <= 8'h10 ;
			data[5515] <= 8'h10 ;
			data[5516] <= 8'h10 ;
			data[5517] <= 8'h10 ;
			data[5518] <= 8'h10 ;
			data[5519] <= 8'h10 ;
			data[5520] <= 8'h10 ;
			data[5521] <= 8'h10 ;
			data[5522] <= 8'h10 ;
			data[5523] <= 8'h10 ;
			data[5524] <= 8'h10 ;
			data[5525] <= 8'h10 ;
			data[5526] <= 8'h10 ;
			data[5527] <= 8'h10 ;
			data[5528] <= 8'h10 ;
			data[5529] <= 8'h10 ;
			data[5530] <= 8'h10 ;
			data[5531] <= 8'h10 ;
			data[5532] <= 8'h10 ;
			data[5533] <= 8'h10 ;
			data[5534] <= 8'h10 ;
			data[5535] <= 8'h10 ;
			data[5536] <= 8'h10 ;
			data[5537] <= 8'h10 ;
			data[5538] <= 8'h10 ;
			data[5539] <= 8'h10 ;
			data[5540] <= 8'h10 ;
			data[5541] <= 8'h10 ;
			data[5542] <= 8'h10 ;
			data[5543] <= 8'h10 ;
			data[5544] <= 8'h10 ;
			data[5545] <= 8'h10 ;
			data[5546] <= 8'h10 ;
			data[5547] <= 8'h10 ;
			data[5548] <= 8'h10 ;
			data[5549] <= 8'h10 ;
			data[5550] <= 8'h10 ;
			data[5551] <= 8'h10 ;
			data[5552] <= 8'h10 ;
			data[5553] <= 8'h10 ;
			data[5554] <= 8'h10 ;
			data[5555] <= 8'h10 ;
			data[5556] <= 8'h10 ;
			data[5557] <= 8'h10 ;
			data[5558] <= 8'h10 ;
			data[5559] <= 8'h10 ;
			data[5560] <= 8'h10 ;
			data[5561] <= 8'h10 ;
			data[5562] <= 8'h10 ;
			data[5563] <= 8'h10 ;
			data[5564] <= 8'h10 ;
			data[5565] <= 8'h10 ;
			data[5566] <= 8'h10 ;
			data[5567] <= 8'h10 ;
			data[5568] <= 8'h10 ;
			data[5569] <= 8'h10 ;
			data[5570] <= 8'h10 ;
			data[5571] <= 8'h10 ;
			data[5572] <= 8'h10 ;
			data[5573] <= 8'h10 ;
			data[5574] <= 8'h10 ;
			data[5575] <= 8'h10 ;
			data[5576] <= 8'h10 ;
			data[5577] <= 8'h10 ;
			data[5578] <= 8'h10 ;
			data[5579] <= 8'h10 ;
			data[5580] <= 8'h10 ;
			data[5581] <= 8'h10 ;
			data[5582] <= 8'h10 ;
			data[5583] <= 8'h10 ;
			data[5584] <= 8'h10 ;
			data[5585] <= 8'h10 ;
			data[5586] <= 8'h10 ;
			data[5587] <= 8'h10 ;
			data[5588] <= 8'h10 ;
			data[5589] <= 8'h10 ;
			data[5590] <= 8'h10 ;
			data[5591] <= 8'h10 ;
			data[5592] <= 8'h10 ;
			data[5593] <= 8'h10 ;
			data[5594] <= 8'h10 ;
			data[5595] <= 8'h10 ;
			data[5596] <= 8'h10 ;
			data[5597] <= 8'h10 ;
			data[5598] <= 8'h10 ;
			data[5599] <= 8'h10 ;
			data[5600] <= 8'h10 ;
			data[5601] <= 8'h10 ;
			data[5602] <= 8'h10 ;
			data[5603] <= 8'h10 ;
			data[5604] <= 8'h10 ;
			data[5605] <= 8'h10 ;
			data[5606] <= 8'h10 ;
			data[5607] <= 8'h10 ;
			data[5608] <= 8'h10 ;
			data[5609] <= 8'h10 ;
			data[5610] <= 8'h10 ;
			data[5611] <= 8'h10 ;
			data[5612] <= 8'h10 ;
			data[5613] <= 8'h10 ;
			data[5614] <= 8'h10 ;
			data[5615] <= 8'h10 ;
			data[5616] <= 8'h10 ;
			data[5617] <= 8'h10 ;
			data[5618] <= 8'h10 ;
			data[5619] <= 8'h10 ;
			data[5620] <= 8'h10 ;
			data[5621] <= 8'h10 ;
			data[5622] <= 8'h10 ;
			data[5623] <= 8'h10 ;
			data[5624] <= 8'h10 ;
			data[5625] <= 8'h10 ;
			data[5626] <= 8'h10 ;
			data[5627] <= 8'h10 ;
			data[5628] <= 8'h10 ;
			data[5629] <= 8'h10 ;
			data[5630] <= 8'h10 ;
			data[5631] <= 8'h10 ;
			data[5632] <= 8'h10 ;
			data[5633] <= 8'h10 ;
			data[5634] <= 8'h10 ;
			data[5635] <= 8'h10 ;
			data[5636] <= 8'h10 ;
			data[5637] <= 8'h10 ;
			data[5638] <= 8'h10 ;
			data[5639] <= 8'h10 ;
			data[5640] <= 8'h10 ;
			data[5641] <= 8'h10 ;
			data[5642] <= 8'h10 ;
			data[5643] <= 8'h10 ;
			data[5644] <= 8'h10 ;
			data[5645] <= 8'h10 ;
			data[5646] <= 8'h10 ;
			data[5647] <= 8'h10 ;
			data[5648] <= 8'h10 ;
			data[5649] <= 8'h10 ;
			data[5650] <= 8'h10 ;
			data[5651] <= 8'h10 ;
			data[5652] <= 8'h10 ;
			data[5653] <= 8'h10 ;
			data[5654] <= 8'h10 ;
			data[5655] <= 8'h10 ;
			data[5656] <= 8'h10 ;
			data[5657] <= 8'h10 ;
			data[5658] <= 8'h10 ;
			data[5659] <= 8'h10 ;
			data[5660] <= 8'h10 ;
			data[5661] <= 8'h10 ;
			data[5662] <= 8'h10 ;
			data[5663] <= 8'h10 ;
			data[5664] <= 8'h10 ;
			data[5665] <= 8'h10 ;
			data[5666] <= 8'h10 ;
			data[5667] <= 8'h10 ;
			data[5668] <= 8'h10 ;
			data[5669] <= 8'h10 ;
			data[5670] <= 8'h10 ;
			data[5671] <= 8'h10 ;
			data[5672] <= 8'h10 ;
			data[5673] <= 8'h10 ;
			data[5674] <= 8'h10 ;
			data[5675] <= 8'h10 ;
			data[5676] <= 8'h10 ;
			data[5677] <= 8'h10 ;
			data[5678] <= 8'h10 ;
			data[5679] <= 8'h10 ;
			data[5680] <= 8'h10 ;
			data[5681] <= 8'h10 ;
			data[5682] <= 8'h10 ;
			data[5683] <= 8'h10 ;
			data[5684] <= 8'h10 ;
			data[5685] <= 8'h10 ;
			data[5686] <= 8'h10 ;
			data[5687] <= 8'h10 ;
			data[5688] <= 8'h10 ;
			data[5689] <= 8'h10 ;
			data[5690] <= 8'h10 ;
			data[5691] <= 8'h10 ;
			data[5692] <= 8'h10 ;
			data[5693] <= 8'h10 ;
			data[5694] <= 8'h10 ;
			data[5695] <= 8'h10 ;
			data[5696] <= 8'h10 ;
			data[5697] <= 8'h10 ;
			data[5698] <= 8'h10 ;
			data[5699] <= 8'h10 ;
			data[5700] <= 8'h10 ;
			data[5701] <= 8'h10 ;
			data[5702] <= 8'h10 ;
			data[5703] <= 8'h10 ;
			data[5704] <= 8'h10 ;
			data[5705] <= 8'h10 ;
			data[5706] <= 8'h10 ;
			data[5707] <= 8'h10 ;
			data[5708] <= 8'h10 ;
			data[5709] <= 8'h10 ;
			data[5710] <= 8'h10 ;
			data[5711] <= 8'h10 ;
			data[5712] <= 8'h10 ;
			data[5713] <= 8'h10 ;
			data[5714] <= 8'h10 ;
			data[5715] <= 8'h10 ;
			data[5716] <= 8'h10 ;
			data[5717] <= 8'h10 ;
			data[5718] <= 8'h10 ;
			data[5719] <= 8'h10 ;
			data[5720] <= 8'h10 ;
			data[5721] <= 8'h10 ;
			data[5722] <= 8'h10 ;
			data[5723] <= 8'h10 ;
			data[5724] <= 8'h10 ;
			data[5725] <= 8'h10 ;
			data[5726] <= 8'h10 ;
			data[5727] <= 8'h10 ;
			data[5728] <= 8'h10 ;
			data[5729] <= 8'h10 ;
			data[5730] <= 8'h10 ;
			data[5731] <= 8'h10 ;
			data[5732] <= 8'h10 ;
			data[5733] <= 8'h10 ;
			data[5734] <= 8'h10 ;
			data[5735] <= 8'h10 ;
			data[5736] <= 8'h10 ;
			data[5737] <= 8'h10 ;
			data[5738] <= 8'h10 ;
			data[5739] <= 8'h10 ;
			data[5740] <= 8'h10 ;
			data[5741] <= 8'h10 ;
			data[5742] <= 8'h10 ;
			data[5743] <= 8'h10 ;
			data[5744] <= 8'h10 ;
			data[5745] <= 8'h10 ;
			data[5746] <= 8'h10 ;
			data[5747] <= 8'h10 ;
			data[5748] <= 8'h10 ;
			data[5749] <= 8'h10 ;
			data[5750] <= 8'h10 ;
			data[5751] <= 8'h10 ;
			data[5752] <= 8'h10 ;
			data[5753] <= 8'h10 ;
			data[5754] <= 8'h10 ;
			data[5755] <= 8'h10 ;
			data[5756] <= 8'h10 ;
			data[5757] <= 8'h10 ;
			data[5758] <= 8'h10 ;
			data[5759] <= 8'h10 ;
			data[5760] <= 8'h10 ;
			data[5761] <= 8'h10 ;
			data[5762] <= 8'h10 ;
			data[5763] <= 8'h10 ;
			data[5764] <= 8'h10 ;
			data[5765] <= 8'h10 ;
			data[5766] <= 8'h10 ;
			data[5767] <= 8'h10 ;
			data[5768] <= 8'h10 ;
			data[5769] <= 8'h10 ;
			data[5770] <= 8'h10 ;
			data[5771] <= 8'h10 ;
			data[5772] <= 8'h10 ;
			data[5773] <= 8'h10 ;
			data[5774] <= 8'h10 ;
			data[5775] <= 8'h10 ;
			data[5776] <= 8'h10 ;
			data[5777] <= 8'h10 ;
			data[5778] <= 8'h10 ;
			data[5779] <= 8'h10 ;
			data[5780] <= 8'h10 ;
			data[5781] <= 8'h10 ;
			data[5782] <= 8'h10 ;
			data[5783] <= 8'h10 ;
			data[5784] <= 8'h10 ;
			data[5785] <= 8'h10 ;
			data[5786] <= 8'h10 ;
			data[5787] <= 8'h10 ;
			data[5788] <= 8'h10 ;
			data[5789] <= 8'h10 ;
			data[5790] <= 8'h10 ;
			data[5791] <= 8'h10 ;
			data[5792] <= 8'h10 ;
			data[5793] <= 8'h10 ;
			data[5794] <= 8'h10 ;
			data[5795] <= 8'h10 ;
			data[5796] <= 8'h10 ;
			data[5797] <= 8'h10 ;
			data[5798] <= 8'h10 ;
			data[5799] <= 8'h10 ;
			data[5800] <= 8'h10 ;
			data[5801] <= 8'h10 ;
			data[5802] <= 8'h10 ;
			data[5803] <= 8'h10 ;
			data[5804] <= 8'h10 ;
			data[5805] <= 8'h10 ;
			data[5806] <= 8'h10 ;
			data[5807] <= 8'h10 ;
			data[5808] <= 8'h10 ;
			data[5809] <= 8'h10 ;
			data[5810] <= 8'h10 ;
			data[5811] <= 8'h10 ;
			data[5812] <= 8'h10 ;
			data[5813] <= 8'h10 ;
			data[5814] <= 8'h10 ;
			data[5815] <= 8'h10 ;
			data[5816] <= 8'h10 ;
			data[5817] <= 8'h10 ;
			data[5818] <= 8'h10 ;
			data[5819] <= 8'h10 ;
			data[5820] <= 8'h10 ;
			data[5821] <= 8'h10 ;
			data[5822] <= 8'h10 ;
			data[5823] <= 8'h10 ;
			data[5824] <= 8'h10 ;
			data[5825] <= 8'h10 ;
			data[5826] <= 8'h10 ;
			data[5827] <= 8'h10 ;
			data[5828] <= 8'h10 ;
			data[5829] <= 8'h10 ;
			data[5830] <= 8'h10 ;
			data[5831] <= 8'h10 ;
			data[5832] <= 8'h10 ;
			data[5833] <= 8'h10 ;
			data[5834] <= 8'h10 ;
			data[5835] <= 8'h10 ;
			data[5836] <= 8'h10 ;
			data[5837] <= 8'h10 ;
			data[5838] <= 8'h10 ;
			data[5839] <= 8'h10 ;
			data[5840] <= 8'h10 ;
			data[5841] <= 8'h10 ;
			data[5842] <= 8'h10 ;
			data[5843] <= 8'h10 ;
			data[5844] <= 8'h10 ;
			data[5845] <= 8'h10 ;
			data[5846] <= 8'h10 ;
			data[5847] <= 8'h10 ;
			data[5848] <= 8'h10 ;
			data[5849] <= 8'h10 ;
			data[5850] <= 8'h10 ;
			data[5851] <= 8'h10 ;
			data[5852] <= 8'h10 ;
			data[5853] <= 8'h10 ;
			data[5854] <= 8'h10 ;
			data[5855] <= 8'h10 ;
			data[5856] <= 8'h10 ;
			data[5857] <= 8'h10 ;
			data[5858] <= 8'h10 ;
			data[5859] <= 8'h10 ;
			data[5860] <= 8'h10 ;
			data[5861] <= 8'h10 ;
			data[5862] <= 8'h10 ;
			data[5863] <= 8'h10 ;
			data[5864] <= 8'h10 ;
			data[5865] <= 8'h10 ;
			data[5866] <= 8'h10 ;
			data[5867] <= 8'h10 ;
			data[5868] <= 8'h10 ;
			data[5869] <= 8'h10 ;
			data[5870] <= 8'h10 ;
			data[5871] <= 8'h10 ;
			data[5872] <= 8'h10 ;
			data[5873] <= 8'h10 ;
			data[5874] <= 8'h10 ;
			data[5875] <= 8'h10 ;
			data[5876] <= 8'h10 ;
			data[5877] <= 8'h10 ;
			data[5878] <= 8'h10 ;
			data[5879] <= 8'h10 ;
			data[5880] <= 8'h10 ;
			data[5881] <= 8'h10 ;
			data[5882] <= 8'h10 ;
			data[5883] <= 8'h10 ;
			data[5884] <= 8'h10 ;
			data[5885] <= 8'h10 ;
			data[5886] <= 8'h10 ;
			data[5887] <= 8'h10 ;
			data[5888] <= 8'h10 ;
			data[5889] <= 8'h10 ;
			data[5890] <= 8'h10 ;
			data[5891] <= 8'h10 ;
			data[5892] <= 8'h10 ;
			data[5893] <= 8'h10 ;
			data[5894] <= 8'h10 ;
			data[5895] <= 8'h10 ;
			data[5896] <= 8'h10 ;
			data[5897] <= 8'h10 ;
			data[5898] <= 8'h10 ;
			data[5899] <= 8'h10 ;
			data[5900] <= 8'h10 ;
			data[5901] <= 8'h10 ;
			data[5902] <= 8'h10 ;
			data[5903] <= 8'h10 ;
			data[5904] <= 8'h10 ;
			data[5905] <= 8'h10 ;
			data[5906] <= 8'h10 ;
			data[5907] <= 8'h10 ;
			data[5908] <= 8'h10 ;
			data[5909] <= 8'h10 ;
			data[5910] <= 8'h10 ;
			data[5911] <= 8'h10 ;
			data[5912] <= 8'h10 ;
			data[5913] <= 8'h10 ;
			data[5914] <= 8'h10 ;
			data[5915] <= 8'h10 ;
			data[5916] <= 8'h10 ;
			data[5917] <= 8'h10 ;
			data[5918] <= 8'h10 ;
			data[5919] <= 8'h10 ;
			data[5920] <= 8'h10 ;
			data[5921] <= 8'h10 ;
			data[5922] <= 8'h10 ;
			data[5923] <= 8'h10 ;
			data[5924] <= 8'h10 ;
			data[5925] <= 8'h10 ;
			data[5926] <= 8'h10 ;
			data[5927] <= 8'h10 ;
			data[5928] <= 8'h10 ;
			data[5929] <= 8'h10 ;
			data[5930] <= 8'h10 ;
			data[5931] <= 8'h10 ;
			data[5932] <= 8'h10 ;
			data[5933] <= 8'h10 ;
			data[5934] <= 8'h10 ;
			data[5935] <= 8'h10 ;
			data[5936] <= 8'h10 ;
			data[5937] <= 8'h10 ;
			data[5938] <= 8'h10 ;
			data[5939] <= 8'h10 ;
			data[5940] <= 8'h10 ;
			data[5941] <= 8'h10 ;
			data[5942] <= 8'h10 ;
			data[5943] <= 8'h10 ;
			data[5944] <= 8'h10 ;
			data[5945] <= 8'h10 ;
			data[5946] <= 8'h10 ;
			data[5947] <= 8'h10 ;
			data[5948] <= 8'h10 ;
			data[5949] <= 8'h10 ;
			data[5950] <= 8'h10 ;
			data[5951] <= 8'h10 ;
			data[5952] <= 8'h10 ;
			data[5953] <= 8'h10 ;
			data[5954] <= 8'h10 ;
			data[5955] <= 8'h10 ;
			data[5956] <= 8'h10 ;
			data[5957] <= 8'h10 ;
			data[5958] <= 8'h10 ;
			data[5959] <= 8'h10 ;
			data[5960] <= 8'h10 ;
			data[5961] <= 8'h10 ;
			data[5962] <= 8'h10 ;
			data[5963] <= 8'h10 ;
			data[5964] <= 8'h10 ;
			data[5965] <= 8'h10 ;
			data[5966] <= 8'h10 ;
			data[5967] <= 8'h10 ;
			data[5968] <= 8'h10 ;
			data[5969] <= 8'h10 ;
			data[5970] <= 8'h10 ;
			data[5971] <= 8'h10 ;
			data[5972] <= 8'h10 ;
			data[5973] <= 8'h10 ;
			data[5974] <= 8'h10 ;
			data[5975] <= 8'h10 ;
			data[5976] <= 8'h10 ;
			data[5977] <= 8'h10 ;
			data[5978] <= 8'h10 ;
			data[5979] <= 8'h10 ;
			data[5980] <= 8'h10 ;
			data[5981] <= 8'h10 ;
			data[5982] <= 8'h10 ;
			data[5983] <= 8'h10 ;
			data[5984] <= 8'h10 ;
			data[5985] <= 8'h10 ;
			data[5986] <= 8'h10 ;
			data[5987] <= 8'h10 ;
			data[5988] <= 8'h10 ;
			data[5989] <= 8'h10 ;
			data[5990] <= 8'h10 ;
			data[5991] <= 8'h10 ;
			data[5992] <= 8'h10 ;
			data[5993] <= 8'h10 ;
			data[5994] <= 8'h10 ;
			data[5995] <= 8'h10 ;
			data[5996] <= 8'h10 ;
			data[5997] <= 8'h10 ;
			data[5998] <= 8'h10 ;
			data[5999] <= 8'h10 ;
			data[6000] <= 8'h10 ;
			data[6001] <= 8'h10 ;
			data[6002] <= 8'h10 ;
			data[6003] <= 8'h10 ;
			data[6004] <= 8'h10 ;
			data[6005] <= 8'h10 ;
			data[6006] <= 8'h10 ;
			data[6007] <= 8'h10 ;
			data[6008] <= 8'h10 ;
			data[6009] <= 8'h10 ;
			data[6010] <= 8'h10 ;
			data[6011] <= 8'h10 ;
			data[6012] <= 8'h10 ;
			data[6013] <= 8'h10 ;
			data[6014] <= 8'h10 ;
			data[6015] <= 8'h10 ;
			data[6016] <= 8'h10 ;
			data[6017] <= 8'h10 ;
			data[6018] <= 8'h10 ;
			data[6019] <= 8'h10 ;
			data[6020] <= 8'h10 ;
			data[6021] <= 8'h10 ;
			data[6022] <= 8'h10 ;
			data[6023] <= 8'h10 ;
			data[6024] <= 8'h10 ;
			data[6025] <= 8'h10 ;
			data[6026] <= 8'h10 ;
			data[6027] <= 8'h10 ;
			data[6028] <= 8'h10 ;
			data[6029] <= 8'h10 ;
			data[6030] <= 8'h10 ;
			data[6031] <= 8'h10 ;
			data[6032] <= 8'h10 ;
			data[6033] <= 8'h10 ;
			data[6034] <= 8'h10 ;
			data[6035] <= 8'h10 ;
			data[6036] <= 8'h10 ;
			data[6037] <= 8'h10 ;
			data[6038] <= 8'h10 ;
			data[6039] <= 8'h10 ;
			data[6040] <= 8'h10 ;
			data[6041] <= 8'h10 ;
			data[6042] <= 8'h10 ;
			data[6043] <= 8'h10 ;
			data[6044] <= 8'h10 ;
			data[6045] <= 8'h10 ;
			data[6046] <= 8'h10 ;
			data[6047] <= 8'h10 ;
			data[6048] <= 8'h10 ;
			data[6049] <= 8'h10 ;
			data[6050] <= 8'h10 ;
			data[6051] <= 8'h10 ;
			data[6052] <= 8'h10 ;
			data[6053] <= 8'h10 ;
			data[6054] <= 8'h10 ;
			data[6055] <= 8'h10 ;
			data[6056] <= 8'h10 ;
			data[6057] <= 8'h10 ;
			data[6058] <= 8'h10 ;
			data[6059] <= 8'h10 ;
			data[6060] <= 8'h10 ;
			data[6061] <= 8'h10 ;
			data[6062] <= 8'h10 ;
			data[6063] <= 8'h10 ;
			data[6064] <= 8'h10 ;
			data[6065] <= 8'h10 ;
			data[6066] <= 8'h10 ;
			data[6067] <= 8'h10 ;
			data[6068] <= 8'h10 ;
			data[6069] <= 8'h10 ;
			data[6070] <= 8'h10 ;
			data[6071] <= 8'h10 ;
			data[6072] <= 8'h10 ;
			data[6073] <= 8'h10 ;
			data[6074] <= 8'h10 ;
			data[6075] <= 8'h10 ;
			data[6076] <= 8'h10 ;
			data[6077] <= 8'h10 ;
			data[6078] <= 8'h10 ;
			data[6079] <= 8'h10 ;
			data[6080] <= 8'h10 ;
			data[6081] <= 8'h10 ;
			data[6082] <= 8'h10 ;
			data[6083] <= 8'h10 ;
			data[6084] <= 8'h10 ;
			data[6085] <= 8'h10 ;
			data[6086] <= 8'h10 ;
			data[6087] <= 8'h10 ;
			data[6088] <= 8'h10 ;
			data[6089] <= 8'h10 ;
			data[6090] <= 8'h10 ;
			data[6091] <= 8'h10 ;
			data[6092] <= 8'h10 ;
			data[6093] <= 8'h10 ;
			data[6094] <= 8'h10 ;
			data[6095] <= 8'h10 ;
			data[6096] <= 8'h10 ;
			data[6097] <= 8'h10 ;
			data[6098] <= 8'h10 ;
			data[6099] <= 8'h10 ;
			data[6100] <= 8'h10 ;
			data[6101] <= 8'h10 ;
			data[6102] <= 8'h10 ;
			data[6103] <= 8'h10 ;
			data[6104] <= 8'h10 ;
			data[6105] <= 8'h10 ;
			data[6106] <= 8'h10 ;
			data[6107] <= 8'h10 ;
			data[6108] <= 8'h10 ;
			data[6109] <= 8'h10 ;
			data[6110] <= 8'h10 ;
			data[6111] <= 8'h10 ;
			data[6112] <= 8'h10 ;
			data[6113] <= 8'h10 ;
			data[6114] <= 8'h10 ;
			data[6115] <= 8'h10 ;
			data[6116] <= 8'h10 ;
			data[6117] <= 8'h10 ;
			data[6118] <= 8'h10 ;
			data[6119] <= 8'h10 ;
			data[6120] <= 8'h10 ;
			data[6121] <= 8'h10 ;
			data[6122] <= 8'h10 ;
			data[6123] <= 8'h10 ;
			data[6124] <= 8'h10 ;
			data[6125] <= 8'h10 ;
			data[6126] <= 8'h10 ;
			data[6127] <= 8'h10 ;
			data[6128] <= 8'h10 ;
			data[6129] <= 8'h10 ;
			data[6130] <= 8'h10 ;
			data[6131] <= 8'h10 ;
			data[6132] <= 8'h10 ;
			data[6133] <= 8'h10 ;
			data[6134] <= 8'h10 ;
			data[6135] <= 8'h10 ;
			data[6136] <= 8'h10 ;
			data[6137] <= 8'h10 ;
			data[6138] <= 8'h10 ;
			data[6139] <= 8'h10 ;
			data[6140] <= 8'h10 ;
			data[6141] <= 8'h10 ;
			data[6142] <= 8'h10 ;
			data[6143] <= 8'h10 ;
			data[6144] <= 8'h10 ;
			data[6145] <= 8'h10 ;
			data[6146] <= 8'h10 ;
			data[6147] <= 8'h10 ;
			data[6148] <= 8'h10 ;
			data[6149] <= 8'h10 ;
			data[6150] <= 8'h10 ;
			data[6151] <= 8'h10 ;
			data[6152] <= 8'h10 ;
			data[6153] <= 8'h10 ;
			data[6154] <= 8'h10 ;
			data[6155] <= 8'h10 ;
			data[6156] <= 8'h10 ;
			data[6157] <= 8'h10 ;
			data[6158] <= 8'h10 ;
			data[6159] <= 8'h10 ;
			data[6160] <= 8'h10 ;
			data[6161] <= 8'h10 ;
			data[6162] <= 8'h10 ;
			data[6163] <= 8'h10 ;
			data[6164] <= 8'h10 ;
			data[6165] <= 8'h10 ;
			data[6166] <= 8'h10 ;
			data[6167] <= 8'h10 ;
			data[6168] <= 8'h10 ;
			data[6169] <= 8'h10 ;
			data[6170] <= 8'h10 ;
			data[6171] <= 8'h10 ;
			data[6172] <= 8'h10 ;
			data[6173] <= 8'h10 ;
			data[6174] <= 8'h10 ;
			data[6175] <= 8'h10 ;
			data[6176] <= 8'h10 ;
			data[6177] <= 8'h10 ;
			data[6178] <= 8'h10 ;
			data[6179] <= 8'h10 ;
			data[6180] <= 8'h10 ;
			data[6181] <= 8'h10 ;
			data[6182] <= 8'h10 ;
			data[6183] <= 8'h10 ;
			data[6184] <= 8'h10 ;
			data[6185] <= 8'h10 ;
			data[6186] <= 8'h10 ;
			data[6187] <= 8'h10 ;
			data[6188] <= 8'h10 ;
			data[6189] <= 8'h10 ;
			data[6190] <= 8'h10 ;
			data[6191] <= 8'h10 ;
			data[6192] <= 8'h10 ;
			data[6193] <= 8'h10 ;
			data[6194] <= 8'h10 ;
			data[6195] <= 8'h10 ;
			data[6196] <= 8'h10 ;
			data[6197] <= 8'h10 ;
			data[6198] <= 8'h10 ;
			data[6199] <= 8'h10 ;
			data[6200] <= 8'h10 ;
			data[6201] <= 8'h10 ;
			data[6202] <= 8'h10 ;
			data[6203] <= 8'h10 ;
			data[6204] <= 8'h10 ;
			data[6205] <= 8'h10 ;
			data[6206] <= 8'h10 ;
			data[6207] <= 8'h10 ;
			data[6208] <= 8'h10 ;
			data[6209] <= 8'h10 ;
			data[6210] <= 8'h10 ;
			data[6211] <= 8'h10 ;
			data[6212] <= 8'h10 ;
			data[6213] <= 8'h10 ;
			data[6214] <= 8'h10 ;
			data[6215] <= 8'h10 ;
			data[6216] <= 8'h10 ;
			data[6217] <= 8'h10 ;
			data[6218] <= 8'h10 ;
			data[6219] <= 8'h10 ;
			data[6220] <= 8'h10 ;
			data[6221] <= 8'h10 ;
			data[6222] <= 8'h10 ;
			data[6223] <= 8'h10 ;
			data[6224] <= 8'h10 ;
			data[6225] <= 8'h10 ;
			data[6226] <= 8'h10 ;
			data[6227] <= 8'h10 ;
			data[6228] <= 8'h10 ;
			data[6229] <= 8'h10 ;
			data[6230] <= 8'h10 ;
			data[6231] <= 8'h10 ;
			data[6232] <= 8'h10 ;
			data[6233] <= 8'h10 ;
			data[6234] <= 8'h10 ;
			data[6235] <= 8'h10 ;
			data[6236] <= 8'h10 ;
			data[6237] <= 8'h10 ;
			data[6238] <= 8'h10 ;
			data[6239] <= 8'h10 ;
			data[6240] <= 8'h10 ;
			data[6241] <= 8'h10 ;
			data[6242] <= 8'h10 ;
			data[6243] <= 8'h10 ;
			data[6244] <= 8'h10 ;
			data[6245] <= 8'h10 ;
			data[6246] <= 8'h10 ;
			data[6247] <= 8'h10 ;
			data[6248] <= 8'h10 ;
			data[6249] <= 8'h10 ;
			data[6250] <= 8'h10 ;
			data[6251] <= 8'h10 ;
			data[6252] <= 8'h10 ;
			data[6253] <= 8'h10 ;
			data[6254] <= 8'h10 ;
			data[6255] <= 8'h10 ;
			data[6256] <= 8'h10 ;
			data[6257] <= 8'h10 ;
			data[6258] <= 8'h10 ;
			data[6259] <= 8'h10 ;
			data[6260] <= 8'h10 ;
			data[6261] <= 8'h10 ;
			data[6262] <= 8'h10 ;
			data[6263] <= 8'h10 ;
			data[6264] <= 8'h10 ;
			data[6265] <= 8'h10 ;
			data[6266] <= 8'h10 ;
			data[6267] <= 8'h10 ;
			data[6268] <= 8'h10 ;
			data[6269] <= 8'h10 ;
			data[6270] <= 8'h10 ;
			data[6271] <= 8'h10 ;
			data[6272] <= 8'h10 ;
			data[6273] <= 8'h10 ;
			data[6274] <= 8'h10 ;
			data[6275] <= 8'h10 ;
			data[6276] <= 8'h10 ;
			data[6277] <= 8'h10 ;
			data[6278] <= 8'h10 ;
			data[6279] <= 8'h10 ;
			data[6280] <= 8'h10 ;
			data[6281] <= 8'h10 ;
			data[6282] <= 8'h10 ;
			data[6283] <= 8'h10 ;
			data[6284] <= 8'h10 ;
			data[6285] <= 8'h10 ;
			data[6286] <= 8'h10 ;
			data[6287] <= 8'h10 ;
			data[6288] <= 8'h10 ;
			data[6289] <= 8'h10 ;
			data[6290] <= 8'h10 ;
			data[6291] <= 8'h10 ;
			data[6292] <= 8'h10 ;
			data[6293] <= 8'h10 ;
			data[6294] <= 8'h10 ;
			data[6295] <= 8'h10 ;
			data[6296] <= 8'h10 ;
			data[6297] <= 8'h10 ;
			data[6298] <= 8'h10 ;
			data[6299] <= 8'h10 ;
			data[6300] <= 8'h10 ;
			data[6301] <= 8'h10 ;
			data[6302] <= 8'h10 ;
			data[6303] <= 8'h10 ;
			data[6304] <= 8'h10 ;
			data[6305] <= 8'h10 ;
			data[6306] <= 8'h10 ;
			data[6307] <= 8'h10 ;
			data[6308] <= 8'h10 ;
			data[6309] <= 8'h10 ;
			data[6310] <= 8'h10 ;
			data[6311] <= 8'h10 ;
			data[6312] <= 8'h10 ;
			data[6313] <= 8'h10 ;
			data[6314] <= 8'h10 ;
			data[6315] <= 8'h10 ;
			data[6316] <= 8'h10 ;
			data[6317] <= 8'h10 ;
			data[6318] <= 8'h10 ;
			data[6319] <= 8'h10 ;
			data[6320] <= 8'h10 ;
			data[6321] <= 8'h10 ;
			data[6322] <= 8'h10 ;
			data[6323] <= 8'h10 ;
			data[6324] <= 8'h10 ;
			data[6325] <= 8'h10 ;
			data[6326] <= 8'h10 ;
			data[6327] <= 8'h10 ;
			data[6328] <= 8'h10 ;
			data[6329] <= 8'h10 ;
			data[6330] <= 8'h10 ;
			data[6331] <= 8'h10 ;
			data[6332] <= 8'h10 ;
			data[6333] <= 8'h10 ;
			data[6334] <= 8'h10 ;
			data[6335] <= 8'h10 ;
			data[6336] <= 8'h10 ;
			data[6337] <= 8'h10 ;
			data[6338] <= 8'h10 ;
			data[6339] <= 8'h10 ;
			data[6340] <= 8'h10 ;
			data[6341] <= 8'h10 ;
			data[6342] <= 8'h10 ;
			data[6343] <= 8'h10 ;
			data[6344] <= 8'h10 ;
			data[6345] <= 8'h10 ;
			data[6346] <= 8'h10 ;
			data[6347] <= 8'h10 ;
			data[6348] <= 8'h10 ;
			data[6349] <= 8'h10 ;
			data[6350] <= 8'h10 ;
			data[6351] <= 8'h10 ;
			data[6352] <= 8'h10 ;
			data[6353] <= 8'h10 ;
			data[6354] <= 8'h10 ;
			data[6355] <= 8'h10 ;
			data[6356] <= 8'h10 ;
			data[6357] <= 8'h10 ;
			data[6358] <= 8'h10 ;
			data[6359] <= 8'h10 ;
			data[6360] <= 8'h10 ;
			data[6361] <= 8'h10 ;
			data[6362] <= 8'h10 ;
			data[6363] <= 8'h10 ;
			data[6364] <= 8'h10 ;
			data[6365] <= 8'h10 ;
			data[6366] <= 8'h10 ;
			data[6367] <= 8'h10 ;
			data[6368] <= 8'h10 ;
			data[6369] <= 8'h10 ;
			data[6370] <= 8'h10 ;
			data[6371] <= 8'h10 ;
			data[6372] <= 8'h10 ;
			data[6373] <= 8'h10 ;
			data[6374] <= 8'h10 ;
			data[6375] <= 8'h10 ;
			data[6376] <= 8'h10 ;
			data[6377] <= 8'h10 ;
			data[6378] <= 8'h10 ;
			data[6379] <= 8'h10 ;
			data[6380] <= 8'h10 ;
			data[6381] <= 8'h10 ;
			data[6382] <= 8'h10 ;
			data[6383] <= 8'h10 ;
			data[6384] <= 8'h10 ;
			data[6385] <= 8'h10 ;
			data[6386] <= 8'h10 ;
			data[6387] <= 8'h10 ;
			data[6388] <= 8'h10 ;
			data[6389] <= 8'h10 ;
			data[6390] <= 8'h10 ;
			data[6391] <= 8'h10 ;
			data[6392] <= 8'h10 ;
			data[6393] <= 8'h10 ;
			data[6394] <= 8'h10 ;
			data[6395] <= 8'h10 ;
			data[6396] <= 8'h10 ;
			data[6397] <= 8'h10 ;
			data[6398] <= 8'h10 ;
			data[6399] <= 8'h10 ;
			data[6400] <= 8'h10 ;
			data[6401] <= 8'h10 ;
			data[6402] <= 8'h10 ;
			data[6403] <= 8'h10 ;
			data[6404] <= 8'h10 ;
			data[6405] <= 8'h10 ;
			data[6406] <= 8'h10 ;
			data[6407] <= 8'h10 ;
			data[6408] <= 8'h10 ;
			data[6409] <= 8'h10 ;
			data[6410] <= 8'h10 ;
			data[6411] <= 8'h10 ;
			data[6412] <= 8'h10 ;
			data[6413] <= 8'h10 ;
			data[6414] <= 8'h10 ;
			data[6415] <= 8'h10 ;
			data[6416] <= 8'h10 ;
			data[6417] <= 8'h10 ;
			data[6418] <= 8'h10 ;
			data[6419] <= 8'h10 ;
			data[6420] <= 8'h10 ;
			data[6421] <= 8'h10 ;
			data[6422] <= 8'h10 ;
			data[6423] <= 8'h10 ;
			data[6424] <= 8'h10 ;
			data[6425] <= 8'h10 ;
			data[6426] <= 8'h10 ;
			data[6427] <= 8'h10 ;
			data[6428] <= 8'h10 ;
			data[6429] <= 8'h10 ;
			data[6430] <= 8'h10 ;
			data[6431] <= 8'h10 ;
			data[6432] <= 8'h10 ;
			data[6433] <= 8'h10 ;
			data[6434] <= 8'h10 ;
			data[6435] <= 8'h10 ;
			data[6436] <= 8'h10 ;
			data[6437] <= 8'h10 ;
			data[6438] <= 8'h10 ;
			data[6439] <= 8'h10 ;
			data[6440] <= 8'h10 ;
			data[6441] <= 8'h10 ;
			data[6442] <= 8'h10 ;
			data[6443] <= 8'h10 ;
			data[6444] <= 8'h10 ;
			data[6445] <= 8'h10 ;
			data[6446] <= 8'h10 ;
			data[6447] <= 8'h10 ;
			data[6448] <= 8'h10 ;
			data[6449] <= 8'h10 ;
			data[6450] <= 8'h10 ;
			data[6451] <= 8'h10 ;
			data[6452] <= 8'h10 ;
			data[6453] <= 8'h10 ;
			data[6454] <= 8'h10 ;
			data[6455] <= 8'h10 ;
			data[6456] <= 8'h10 ;
			data[6457] <= 8'h10 ;
			data[6458] <= 8'h10 ;
			data[6459] <= 8'h10 ;
			data[6460] <= 8'h10 ;
			data[6461] <= 8'h10 ;
			data[6462] <= 8'h10 ;
			data[6463] <= 8'h10 ;
			data[6464] <= 8'h10 ;
			data[6465] <= 8'h10 ;
			data[6466] <= 8'h10 ;
			data[6467] <= 8'h10 ;
			data[6468] <= 8'h10 ;
			data[6469] <= 8'h10 ;
			data[6470] <= 8'h10 ;
			data[6471] <= 8'h10 ;
			data[6472] <= 8'h10 ;
			data[6473] <= 8'h10 ;
			data[6474] <= 8'h10 ;
			data[6475] <= 8'h10 ;
			data[6476] <= 8'h10 ;
			data[6477] <= 8'h10 ;
			data[6478] <= 8'h10 ;
			data[6479] <= 8'h10 ;
			data[6480] <= 8'h10 ;
			data[6481] <= 8'h10 ;
			data[6482] <= 8'h10 ;
			data[6483] <= 8'h10 ;
			data[6484] <= 8'h10 ;
			data[6485] <= 8'h10 ;
			data[6486] <= 8'h10 ;
			data[6487] <= 8'h10 ;
			data[6488] <= 8'h10 ;
			data[6489] <= 8'h10 ;
			data[6490] <= 8'h10 ;
			data[6491] <= 8'h10 ;
			data[6492] <= 8'h10 ;
			data[6493] <= 8'h10 ;
			data[6494] <= 8'h10 ;
			data[6495] <= 8'h10 ;
			data[6496] <= 8'h10 ;
			data[6497] <= 8'h10 ;
			data[6498] <= 8'h10 ;
			data[6499] <= 8'h10 ;
			data[6500] <= 8'h10 ;
			data[6501] <= 8'h10 ;
			data[6502] <= 8'h10 ;
			data[6503] <= 8'h10 ;
			data[6504] <= 8'h10 ;
			data[6505] <= 8'h10 ;
			data[6506] <= 8'h10 ;
			data[6507] <= 8'h10 ;
			data[6508] <= 8'h10 ;
			data[6509] <= 8'h10 ;
			data[6510] <= 8'h10 ;
			data[6511] <= 8'h10 ;
			data[6512] <= 8'h10 ;
			data[6513] <= 8'h10 ;
			data[6514] <= 8'h10 ;
			data[6515] <= 8'h10 ;
			data[6516] <= 8'h10 ;
			data[6517] <= 8'h10 ;
			data[6518] <= 8'h10 ;
			data[6519] <= 8'h10 ;
			data[6520] <= 8'h10 ;
			data[6521] <= 8'h10 ;
			data[6522] <= 8'h10 ;
			data[6523] <= 8'h10 ;
			data[6524] <= 8'h10 ;
			data[6525] <= 8'h10 ;
			data[6526] <= 8'h10 ;
			data[6527] <= 8'h10 ;
			data[6528] <= 8'h10 ;
			data[6529] <= 8'h10 ;
			data[6530] <= 8'h10 ;
			data[6531] <= 8'h10 ;
			data[6532] <= 8'h10 ;
			data[6533] <= 8'h10 ;
			data[6534] <= 8'h10 ;
			data[6535] <= 8'h10 ;
			data[6536] <= 8'h10 ;
			data[6537] <= 8'h10 ;
			data[6538] <= 8'h10 ;
			data[6539] <= 8'h10 ;
			data[6540] <= 8'h10 ;
			data[6541] <= 8'h10 ;
			data[6542] <= 8'h10 ;
			data[6543] <= 8'h10 ;
			data[6544] <= 8'h10 ;
			data[6545] <= 8'h10 ;
			data[6546] <= 8'h10 ;
			data[6547] <= 8'h10 ;
			data[6548] <= 8'h10 ;
			data[6549] <= 8'h10 ;
			data[6550] <= 8'h10 ;
			data[6551] <= 8'h10 ;
			data[6552] <= 8'h10 ;
			data[6553] <= 8'h10 ;
			data[6554] <= 8'h10 ;
			data[6555] <= 8'h10 ;
			data[6556] <= 8'h10 ;
			data[6557] <= 8'h10 ;
			data[6558] <= 8'h10 ;
			data[6559] <= 8'h10 ;
			data[6560] <= 8'h10 ;
			data[6561] <= 8'h10 ;
			data[6562] <= 8'h10 ;
			data[6563] <= 8'h10 ;
			data[6564] <= 8'h10 ;
			data[6565] <= 8'h10 ;
			data[6566] <= 8'h10 ;
			data[6567] <= 8'h10 ;
			data[6568] <= 8'h10 ;
			data[6569] <= 8'h10 ;
			data[6570] <= 8'h10 ;
			data[6571] <= 8'h10 ;
			data[6572] <= 8'h10 ;
			data[6573] <= 8'h10 ;
			data[6574] <= 8'h10 ;
			data[6575] <= 8'h10 ;
			data[6576] <= 8'h10 ;
			data[6577] <= 8'h10 ;
			data[6578] <= 8'h10 ;
			data[6579] <= 8'h10 ;
			data[6580] <= 8'h10 ;
			data[6581] <= 8'h10 ;
			data[6582] <= 8'h10 ;
			data[6583] <= 8'h10 ;
			data[6584] <= 8'h10 ;
			data[6585] <= 8'h10 ;
			data[6586] <= 8'h10 ;
			data[6587] <= 8'h10 ;
			data[6588] <= 8'h10 ;
			data[6589] <= 8'h10 ;
			data[6590] <= 8'h10 ;
			data[6591] <= 8'h10 ;
			data[6592] <= 8'h10 ;
			data[6593] <= 8'h10 ;
			data[6594] <= 8'h10 ;
			data[6595] <= 8'h10 ;
			data[6596] <= 8'h10 ;
			data[6597] <= 8'h10 ;
			data[6598] <= 8'h10 ;
			data[6599] <= 8'h10 ;
			data[6600] <= 8'h10 ;
			data[6601] <= 8'h10 ;
			data[6602] <= 8'h10 ;
			data[6603] <= 8'h10 ;
			data[6604] <= 8'h10 ;
			data[6605] <= 8'h10 ;
			data[6606] <= 8'h10 ;
			data[6607] <= 8'h10 ;
			data[6608] <= 8'h10 ;
			data[6609] <= 8'h10 ;
			data[6610] <= 8'h10 ;
			data[6611] <= 8'h10 ;
			data[6612] <= 8'h10 ;
			data[6613] <= 8'h10 ;
			data[6614] <= 8'h10 ;
			data[6615] <= 8'h10 ;
			data[6616] <= 8'h10 ;
			data[6617] <= 8'h10 ;
			data[6618] <= 8'h10 ;
			data[6619] <= 8'h10 ;
			data[6620] <= 8'h10 ;
			data[6621] <= 8'h10 ;
			data[6622] <= 8'h10 ;
			data[6623] <= 8'h10 ;
			data[6624] <= 8'h10 ;
			data[6625] <= 8'h10 ;
			data[6626] <= 8'h10 ;
			data[6627] <= 8'h10 ;
			data[6628] <= 8'h10 ;
			data[6629] <= 8'h10 ;
			data[6630] <= 8'h10 ;
			data[6631] <= 8'h10 ;
			data[6632] <= 8'h10 ;
			data[6633] <= 8'h10 ;
			data[6634] <= 8'h10 ;
			data[6635] <= 8'h10 ;
			data[6636] <= 8'h10 ;
			data[6637] <= 8'h10 ;
			data[6638] <= 8'h10 ;
			data[6639] <= 8'h10 ;
			data[6640] <= 8'h10 ;
			data[6641] <= 8'h10 ;
			data[6642] <= 8'h10 ;
			data[6643] <= 8'h10 ;
			data[6644] <= 8'h10 ;
			data[6645] <= 8'h10 ;
			data[6646] <= 8'h10 ;
			data[6647] <= 8'h10 ;
			data[6648] <= 8'h10 ;
			data[6649] <= 8'h10 ;
			data[6650] <= 8'h10 ;
			data[6651] <= 8'h10 ;
			data[6652] <= 8'h10 ;
			data[6653] <= 8'h10 ;
			data[6654] <= 8'h10 ;
			data[6655] <= 8'h10 ;
			data[6656] <= 8'h10 ;
			data[6657] <= 8'h10 ;
			data[6658] <= 8'h10 ;
			data[6659] <= 8'h10 ;
			data[6660] <= 8'h10 ;
			data[6661] <= 8'h10 ;
			data[6662] <= 8'h10 ;
			data[6663] <= 8'h10 ;
			data[6664] <= 8'h10 ;
			data[6665] <= 8'h10 ;
			data[6666] <= 8'h10 ;
			data[6667] <= 8'h10 ;
			data[6668] <= 8'h10 ;
			data[6669] <= 8'h10 ;
			data[6670] <= 8'h10 ;
			data[6671] <= 8'h10 ;
			data[6672] <= 8'h10 ;
			data[6673] <= 8'h10 ;
			data[6674] <= 8'h10 ;
			data[6675] <= 8'h10 ;
			data[6676] <= 8'h10 ;
			data[6677] <= 8'h10 ;
			data[6678] <= 8'h10 ;
			data[6679] <= 8'h10 ;
			data[6680] <= 8'h10 ;
			data[6681] <= 8'h10 ;
			data[6682] <= 8'h10 ;
			data[6683] <= 8'h10 ;
			data[6684] <= 8'h10 ;
			data[6685] <= 8'h10 ;
			data[6686] <= 8'h10 ;
			data[6687] <= 8'h10 ;
			data[6688] <= 8'h10 ;
			data[6689] <= 8'h10 ;
			data[6690] <= 8'h10 ;
			data[6691] <= 8'h10 ;
			data[6692] <= 8'h10 ;
			data[6693] <= 8'h10 ;
			data[6694] <= 8'h10 ;
			data[6695] <= 8'h10 ;
			data[6696] <= 8'h10 ;
			data[6697] <= 8'h10 ;
			data[6698] <= 8'h10 ;
			data[6699] <= 8'h10 ;
			data[6700] <= 8'h10 ;
			data[6701] <= 8'h10 ;
			data[6702] <= 8'h10 ;
			data[6703] <= 8'h10 ;
			data[6704] <= 8'h10 ;
			data[6705] <= 8'h10 ;
			data[6706] <= 8'h10 ;
			data[6707] <= 8'h10 ;
			data[6708] <= 8'h10 ;
			data[6709] <= 8'h10 ;
			data[6710] <= 8'h10 ;
			data[6711] <= 8'h10 ;
			data[6712] <= 8'h10 ;
			data[6713] <= 8'h10 ;
			data[6714] <= 8'h10 ;
			data[6715] <= 8'h10 ;
			data[6716] <= 8'h10 ;
			data[6717] <= 8'h10 ;
			data[6718] <= 8'h10 ;
			data[6719] <= 8'h10 ;
			data[6720] <= 8'h10 ;
			data[6721] <= 8'h10 ;
			data[6722] <= 8'h10 ;
			data[6723] <= 8'h10 ;
			data[6724] <= 8'h10 ;
			data[6725] <= 8'h10 ;
			data[6726] <= 8'h10 ;
			data[6727] <= 8'h10 ;
			data[6728] <= 8'h10 ;
			data[6729] <= 8'h10 ;
			data[6730] <= 8'h10 ;
			data[6731] <= 8'h10 ;
			data[6732] <= 8'h10 ;
			data[6733] <= 8'h10 ;
			data[6734] <= 8'h10 ;
			data[6735] <= 8'h10 ;
			data[6736] <= 8'h10 ;
			data[6737] <= 8'h10 ;
			data[6738] <= 8'h10 ;
			data[6739] <= 8'h10 ;
			data[6740] <= 8'h10 ;
			data[6741] <= 8'h10 ;
			data[6742] <= 8'h10 ;
			data[6743] <= 8'h10 ;
			data[6744] <= 8'h10 ;
			data[6745] <= 8'h10 ;
			data[6746] <= 8'h10 ;
			data[6747] <= 8'h10 ;
			data[6748] <= 8'h10 ;
			data[6749] <= 8'h10 ;
			data[6750] <= 8'h10 ;
			data[6751] <= 8'h10 ;
			data[6752] <= 8'h10 ;
			data[6753] <= 8'h10 ;
			data[6754] <= 8'h10 ;
			data[6755] <= 8'h10 ;
			data[6756] <= 8'h10 ;
			data[6757] <= 8'h10 ;
			data[6758] <= 8'h10 ;
			data[6759] <= 8'h10 ;
			data[6760] <= 8'h10 ;
			data[6761] <= 8'h10 ;
			data[6762] <= 8'h10 ;
			data[6763] <= 8'h10 ;
			data[6764] <= 8'h10 ;
			data[6765] <= 8'h10 ;
			data[6766] <= 8'h10 ;
			data[6767] <= 8'h10 ;
			data[6768] <= 8'h10 ;
			data[6769] <= 8'h10 ;
			data[6770] <= 8'h10 ;
			data[6771] <= 8'h10 ;
			data[6772] <= 8'h10 ;
			data[6773] <= 8'h10 ;
			data[6774] <= 8'h10 ;
			data[6775] <= 8'h10 ;
			data[6776] <= 8'h10 ;
			data[6777] <= 8'h10 ;
			data[6778] <= 8'h10 ;
			data[6779] <= 8'h10 ;
			data[6780] <= 8'h10 ;
			data[6781] <= 8'h10 ;
			data[6782] <= 8'h10 ;
			data[6783] <= 8'h10 ;
			data[6784] <= 8'h10 ;
			data[6785] <= 8'h10 ;
			data[6786] <= 8'h10 ;
			data[6787] <= 8'h10 ;
			data[6788] <= 8'h10 ;
			data[6789] <= 8'h10 ;
			data[6790] <= 8'h10 ;
			data[6791] <= 8'h10 ;
			data[6792] <= 8'h10 ;
			data[6793] <= 8'h10 ;
			data[6794] <= 8'h10 ;
			data[6795] <= 8'h10 ;
			data[6796] <= 8'h10 ;
			data[6797] <= 8'h10 ;
			data[6798] <= 8'h10 ;
			data[6799] <= 8'h10 ;
			data[6800] <= 8'h10 ;
			data[6801] <= 8'h10 ;
			data[6802] <= 8'h10 ;
			data[6803] <= 8'h10 ;
			data[6804] <= 8'h10 ;
			data[6805] <= 8'h10 ;
			data[6806] <= 8'h10 ;
			data[6807] <= 8'h10 ;
			data[6808] <= 8'h10 ;
			data[6809] <= 8'h10 ;
			data[6810] <= 8'h10 ;
			data[6811] <= 8'h10 ;
			data[6812] <= 8'h10 ;
			data[6813] <= 8'h10 ;
			data[6814] <= 8'h10 ;
			data[6815] <= 8'h10 ;
			data[6816] <= 8'h10 ;
			data[6817] <= 8'h10 ;
			data[6818] <= 8'h10 ;
			data[6819] <= 8'h10 ;
			data[6820] <= 8'h10 ;
			data[6821] <= 8'h10 ;
			data[6822] <= 8'h10 ;
			data[6823] <= 8'h10 ;
			data[6824] <= 8'h10 ;
			data[6825] <= 8'h10 ;
			data[6826] <= 8'h10 ;
			data[6827] <= 8'h10 ;
			data[6828] <= 8'h10 ;
			data[6829] <= 8'h10 ;
			data[6830] <= 8'h10 ;
			data[6831] <= 8'h10 ;
			data[6832] <= 8'h10 ;
			data[6833] <= 8'h10 ;
			data[6834] <= 8'h10 ;
			data[6835] <= 8'h10 ;
			data[6836] <= 8'h10 ;
			data[6837] <= 8'h10 ;
			data[6838] <= 8'h10 ;
			data[6839] <= 8'h10 ;
			data[6840] <= 8'h10 ;
			data[6841] <= 8'h10 ;
			data[6842] <= 8'h10 ;
			data[6843] <= 8'h10 ;
			data[6844] <= 8'h10 ;
			data[6845] <= 8'h10 ;
			data[6846] <= 8'h10 ;
			data[6847] <= 8'h10 ;
			data[6848] <= 8'h10 ;
			data[6849] <= 8'h10 ;
			data[6850] <= 8'h10 ;
			data[6851] <= 8'h10 ;
			data[6852] <= 8'h10 ;
			data[6853] <= 8'h10 ;
			data[6854] <= 8'h10 ;
			data[6855] <= 8'h10 ;
			data[6856] <= 8'h10 ;
			data[6857] <= 8'h10 ;
			data[6858] <= 8'h10 ;
			data[6859] <= 8'h10 ;
			data[6860] <= 8'h10 ;
			data[6861] <= 8'h10 ;
			data[6862] <= 8'h10 ;
			data[6863] <= 8'h10 ;
			data[6864] <= 8'h10 ;
			data[6865] <= 8'h10 ;
			data[6866] <= 8'h10 ;
			data[6867] <= 8'h10 ;
			data[6868] <= 8'h10 ;
			data[6869] <= 8'h10 ;
			data[6870] <= 8'h10 ;
			data[6871] <= 8'h10 ;
			data[6872] <= 8'h10 ;
			data[6873] <= 8'h10 ;
			data[6874] <= 8'h10 ;
			data[6875] <= 8'h10 ;
			data[6876] <= 8'h10 ;
			data[6877] <= 8'h10 ;
			data[6878] <= 8'h10 ;
			data[6879] <= 8'h10 ;
			data[6880] <= 8'h10 ;
			data[6881] <= 8'h10 ;
			data[6882] <= 8'h10 ;
			data[6883] <= 8'h10 ;
			data[6884] <= 8'h10 ;
			data[6885] <= 8'h10 ;
			data[6886] <= 8'h10 ;
			data[6887] <= 8'h10 ;
			data[6888] <= 8'h10 ;
			data[6889] <= 8'h10 ;
			data[6890] <= 8'h10 ;
			data[6891] <= 8'h10 ;
			data[6892] <= 8'h10 ;
			data[6893] <= 8'h10 ;
			data[6894] <= 8'h10 ;
			data[6895] <= 8'h10 ;
			data[6896] <= 8'h10 ;
			data[6897] <= 8'h10 ;
			data[6898] <= 8'h10 ;
			data[6899] <= 8'h10 ;
			data[6900] <= 8'h10 ;
			data[6901] <= 8'h10 ;
			data[6902] <= 8'h10 ;
			data[6903] <= 8'h10 ;
			data[6904] <= 8'h10 ;
			data[6905] <= 8'h10 ;
			data[6906] <= 8'h10 ;
			data[6907] <= 8'h10 ;
			data[6908] <= 8'h10 ;
			data[6909] <= 8'h10 ;
			data[6910] <= 8'h10 ;
			data[6911] <= 8'h10 ;
			data[6912] <= 8'h10 ;
			data[6913] <= 8'h10 ;
			data[6914] <= 8'h10 ;
			data[6915] <= 8'h10 ;
			data[6916] <= 8'h10 ;
			data[6917] <= 8'h10 ;
			data[6918] <= 8'h10 ;
			data[6919] <= 8'h10 ;
			data[6920] <= 8'h10 ;
			data[6921] <= 8'h10 ;
			data[6922] <= 8'h10 ;
			data[6923] <= 8'h10 ;
			data[6924] <= 8'h10 ;
			data[6925] <= 8'h10 ;
			data[6926] <= 8'h10 ;
			data[6927] <= 8'h10 ;
			data[6928] <= 8'h10 ;
			data[6929] <= 8'h10 ;
			data[6930] <= 8'h10 ;
			data[6931] <= 8'h10 ;
			data[6932] <= 8'h10 ;
			data[6933] <= 8'h10 ;
			data[6934] <= 8'h10 ;
			data[6935] <= 8'h10 ;
			data[6936] <= 8'h10 ;
			data[6937] <= 8'h10 ;
			data[6938] <= 8'h10 ;
			data[6939] <= 8'h10 ;
			data[6940] <= 8'h10 ;
			data[6941] <= 8'h10 ;
			data[6942] <= 8'h10 ;
			data[6943] <= 8'h10 ;
			data[6944] <= 8'h10 ;
			data[6945] <= 8'h10 ;
			data[6946] <= 8'h10 ;
			data[6947] <= 8'h10 ;
			data[6948] <= 8'h10 ;
			data[6949] <= 8'h10 ;
			data[6950] <= 8'h10 ;
			data[6951] <= 8'h10 ;
			data[6952] <= 8'h10 ;
			data[6953] <= 8'h10 ;
			data[6954] <= 8'h10 ;
			data[6955] <= 8'h10 ;
			data[6956] <= 8'h10 ;
			data[6957] <= 8'h10 ;
			data[6958] <= 8'h10 ;
			data[6959] <= 8'h10 ;
			data[6960] <= 8'h10 ;
			data[6961] <= 8'h10 ;
			data[6962] <= 8'h10 ;
			data[6963] <= 8'h10 ;
			data[6964] <= 8'h10 ;
			data[6965] <= 8'h10 ;
			data[6966] <= 8'h10 ;
			data[6967] <= 8'h10 ;
			data[6968] <= 8'h10 ;
			data[6969] <= 8'h10 ;
			data[6970] <= 8'h10 ;
			data[6971] <= 8'h10 ;
			data[6972] <= 8'h10 ;
			data[6973] <= 8'h10 ;
			data[6974] <= 8'h10 ;
			data[6975] <= 8'h10 ;
			data[6976] <= 8'h10 ;
			data[6977] <= 8'h10 ;
			data[6978] <= 8'h10 ;
			data[6979] <= 8'h10 ;
			data[6980] <= 8'h10 ;
			data[6981] <= 8'h10 ;
			data[6982] <= 8'h10 ;
			data[6983] <= 8'h10 ;
			data[6984] <= 8'h10 ;
			data[6985] <= 8'h10 ;
			data[6986] <= 8'h10 ;
			data[6987] <= 8'h10 ;
			data[6988] <= 8'h10 ;
			data[6989] <= 8'h10 ;
			data[6990] <= 8'h10 ;
			data[6991] <= 8'h10 ;
			data[6992] <= 8'h10 ;
			data[6993] <= 8'h10 ;
			data[6994] <= 8'h10 ;
			data[6995] <= 8'h10 ;
			data[6996] <= 8'h10 ;
			data[6997] <= 8'h10 ;
			data[6998] <= 8'h10 ;
			data[6999] <= 8'h10 ;
			data[7000] <= 8'h10 ;
			data[7001] <= 8'h10 ;
			data[7002] <= 8'h10 ;
			data[7003] <= 8'h10 ;
			data[7004] <= 8'h10 ;
			data[7005] <= 8'h10 ;
			data[7006] <= 8'h10 ;
			data[7007] <= 8'h10 ;
			data[7008] <= 8'h10 ;
			data[7009] <= 8'h10 ;
			data[7010] <= 8'h10 ;
			data[7011] <= 8'h10 ;
			data[7012] <= 8'h10 ;
			data[7013] <= 8'h10 ;
			data[7014] <= 8'h10 ;
			data[7015] <= 8'h10 ;
			data[7016] <= 8'h10 ;
			data[7017] <= 8'h10 ;
			data[7018] <= 8'h10 ;
			data[7019] <= 8'h10 ;
			data[7020] <= 8'h10 ;
			data[7021] <= 8'h10 ;
			data[7022] <= 8'h10 ;
			data[7023] <= 8'h10 ;
			data[7024] <= 8'h10 ;
			data[7025] <= 8'h10 ;
			data[7026] <= 8'h10 ;
			data[7027] <= 8'h10 ;
			data[7028] <= 8'h10 ;
			data[7029] <= 8'h10 ;
			data[7030] <= 8'h10 ;
			data[7031] <= 8'h10 ;
			data[7032] <= 8'h10 ;
			data[7033] <= 8'h10 ;
			data[7034] <= 8'h10 ;
			data[7035] <= 8'h10 ;
			data[7036] <= 8'h10 ;
			data[7037] <= 8'h10 ;
			data[7038] <= 8'h10 ;
			data[7039] <= 8'h10 ;
			data[7040] <= 8'h10 ;
			data[7041] <= 8'h10 ;
			data[7042] <= 8'h10 ;
			data[7043] <= 8'h10 ;
			data[7044] <= 8'h10 ;
			data[7045] <= 8'h10 ;
			data[7046] <= 8'h10 ;
			data[7047] <= 8'h10 ;
			data[7048] <= 8'h10 ;
			data[7049] <= 8'h10 ;
			data[7050] <= 8'h10 ;
			data[7051] <= 8'h10 ;
			data[7052] <= 8'h10 ;
			data[7053] <= 8'h10 ;
			data[7054] <= 8'h10 ;
			data[7055] <= 8'h10 ;
			data[7056] <= 8'h10 ;
			data[7057] <= 8'h10 ;
			data[7058] <= 8'h10 ;
			data[7059] <= 8'h10 ;
			data[7060] <= 8'h10 ;
			data[7061] <= 8'h10 ;
			data[7062] <= 8'h10 ;
			data[7063] <= 8'h10 ;
			data[7064] <= 8'h10 ;
			data[7065] <= 8'h10 ;
			data[7066] <= 8'h10 ;
			data[7067] <= 8'h10 ;
			data[7068] <= 8'h10 ;
			data[7069] <= 8'h10 ;
			data[7070] <= 8'h10 ;
			data[7071] <= 8'h10 ;
			data[7072] <= 8'h10 ;
			data[7073] <= 8'h10 ;
			data[7074] <= 8'h10 ;
			data[7075] <= 8'h10 ;
			data[7076] <= 8'h10 ;
			data[7077] <= 8'h10 ;
			data[7078] <= 8'h10 ;
			data[7079] <= 8'h10 ;
			data[7080] <= 8'h10 ;
			data[7081] <= 8'h10 ;
			data[7082] <= 8'h10 ;
			data[7083] <= 8'h10 ;
			data[7084] <= 8'h10 ;
			data[7085] <= 8'h10 ;
			data[7086] <= 8'h10 ;
			data[7087] <= 8'h10 ;
			data[7088] <= 8'h10 ;
			data[7089] <= 8'h10 ;
			data[7090] <= 8'h10 ;
			data[7091] <= 8'h10 ;
			data[7092] <= 8'h10 ;
			data[7093] <= 8'h10 ;
			data[7094] <= 8'h10 ;
			data[7095] <= 8'h10 ;
			data[7096] <= 8'h10 ;
			data[7097] <= 8'h10 ;
			data[7098] <= 8'h10 ;
			data[7099] <= 8'h10 ;
			data[7100] <= 8'h10 ;
			data[7101] <= 8'h10 ;
			data[7102] <= 8'h10 ;
			data[7103] <= 8'h10 ;
			data[7104] <= 8'h10 ;
			data[7105] <= 8'h10 ;
			data[7106] <= 8'h10 ;
			data[7107] <= 8'h10 ;
			data[7108] <= 8'h10 ;
			data[7109] <= 8'h10 ;
			data[7110] <= 8'h10 ;
			data[7111] <= 8'h10 ;
			data[7112] <= 8'h10 ;
			data[7113] <= 8'h10 ;
			data[7114] <= 8'h10 ;
			data[7115] <= 8'h10 ;
			data[7116] <= 8'h10 ;
			data[7117] <= 8'h10 ;
			data[7118] <= 8'h10 ;
			data[7119] <= 8'h10 ;
			data[7120] <= 8'h10 ;
			data[7121] <= 8'h10 ;
			data[7122] <= 8'h10 ;
			data[7123] <= 8'h10 ;
			data[7124] <= 8'h10 ;
			data[7125] <= 8'h10 ;
			data[7126] <= 8'h10 ;
			data[7127] <= 8'h10 ;
			data[7128] <= 8'h10 ;
			data[7129] <= 8'h10 ;
			data[7130] <= 8'h10 ;
			data[7131] <= 8'h10 ;
			data[7132] <= 8'h10 ;
			data[7133] <= 8'h10 ;
			data[7134] <= 8'h10 ;
			data[7135] <= 8'h10 ;
			data[7136] <= 8'h10 ;
			data[7137] <= 8'h10 ;
			data[7138] <= 8'h10 ;
			data[7139] <= 8'h10 ;
			data[7140] <= 8'h10 ;
			data[7141] <= 8'h10 ;
			data[7142] <= 8'h10 ;
			data[7143] <= 8'h10 ;
			data[7144] <= 8'h10 ;
			data[7145] <= 8'h10 ;
			data[7146] <= 8'h10 ;
			data[7147] <= 8'h10 ;
			data[7148] <= 8'h10 ;
			data[7149] <= 8'h10 ;
			data[7150] <= 8'h10 ;
			data[7151] <= 8'h10 ;
			data[7152] <= 8'h10 ;
			data[7153] <= 8'h10 ;
			data[7154] <= 8'h10 ;
			data[7155] <= 8'h10 ;
			data[7156] <= 8'h10 ;
			data[7157] <= 8'h10 ;
			data[7158] <= 8'h10 ;
			data[7159] <= 8'h10 ;
			data[7160] <= 8'h10 ;
			data[7161] <= 8'h10 ;
			data[7162] <= 8'h10 ;
			data[7163] <= 8'h10 ;
			data[7164] <= 8'h10 ;
			data[7165] <= 8'h10 ;
			data[7166] <= 8'h10 ;
			data[7167] <= 8'h10 ;
			data[7168] <= 8'h10 ;
			data[7169] <= 8'h10 ;
			data[7170] <= 8'h10 ;
			data[7171] <= 8'h10 ;
			data[7172] <= 8'h10 ;
			data[7173] <= 8'h10 ;
			data[7174] <= 8'h10 ;
			data[7175] <= 8'h10 ;
			data[7176] <= 8'h10 ;
			data[7177] <= 8'h10 ;
			data[7178] <= 8'h10 ;
			data[7179] <= 8'h10 ;
			data[7180] <= 8'h10 ;
			data[7181] <= 8'h10 ;
			data[7182] <= 8'h10 ;
			data[7183] <= 8'h10 ;
			data[7184] <= 8'h10 ;
			data[7185] <= 8'h10 ;
			data[7186] <= 8'h10 ;
			data[7187] <= 8'h10 ;
			data[7188] <= 8'h10 ;
			data[7189] <= 8'h10 ;
			data[7190] <= 8'h10 ;
			data[7191] <= 8'h10 ;
			data[7192] <= 8'h10 ;
			data[7193] <= 8'h10 ;
			data[7194] <= 8'h10 ;
			data[7195] <= 8'h10 ;
			data[7196] <= 8'h10 ;
			data[7197] <= 8'h10 ;
			data[7198] <= 8'h10 ;
			data[7199] <= 8'h10 ;
			data[7200] <= 8'h10 ;
			data[7201] <= 8'h10 ;
			data[7202] <= 8'h10 ;
			data[7203] <= 8'h10 ;
			data[7204] <= 8'h10 ;
			data[7205] <= 8'h10 ;
			data[7206] <= 8'h10 ;
			data[7207] <= 8'h10 ;
			data[7208] <= 8'h10 ;
			data[7209] <= 8'h10 ;
			data[7210] <= 8'h10 ;
			data[7211] <= 8'h10 ;
			data[7212] <= 8'h10 ;
			data[7213] <= 8'h10 ;
			data[7214] <= 8'h10 ;
			data[7215] <= 8'h10 ;
			data[7216] <= 8'h10 ;
			data[7217] <= 8'h10 ;
			data[7218] <= 8'h10 ;
			data[7219] <= 8'h10 ;
			data[7220] <= 8'h10 ;
			data[7221] <= 8'h10 ;
			data[7222] <= 8'h10 ;
			data[7223] <= 8'h10 ;
			data[7224] <= 8'h10 ;
			data[7225] <= 8'h10 ;
			data[7226] <= 8'h10 ;
			data[7227] <= 8'h10 ;
			data[7228] <= 8'h10 ;
			data[7229] <= 8'h10 ;
			data[7230] <= 8'h10 ;
			data[7231] <= 8'h10 ;
			data[7232] <= 8'h10 ;
			data[7233] <= 8'h10 ;
			data[7234] <= 8'h10 ;
			data[7235] <= 8'h10 ;
			data[7236] <= 8'h10 ;
			data[7237] <= 8'h10 ;
			data[7238] <= 8'h10 ;
			data[7239] <= 8'h10 ;
			data[7240] <= 8'h10 ;
			data[7241] <= 8'h10 ;
			data[7242] <= 8'h10 ;
			data[7243] <= 8'h10 ;
			data[7244] <= 8'h10 ;
			data[7245] <= 8'h10 ;
			data[7246] <= 8'h10 ;
			data[7247] <= 8'h10 ;
			data[7248] <= 8'h10 ;
			data[7249] <= 8'h10 ;
			data[7250] <= 8'h10 ;
			data[7251] <= 8'h10 ;
			data[7252] <= 8'h10 ;
			data[7253] <= 8'h10 ;
			data[7254] <= 8'h10 ;
			data[7255] <= 8'h10 ;
			data[7256] <= 8'h10 ;
			data[7257] <= 8'h10 ;
			data[7258] <= 8'h10 ;
			data[7259] <= 8'h10 ;
			data[7260] <= 8'h10 ;
			data[7261] <= 8'h10 ;
			data[7262] <= 8'h10 ;
			data[7263] <= 8'h10 ;
			data[7264] <= 8'h10 ;
			data[7265] <= 8'h10 ;
			data[7266] <= 8'h10 ;
			data[7267] <= 8'h10 ;
			data[7268] <= 8'h10 ;
			data[7269] <= 8'h10 ;
			data[7270] <= 8'h10 ;
			data[7271] <= 8'h10 ;
			data[7272] <= 8'h10 ;
			data[7273] <= 8'h10 ;
			data[7274] <= 8'h10 ;
			data[7275] <= 8'h10 ;
			data[7276] <= 8'h10 ;
			data[7277] <= 8'h10 ;
			data[7278] <= 8'h10 ;
			data[7279] <= 8'h10 ;
			data[7280] <= 8'h10 ;
			data[7281] <= 8'h10 ;
			data[7282] <= 8'h10 ;
			data[7283] <= 8'h10 ;
			data[7284] <= 8'h10 ;
			data[7285] <= 8'h10 ;
			data[7286] <= 8'h10 ;
			data[7287] <= 8'h10 ;
			data[7288] <= 8'h10 ;
			data[7289] <= 8'h10 ;
			data[7290] <= 8'h10 ;
			data[7291] <= 8'h10 ;
			data[7292] <= 8'h10 ;
			data[7293] <= 8'h10 ;
			data[7294] <= 8'h10 ;
			data[7295] <= 8'h10 ;
			data[7296] <= 8'h10 ;
			data[7297] <= 8'h10 ;
			data[7298] <= 8'h10 ;
			data[7299] <= 8'h10 ;
			data[7300] <= 8'h10 ;
			data[7301] <= 8'h10 ;
			data[7302] <= 8'h10 ;
			data[7303] <= 8'h10 ;
			data[7304] <= 8'h10 ;
			data[7305] <= 8'h10 ;
			data[7306] <= 8'h10 ;
			data[7307] <= 8'h10 ;
			data[7308] <= 8'h10 ;
			data[7309] <= 8'h10 ;
			data[7310] <= 8'h10 ;
			data[7311] <= 8'h10 ;
			data[7312] <= 8'h10 ;
			data[7313] <= 8'h10 ;
			data[7314] <= 8'h10 ;
			data[7315] <= 8'h10 ;
			data[7316] <= 8'h10 ;
			data[7317] <= 8'h10 ;
			data[7318] <= 8'h10 ;
			data[7319] <= 8'h10 ;
			data[7320] <= 8'h10 ;
			data[7321] <= 8'h10 ;
			data[7322] <= 8'h10 ;
			data[7323] <= 8'h10 ;
			data[7324] <= 8'h10 ;
			data[7325] <= 8'h10 ;
			data[7326] <= 8'h10 ;
			data[7327] <= 8'h10 ;
			data[7328] <= 8'h10 ;
			data[7329] <= 8'h10 ;
			data[7330] <= 8'h10 ;
			data[7331] <= 8'h10 ;
			data[7332] <= 8'h10 ;
			data[7333] <= 8'h10 ;
			data[7334] <= 8'h10 ;
			data[7335] <= 8'h10 ;
			data[7336] <= 8'h10 ;
			data[7337] <= 8'h10 ;
			data[7338] <= 8'h10 ;
			data[7339] <= 8'h10 ;
			data[7340] <= 8'h10 ;
			data[7341] <= 8'h10 ;
			data[7342] <= 8'h10 ;
			data[7343] <= 8'h10 ;
			data[7344] <= 8'h10 ;
			data[7345] <= 8'h10 ;
			data[7346] <= 8'h10 ;
			data[7347] <= 8'h10 ;
			data[7348] <= 8'h10 ;
			data[7349] <= 8'h10 ;
			data[7350] <= 8'h10 ;
			data[7351] <= 8'h10 ;
			data[7352] <= 8'h10 ;
			data[7353] <= 8'h10 ;
			data[7354] <= 8'h10 ;
			data[7355] <= 8'h10 ;
			data[7356] <= 8'h10 ;
			data[7357] <= 8'h10 ;
			data[7358] <= 8'h10 ;
			data[7359] <= 8'h10 ;
			data[7360] <= 8'h10 ;
			data[7361] <= 8'h10 ;
			data[7362] <= 8'h10 ;
			data[7363] <= 8'h10 ;
			data[7364] <= 8'h10 ;
			data[7365] <= 8'h10 ;
			data[7366] <= 8'h10 ;
			data[7367] <= 8'h10 ;
			data[7368] <= 8'h10 ;
			data[7369] <= 8'h10 ;
			data[7370] <= 8'h10 ;
			data[7371] <= 8'h10 ;
			data[7372] <= 8'h10 ;
			data[7373] <= 8'h10 ;
			data[7374] <= 8'h10 ;
			data[7375] <= 8'h10 ;
			data[7376] <= 8'h10 ;
			data[7377] <= 8'h10 ;
			data[7378] <= 8'h10 ;
			data[7379] <= 8'h10 ;
			data[7380] <= 8'h10 ;
			data[7381] <= 8'h10 ;
			data[7382] <= 8'h10 ;
			data[7383] <= 8'h10 ;
			data[7384] <= 8'h10 ;
			data[7385] <= 8'h10 ;
			data[7386] <= 8'h10 ;
			data[7387] <= 8'h10 ;
			data[7388] <= 8'h10 ;
			data[7389] <= 8'h10 ;
			data[7390] <= 8'h10 ;
			data[7391] <= 8'h10 ;
			data[7392] <= 8'h10 ;
			data[7393] <= 8'h10 ;
			data[7394] <= 8'h10 ;
			data[7395] <= 8'h10 ;
			data[7396] <= 8'h10 ;
			data[7397] <= 8'h10 ;
			data[7398] <= 8'h10 ;
			data[7399] <= 8'h10 ;
			data[7400] <= 8'h10 ;
			data[7401] <= 8'h10 ;
			data[7402] <= 8'h10 ;
			data[7403] <= 8'h10 ;
			data[7404] <= 8'h10 ;
			data[7405] <= 8'h10 ;
			data[7406] <= 8'h10 ;
			data[7407] <= 8'h10 ;
			data[7408] <= 8'h10 ;
			data[7409] <= 8'h10 ;
			data[7410] <= 8'h10 ;
			data[7411] <= 8'h10 ;
			data[7412] <= 8'h10 ;
			data[7413] <= 8'h10 ;
			data[7414] <= 8'h10 ;
			data[7415] <= 8'h10 ;
			data[7416] <= 8'h10 ;
			data[7417] <= 8'h10 ;
			data[7418] <= 8'h10 ;
			data[7419] <= 8'h10 ;
			data[7420] <= 8'h10 ;
			data[7421] <= 8'h10 ;
			data[7422] <= 8'h10 ;
			data[7423] <= 8'h10 ;
			data[7424] <= 8'h10 ;
			data[7425] <= 8'h10 ;
			data[7426] <= 8'h10 ;
			data[7427] <= 8'h10 ;
			data[7428] <= 8'h10 ;
			data[7429] <= 8'h10 ;
			data[7430] <= 8'h10 ;
			data[7431] <= 8'h10 ;
			data[7432] <= 8'h10 ;
			data[7433] <= 8'h10 ;
			data[7434] <= 8'h10 ;
			data[7435] <= 8'h10 ;
			data[7436] <= 8'h10 ;
			data[7437] <= 8'h10 ;
			data[7438] <= 8'h10 ;
			data[7439] <= 8'h10 ;
			data[7440] <= 8'h10 ;
			data[7441] <= 8'h10 ;
			data[7442] <= 8'h10 ;
			data[7443] <= 8'h10 ;
			data[7444] <= 8'h10 ;
			data[7445] <= 8'h10 ;
			data[7446] <= 8'h10 ;
			data[7447] <= 8'h10 ;
			data[7448] <= 8'h10 ;
			data[7449] <= 8'h10 ;
			data[7450] <= 8'h10 ;
			data[7451] <= 8'h10 ;
			data[7452] <= 8'h10 ;
			data[7453] <= 8'h10 ;
			data[7454] <= 8'h10 ;
			data[7455] <= 8'h10 ;
			data[7456] <= 8'h10 ;
			data[7457] <= 8'h10 ;
			data[7458] <= 8'h10 ;
			data[7459] <= 8'h10 ;
			data[7460] <= 8'h10 ;
			data[7461] <= 8'h10 ;
			data[7462] <= 8'h10 ;
			data[7463] <= 8'h10 ;
			data[7464] <= 8'h10 ;
			data[7465] <= 8'h10 ;
			data[7466] <= 8'h10 ;
			data[7467] <= 8'h10 ;
			data[7468] <= 8'h10 ;
			data[7469] <= 8'h10 ;
			data[7470] <= 8'h10 ;
			data[7471] <= 8'h10 ;
			data[7472] <= 8'h10 ;
			data[7473] <= 8'h10 ;
			data[7474] <= 8'h10 ;
			data[7475] <= 8'h10 ;
			data[7476] <= 8'h10 ;
			data[7477] <= 8'h10 ;
			data[7478] <= 8'h10 ;
			data[7479] <= 8'h10 ;
			data[7480] <= 8'h10 ;
			data[7481] <= 8'h10 ;
			data[7482] <= 8'h10 ;
			data[7483] <= 8'h10 ;
			data[7484] <= 8'h10 ;
			data[7485] <= 8'h10 ;
			data[7486] <= 8'h10 ;
			data[7487] <= 8'h10 ;
			data[7488] <= 8'h10 ;
			data[7489] <= 8'h10 ;
			data[7490] <= 8'h10 ;
			data[7491] <= 8'h10 ;
			data[7492] <= 8'h10 ;
			data[7493] <= 8'h10 ;
			data[7494] <= 8'h10 ;
			data[7495] <= 8'h10 ;
			data[7496] <= 8'h10 ;
			data[7497] <= 8'h10 ;
			data[7498] <= 8'h10 ;
			data[7499] <= 8'h10 ;
			data[7500] <= 8'h10 ;
			data[7501] <= 8'h10 ;
			data[7502] <= 8'h10 ;
			data[7503] <= 8'h10 ;
			data[7504] <= 8'h10 ;
			data[7505] <= 8'h10 ;
			data[7506] <= 8'h10 ;
			data[7507] <= 8'h10 ;
			data[7508] <= 8'h10 ;
			data[7509] <= 8'h10 ;
			data[7510] <= 8'h10 ;
			data[7511] <= 8'h10 ;
			data[7512] <= 8'h10 ;
			data[7513] <= 8'h10 ;
			data[7514] <= 8'h10 ;
			data[7515] <= 8'h10 ;
			data[7516] <= 8'h10 ;
			data[7517] <= 8'h10 ;
			data[7518] <= 8'h10 ;
			data[7519] <= 8'h10 ;
			data[7520] <= 8'h10 ;
			data[7521] <= 8'h10 ;
			data[7522] <= 8'h10 ;
			data[7523] <= 8'h10 ;
			data[7524] <= 8'h10 ;
			data[7525] <= 8'h10 ;
			data[7526] <= 8'h10 ;
			data[7527] <= 8'h10 ;
			data[7528] <= 8'h10 ;
			data[7529] <= 8'h10 ;
			data[7530] <= 8'h10 ;
			data[7531] <= 8'h10 ;
			data[7532] <= 8'h10 ;
			data[7533] <= 8'h10 ;
			data[7534] <= 8'h10 ;
			data[7535] <= 8'h10 ;
			data[7536] <= 8'h10 ;
			data[7537] <= 8'h10 ;
			data[7538] <= 8'h10 ;
			data[7539] <= 8'h10 ;
			data[7540] <= 8'h10 ;
			data[7541] <= 8'h10 ;
			data[7542] <= 8'h10 ;
			data[7543] <= 8'h10 ;
			data[7544] <= 8'h10 ;
			data[7545] <= 8'h10 ;
			data[7546] <= 8'h10 ;
			data[7547] <= 8'h10 ;
			data[7548] <= 8'h10 ;
			data[7549] <= 8'h10 ;
			data[7550] <= 8'h10 ;
			data[7551] <= 8'h10 ;
			data[7552] <= 8'h10 ;
			data[7553] <= 8'h10 ;
			data[7554] <= 8'h10 ;
			data[7555] <= 8'h10 ;
			data[7556] <= 8'h10 ;
			data[7557] <= 8'h10 ;
			data[7558] <= 8'h10 ;
			data[7559] <= 8'h10 ;
			data[7560] <= 8'h10 ;
			data[7561] <= 8'h10 ;
			data[7562] <= 8'h10 ;
			data[7563] <= 8'h10 ;
			data[7564] <= 8'h10 ;
			data[7565] <= 8'h10 ;
			data[7566] <= 8'h10 ;
			data[7567] <= 8'h10 ;
			data[7568] <= 8'h10 ;
			data[7569] <= 8'h10 ;
			data[7570] <= 8'h10 ;
			data[7571] <= 8'h10 ;
			data[7572] <= 8'h10 ;
			data[7573] <= 8'h10 ;
			data[7574] <= 8'h10 ;
			data[7575] <= 8'h10 ;
			data[7576] <= 8'h10 ;
			data[7577] <= 8'h10 ;
			data[7578] <= 8'h10 ;
			data[7579] <= 8'h10 ;
			data[7580] <= 8'h10 ;
			data[7581] <= 8'h10 ;
			data[7582] <= 8'h10 ;
			data[7583] <= 8'h10 ;
			data[7584] <= 8'h10 ;
			data[7585] <= 8'h10 ;
			data[7586] <= 8'h10 ;
			data[7587] <= 8'h10 ;
			data[7588] <= 8'h10 ;
			data[7589] <= 8'h10 ;
			data[7590] <= 8'h10 ;
			data[7591] <= 8'h10 ;
			data[7592] <= 8'h10 ;
			data[7593] <= 8'h10 ;
			data[7594] <= 8'h10 ;
			data[7595] <= 8'h10 ;
			data[7596] <= 8'h10 ;
			data[7597] <= 8'h10 ;
			data[7598] <= 8'h10 ;
			data[7599] <= 8'h10 ;
			data[7600] <= 8'h10 ;
			data[7601] <= 8'h10 ;
			data[7602] <= 8'h10 ;
			data[7603] <= 8'h10 ;
			data[7604] <= 8'h10 ;
			data[7605] <= 8'h10 ;
			data[7606] <= 8'h10 ;
			data[7607] <= 8'h10 ;
			data[7608] <= 8'h10 ;
			data[7609] <= 8'h10 ;
			data[7610] <= 8'h10 ;
			data[7611] <= 8'h10 ;
			data[7612] <= 8'h10 ;
			data[7613] <= 8'h10 ;
			data[7614] <= 8'h10 ;
			data[7615] <= 8'h10 ;
			data[7616] <= 8'h10 ;
			data[7617] <= 8'h10 ;
			data[7618] <= 8'h10 ;
			data[7619] <= 8'h10 ;
			data[7620] <= 8'h10 ;
			data[7621] <= 8'h10 ;
			data[7622] <= 8'h10 ;
			data[7623] <= 8'h10 ;
			data[7624] <= 8'h10 ;
			data[7625] <= 8'h10 ;
			data[7626] <= 8'h10 ;
			data[7627] <= 8'h10 ;
			data[7628] <= 8'h10 ;
			data[7629] <= 8'h10 ;
			data[7630] <= 8'h10 ;
			data[7631] <= 8'h10 ;
			data[7632] <= 8'h10 ;
			data[7633] <= 8'h10 ;
			data[7634] <= 8'h10 ;
			data[7635] <= 8'h10 ;
			data[7636] <= 8'h10 ;
			data[7637] <= 8'h10 ;
			data[7638] <= 8'h10 ;
			data[7639] <= 8'h10 ;
			data[7640] <= 8'h10 ;
			data[7641] <= 8'h10 ;
			data[7642] <= 8'h10 ;
			data[7643] <= 8'h10 ;
			data[7644] <= 8'h10 ;
			data[7645] <= 8'h10 ;
			data[7646] <= 8'h10 ;
			data[7647] <= 8'h10 ;
			data[7648] <= 8'h10 ;
			data[7649] <= 8'h10 ;
			data[7650] <= 8'h10 ;
			data[7651] <= 8'h10 ;
			data[7652] <= 8'h10 ;
			data[7653] <= 8'h10 ;
			data[7654] <= 8'h10 ;
			data[7655] <= 8'h10 ;
			data[7656] <= 8'h10 ;
			data[7657] <= 8'h10 ;
			data[7658] <= 8'h10 ;
			data[7659] <= 8'h10 ;
			data[7660] <= 8'h10 ;
			data[7661] <= 8'h10 ;
			data[7662] <= 8'h10 ;
			data[7663] <= 8'h10 ;
			data[7664] <= 8'h10 ;
			data[7665] <= 8'h10 ;
			data[7666] <= 8'h10 ;
			data[7667] <= 8'h10 ;
			data[7668] <= 8'h10 ;
			data[7669] <= 8'h10 ;
			data[7670] <= 8'h10 ;
			data[7671] <= 8'h10 ;
			data[7672] <= 8'h10 ;
			data[7673] <= 8'h10 ;
			data[7674] <= 8'h10 ;
			data[7675] <= 8'h10 ;
			data[7676] <= 8'h10 ;
			data[7677] <= 8'h10 ;
			data[7678] <= 8'h10 ;
			data[7679] <= 8'h10 ;
			data[7680] <= 8'h10 ;
			data[7681] <= 8'h10 ;
			data[7682] <= 8'h10 ;
			data[7683] <= 8'h10 ;
			data[7684] <= 8'h10 ;
			data[7685] <= 8'h10 ;
			data[7686] <= 8'h10 ;
			data[7687] <= 8'h10 ;
			data[7688] <= 8'h10 ;
			data[7689] <= 8'h10 ;
			data[7690] <= 8'h10 ;
			data[7691] <= 8'h10 ;
			data[7692] <= 8'h10 ;
			data[7693] <= 8'h10 ;
			data[7694] <= 8'h10 ;
			data[7695] <= 8'h10 ;
			data[7696] <= 8'h10 ;
			data[7697] <= 8'h10 ;
			data[7698] <= 8'h10 ;
			data[7699] <= 8'h10 ;
			data[7700] <= 8'h10 ;
			data[7701] <= 8'h10 ;
			data[7702] <= 8'h10 ;
			data[7703] <= 8'h10 ;
			data[7704] <= 8'h10 ;
			data[7705] <= 8'h10 ;
			data[7706] <= 8'h10 ;
			data[7707] <= 8'h10 ;
			data[7708] <= 8'h10 ;
			data[7709] <= 8'h10 ;
			data[7710] <= 8'h10 ;
			data[7711] <= 8'h10 ;
			data[7712] <= 8'h10 ;
			data[7713] <= 8'h10 ;
			data[7714] <= 8'h10 ;
			data[7715] <= 8'h10 ;
			data[7716] <= 8'h10 ;
			data[7717] <= 8'h10 ;
			data[7718] <= 8'h10 ;
			data[7719] <= 8'h10 ;
			data[7720] <= 8'h10 ;
			data[7721] <= 8'h10 ;
			data[7722] <= 8'h10 ;
			data[7723] <= 8'h10 ;
			data[7724] <= 8'h10 ;
			data[7725] <= 8'h10 ;
			data[7726] <= 8'h10 ;
			data[7727] <= 8'h10 ;
			data[7728] <= 8'h10 ;
			data[7729] <= 8'h10 ;
			data[7730] <= 8'h10 ;
			data[7731] <= 8'h10 ;
			data[7732] <= 8'h10 ;
			data[7733] <= 8'h10 ;
			data[7734] <= 8'h10 ;
			data[7735] <= 8'h10 ;
			data[7736] <= 8'h10 ;
			data[7737] <= 8'h10 ;
			data[7738] <= 8'h10 ;
			data[7739] <= 8'h10 ;
			data[7740] <= 8'h10 ;
			data[7741] <= 8'h10 ;
			data[7742] <= 8'h10 ;
			data[7743] <= 8'h10 ;
			data[7744] <= 8'h10 ;
			data[7745] <= 8'h10 ;
			data[7746] <= 8'h10 ;
			data[7747] <= 8'h10 ;
			data[7748] <= 8'h10 ;
			data[7749] <= 8'h10 ;
			data[7750] <= 8'h10 ;
			data[7751] <= 8'h10 ;
			data[7752] <= 8'h10 ;
			data[7753] <= 8'h10 ;
			data[7754] <= 8'h10 ;
			data[7755] <= 8'h10 ;
			data[7756] <= 8'h10 ;
			data[7757] <= 8'h10 ;
			data[7758] <= 8'h10 ;
			data[7759] <= 8'h10 ;
			data[7760] <= 8'h10 ;
			data[7761] <= 8'h10 ;
			data[7762] <= 8'h10 ;
			data[7763] <= 8'h10 ;
			data[7764] <= 8'h10 ;
			data[7765] <= 8'h10 ;
			data[7766] <= 8'h10 ;
			data[7767] <= 8'h10 ;
			data[7768] <= 8'h10 ;
			data[7769] <= 8'h10 ;
			data[7770] <= 8'h10 ;
			data[7771] <= 8'h10 ;
			data[7772] <= 8'h10 ;
			data[7773] <= 8'h10 ;
			data[7774] <= 8'h10 ;
			data[7775] <= 8'h10 ;
			data[7776] <= 8'h10 ;
			data[7777] <= 8'h10 ;
			data[7778] <= 8'h10 ;
			data[7779] <= 8'h10 ;
			data[7780] <= 8'h10 ;
			data[7781] <= 8'h10 ;
			data[7782] <= 8'h10 ;
			data[7783] <= 8'h10 ;
			data[7784] <= 8'h10 ;
			data[7785] <= 8'h10 ;
			data[7786] <= 8'h10 ;
			data[7787] <= 8'h10 ;
			data[7788] <= 8'h10 ;
			data[7789] <= 8'h10 ;
			data[7790] <= 8'h10 ;
			data[7791] <= 8'h10 ;
			data[7792] <= 8'h10 ;
			data[7793] <= 8'h10 ;
			data[7794] <= 8'h10 ;
			data[7795] <= 8'h10 ;
			data[7796] <= 8'h10 ;
			data[7797] <= 8'h10 ;
			data[7798] <= 8'h10 ;
			data[7799] <= 8'h10 ;
			data[7800] <= 8'h10 ;
			data[7801] <= 8'h10 ;
			data[7802] <= 8'h10 ;
			data[7803] <= 8'h10 ;
			data[7804] <= 8'h10 ;
			data[7805] <= 8'h10 ;
			data[7806] <= 8'h10 ;
			data[7807] <= 8'h10 ;
			data[7808] <= 8'h10 ;
			data[7809] <= 8'h10 ;
			data[7810] <= 8'h10 ;
			data[7811] <= 8'h10 ;
			data[7812] <= 8'h10 ;
			data[7813] <= 8'h10 ;
			data[7814] <= 8'h10 ;
			data[7815] <= 8'h10 ;
			data[7816] <= 8'h10 ;
			data[7817] <= 8'h10 ;
			data[7818] <= 8'h10 ;
			data[7819] <= 8'h10 ;
			data[7820] <= 8'h10 ;
			data[7821] <= 8'h10 ;
			data[7822] <= 8'h10 ;
			data[7823] <= 8'h10 ;
			data[7824] <= 8'h10 ;
			data[7825] <= 8'h10 ;
			data[7826] <= 8'h10 ;
			data[7827] <= 8'h10 ;
			data[7828] <= 8'h10 ;
			data[7829] <= 8'h10 ;
			data[7830] <= 8'h10 ;
			data[7831] <= 8'h10 ;
			data[7832] <= 8'h10 ;
			data[7833] <= 8'h10 ;
			data[7834] <= 8'h10 ;
			data[7835] <= 8'h10 ;
			data[7836] <= 8'h10 ;
			data[7837] <= 8'h10 ;
			data[7838] <= 8'h10 ;
			data[7839] <= 8'h10 ;
			data[7840] <= 8'h10 ;
			data[7841] <= 8'h10 ;
			data[7842] <= 8'h10 ;
			data[7843] <= 8'h10 ;
			data[7844] <= 8'h10 ;
			data[7845] <= 8'h10 ;
			data[7846] <= 8'h10 ;
			data[7847] <= 8'h10 ;
			data[7848] <= 8'h10 ;
			data[7849] <= 8'h10 ;
			data[7850] <= 8'h10 ;
			data[7851] <= 8'h10 ;
			data[7852] <= 8'h10 ;
			data[7853] <= 8'h10 ;
			data[7854] <= 8'h10 ;
			data[7855] <= 8'h10 ;
			data[7856] <= 8'h10 ;
			data[7857] <= 8'h10 ;
			data[7858] <= 8'h10 ;
			data[7859] <= 8'h10 ;
			data[7860] <= 8'h10 ;
			data[7861] <= 8'h10 ;
			data[7862] <= 8'h10 ;
			data[7863] <= 8'h10 ;
			data[7864] <= 8'h10 ;
			data[7865] <= 8'h10 ;
			data[7866] <= 8'h10 ;
			data[7867] <= 8'h10 ;
			data[7868] <= 8'h10 ;
			data[7869] <= 8'h10 ;
			data[7870] <= 8'h10 ;
			data[7871] <= 8'h10 ;
			data[7872] <= 8'h10 ;
			data[7873] <= 8'h10 ;
			data[7874] <= 8'h10 ;
			data[7875] <= 8'h10 ;
			data[7876] <= 8'h10 ;
			data[7877] <= 8'h10 ;
			data[7878] <= 8'h10 ;
			data[7879] <= 8'h10 ;
			data[7880] <= 8'h10 ;
			data[7881] <= 8'h10 ;
			data[7882] <= 8'h10 ;
			data[7883] <= 8'h10 ;
			data[7884] <= 8'h10 ;
			data[7885] <= 8'h10 ;
			data[7886] <= 8'h10 ;
			data[7887] <= 8'h10 ;
			data[7888] <= 8'h10 ;
			data[7889] <= 8'h10 ;
			data[7890] <= 8'h10 ;
			data[7891] <= 8'h10 ;
			data[7892] <= 8'h10 ;
			data[7893] <= 8'h10 ;
			data[7894] <= 8'h10 ;
			data[7895] <= 8'h10 ;
			data[7896] <= 8'h10 ;
			data[7897] <= 8'h10 ;
			data[7898] <= 8'h10 ;
			data[7899] <= 8'h10 ;
			data[7900] <= 8'h10 ;
			data[7901] <= 8'h10 ;
			data[7902] <= 8'h10 ;
			data[7903] <= 8'h10 ;
			data[7904] <= 8'h10 ;
			data[7905] <= 8'h10 ;
			data[7906] <= 8'h10 ;
			data[7907] <= 8'h10 ;
			data[7908] <= 8'h10 ;
			data[7909] <= 8'h10 ;
			data[7910] <= 8'h10 ;
			data[7911] <= 8'h10 ;
			data[7912] <= 8'h10 ;
			data[7913] <= 8'h10 ;
			data[7914] <= 8'h10 ;
			data[7915] <= 8'h10 ;
			data[7916] <= 8'h10 ;
			data[7917] <= 8'h10 ;
			data[7918] <= 8'h10 ;
			data[7919] <= 8'h10 ;
			data[7920] <= 8'h10 ;
			data[7921] <= 8'h10 ;
			data[7922] <= 8'h10 ;
			data[7923] <= 8'h10 ;
			data[7924] <= 8'h10 ;
			data[7925] <= 8'h10 ;
			data[7926] <= 8'h10 ;
			data[7927] <= 8'h10 ;
			data[7928] <= 8'h10 ;
			data[7929] <= 8'h10 ;
			data[7930] <= 8'h10 ;
			data[7931] <= 8'h10 ;
			data[7932] <= 8'h10 ;
			data[7933] <= 8'h10 ;
			data[7934] <= 8'h10 ;
			data[7935] <= 8'h10 ;
			data[7936] <= 8'h10 ;
			data[7937] <= 8'h10 ;
			data[7938] <= 8'h10 ;
			data[7939] <= 8'h10 ;
			data[7940] <= 8'h10 ;
			data[7941] <= 8'h10 ;
			data[7942] <= 8'h10 ;
			data[7943] <= 8'h10 ;
			data[7944] <= 8'h10 ;
			data[7945] <= 8'h10 ;
			data[7946] <= 8'h10 ;
			data[7947] <= 8'h10 ;
			data[7948] <= 8'h10 ;
			data[7949] <= 8'h10 ;
			data[7950] <= 8'h10 ;
			data[7951] <= 8'h10 ;
			data[7952] <= 8'h10 ;
			data[7953] <= 8'h10 ;
			data[7954] <= 8'h10 ;
			data[7955] <= 8'h10 ;
			data[7956] <= 8'h10 ;
			data[7957] <= 8'h10 ;
			data[7958] <= 8'h10 ;
			data[7959] <= 8'h10 ;
			data[7960] <= 8'h10 ;
			data[7961] <= 8'h10 ;
			data[7962] <= 8'h10 ;
			data[7963] <= 8'h10 ;
			data[7964] <= 8'h10 ;
			data[7965] <= 8'h10 ;
			data[7966] <= 8'h10 ;
			data[7967] <= 8'h10 ;
			data[7968] <= 8'h10 ;
			data[7969] <= 8'h10 ;
			data[7970] <= 8'h10 ;
			data[7971] <= 8'h10 ;
			data[7972] <= 8'h10 ;
			data[7973] <= 8'h10 ;
			data[7974] <= 8'h10 ;
			data[7975] <= 8'h10 ;
			data[7976] <= 8'h10 ;
			data[7977] <= 8'h10 ;
			data[7978] <= 8'h10 ;
			data[7979] <= 8'h10 ;
			data[7980] <= 8'h10 ;
			data[7981] <= 8'h10 ;
			data[7982] <= 8'h10 ;
			data[7983] <= 8'h10 ;
			data[7984] <= 8'h10 ;
			data[7985] <= 8'h10 ;
			data[7986] <= 8'h10 ;
			data[7987] <= 8'h10 ;
			data[7988] <= 8'h10 ;
			data[7989] <= 8'h10 ;
			data[7990] <= 8'h10 ;
			data[7991] <= 8'h10 ;
			data[7992] <= 8'h10 ;
			data[7993] <= 8'h10 ;
			data[7994] <= 8'h10 ;
			data[7995] <= 8'h10 ;
			data[7996] <= 8'h10 ;
			data[7997] <= 8'h10 ;
			data[7998] <= 8'h10 ;
			data[7999] <= 8'h10 ;
			data[8000] <= 8'h10 ;
			data[8001] <= 8'h10 ;
			data[8002] <= 8'h10 ;
			data[8003] <= 8'h10 ;
			data[8004] <= 8'h10 ;
			data[8005] <= 8'h10 ;
			data[8006] <= 8'h10 ;
			data[8007] <= 8'h10 ;
			data[8008] <= 8'h10 ;
			data[8009] <= 8'h10 ;
			data[8010] <= 8'h10 ;
			data[8011] <= 8'h10 ;
			data[8012] <= 8'h10 ;
			data[8013] <= 8'h10 ;
			data[8014] <= 8'h10 ;
			data[8015] <= 8'h10 ;
			data[8016] <= 8'h10 ;
			data[8017] <= 8'h10 ;
			data[8018] <= 8'h10 ;
			data[8019] <= 8'h10 ;
			data[8020] <= 8'h10 ;
			data[8021] <= 8'h10 ;
			data[8022] <= 8'h10 ;
			data[8023] <= 8'h10 ;
			data[8024] <= 8'h10 ;
			data[8025] <= 8'h10 ;
			data[8026] <= 8'h10 ;
			data[8027] <= 8'h10 ;
			data[8028] <= 8'h10 ;
			data[8029] <= 8'h10 ;
			data[8030] <= 8'h10 ;
			data[8031] <= 8'h10 ;
			data[8032] <= 8'h10 ;
			data[8033] <= 8'h10 ;
			data[8034] <= 8'h10 ;
			data[8035] <= 8'h10 ;
			data[8036] <= 8'h10 ;
			data[8037] <= 8'h10 ;
			data[8038] <= 8'h10 ;
			data[8039] <= 8'h10 ;
			data[8040] <= 8'h10 ;
			data[8041] <= 8'h10 ;
			data[8042] <= 8'h10 ;
			data[8043] <= 8'h10 ;
			data[8044] <= 8'h10 ;
			data[8045] <= 8'h10 ;
			data[8046] <= 8'h10 ;
			data[8047] <= 8'h10 ;
			data[8048] <= 8'h10 ;
			data[8049] <= 8'h10 ;
			data[8050] <= 8'h10 ;
			data[8051] <= 8'h10 ;
			data[8052] <= 8'h10 ;
			data[8053] <= 8'h10 ;
			data[8054] <= 8'h10 ;
			data[8055] <= 8'h10 ;
			data[8056] <= 8'h10 ;
			data[8057] <= 8'h10 ;
			data[8058] <= 8'h10 ;
			data[8059] <= 8'h10 ;
			data[8060] <= 8'h10 ;
			data[8061] <= 8'h10 ;
			data[8062] <= 8'h10 ;
			data[8063] <= 8'h10 ;
			data[8064] <= 8'h10 ;
			data[8065] <= 8'h10 ;
			data[8066] <= 8'h10 ;
			data[8067] <= 8'h10 ;
			data[8068] <= 8'h10 ;
			data[8069] <= 8'h10 ;
			data[8070] <= 8'h10 ;
			data[8071] <= 8'h10 ;
			data[8072] <= 8'h10 ;
			data[8073] <= 8'h10 ;
			data[8074] <= 8'h10 ;
			data[8075] <= 8'h10 ;
			data[8076] <= 8'h10 ;
			data[8077] <= 8'h10 ;
			data[8078] <= 8'h10 ;
			data[8079] <= 8'h10 ;
			data[8080] <= 8'h10 ;
			data[8081] <= 8'h10 ;
			data[8082] <= 8'h10 ;
			data[8083] <= 8'h10 ;
			data[8084] <= 8'h10 ;
			data[8085] <= 8'h10 ;
			data[8086] <= 8'h10 ;
			data[8087] <= 8'h10 ;
			data[8088] <= 8'h10 ;
			data[8089] <= 8'h10 ;
			data[8090] <= 8'h10 ;
			data[8091] <= 8'h10 ;
			data[8092] <= 8'h10 ;
			data[8093] <= 8'h10 ;
			data[8094] <= 8'h10 ;
			data[8095] <= 8'h10 ;
			data[8096] <= 8'h10 ;
			data[8097] <= 8'h10 ;
			data[8098] <= 8'h10 ;
			data[8099] <= 8'h10 ;
			data[8100] <= 8'h10 ;
			data[8101] <= 8'h10 ;
			data[8102] <= 8'h10 ;
			data[8103] <= 8'h10 ;
			data[8104] <= 8'h10 ;
			data[8105] <= 8'h10 ;
			data[8106] <= 8'h10 ;
			data[8107] <= 8'h10 ;
			data[8108] <= 8'h10 ;
			data[8109] <= 8'h10 ;
			data[8110] <= 8'h10 ;
			data[8111] <= 8'h10 ;
			data[8112] <= 8'h10 ;
			data[8113] <= 8'h10 ;
			data[8114] <= 8'h10 ;
			data[8115] <= 8'h10 ;
			data[8116] <= 8'h10 ;
			data[8117] <= 8'h10 ;
			data[8118] <= 8'h10 ;
			data[8119] <= 8'h10 ;
			data[8120] <= 8'h10 ;
			data[8121] <= 8'h10 ;
			data[8122] <= 8'h10 ;
			data[8123] <= 8'h10 ;
			data[8124] <= 8'h10 ;
			data[8125] <= 8'h10 ;
			data[8126] <= 8'h10 ;
			data[8127] <= 8'h10 ;
			data[8128] <= 8'h10 ;
			data[8129] <= 8'h10 ;
			data[8130] <= 8'h10 ;
			data[8131] <= 8'h10 ;
			data[8132] <= 8'h10 ;
			data[8133] <= 8'h10 ;
			data[8134] <= 8'h10 ;
			data[8135] <= 8'h10 ;
			data[8136] <= 8'h10 ;
			data[8137] <= 8'h10 ;
			data[8138] <= 8'h10 ;
			data[8139] <= 8'h10 ;
			data[8140] <= 8'h10 ;
			data[8141] <= 8'h10 ;
			data[8142] <= 8'h10 ;
			data[8143] <= 8'h10 ;
			data[8144] <= 8'h10 ;
			data[8145] <= 8'h10 ;
			data[8146] <= 8'h10 ;
			data[8147] <= 8'h10 ;
			data[8148] <= 8'h10 ;
			data[8149] <= 8'h10 ;
			data[8150] <= 8'h10 ;
			data[8151] <= 8'h10 ;
			data[8152] <= 8'h10 ;
			data[8153] <= 8'h10 ;
			data[8154] <= 8'h10 ;
			data[8155] <= 8'h10 ;
			data[8156] <= 8'h10 ;
			data[8157] <= 8'h10 ;
			data[8158] <= 8'h10 ;
			data[8159] <= 8'h10 ;
			data[8160] <= 8'h10 ;
			data[8161] <= 8'h10 ;
			data[8162] <= 8'h10 ;
			data[8163] <= 8'h10 ;
			data[8164] <= 8'h10 ;
			data[8165] <= 8'h10 ;
			data[8166] <= 8'h10 ;
			data[8167] <= 8'h10 ;
			data[8168] <= 8'h10 ;
			data[8169] <= 8'h10 ;
			data[8170] <= 8'h10 ;
			data[8171] <= 8'h10 ;
			data[8172] <= 8'h10 ;
			data[8173] <= 8'h10 ;
			data[8174] <= 8'h10 ;
			data[8175] <= 8'h10 ;
			data[8176] <= 8'h10 ;
			data[8177] <= 8'h10 ;
			data[8178] <= 8'h10 ;
			data[8179] <= 8'h10 ;
			data[8180] <= 8'h10 ;
			data[8181] <= 8'h10 ;
			data[8182] <= 8'h10 ;
			data[8183] <= 8'h10 ;
			data[8184] <= 8'h10 ;
			data[8185] <= 8'h10 ;
			data[8186] <= 8'h10 ;
			data[8187] <= 8'h10 ;
			data[8188] <= 8'h10 ;
			data[8189] <= 8'h10 ;
			data[8190] <= 8'h10 ;
			data[8191] <= 8'h10 ;
			data[8192] <= 8'h10 ;
			data[8193] <= 8'h10 ;
			data[8194] <= 8'h10 ;
			data[8195] <= 8'h10 ;
			data[8196] <= 8'h10 ;
			data[8197] <= 8'h10 ;
			data[8198] <= 8'h10 ;
			data[8199] <= 8'h10 ;
			data[8200] <= 8'h10 ;
			data[8201] <= 8'h10 ;
			data[8202] <= 8'h10 ;
			data[8203] <= 8'h10 ;
			data[8204] <= 8'h10 ;
			data[8205] <= 8'h10 ;
			data[8206] <= 8'h10 ;
			data[8207] <= 8'h10 ;
			data[8208] <= 8'h10 ;
			data[8209] <= 8'h10 ;
			data[8210] <= 8'h10 ;
			data[8211] <= 8'h10 ;
			data[8212] <= 8'h10 ;
			data[8213] <= 8'h10 ;
			data[8214] <= 8'h10 ;
			data[8215] <= 8'h10 ;
			data[8216] <= 8'h10 ;
			data[8217] <= 8'h10 ;
			data[8218] <= 8'h10 ;
			data[8219] <= 8'h10 ;
			data[8220] <= 8'h10 ;
			data[8221] <= 8'h10 ;
			data[8222] <= 8'h10 ;
			data[8223] <= 8'h10 ;
			data[8224] <= 8'h10 ;
			data[8225] <= 8'h10 ;
			data[8226] <= 8'h10 ;
			data[8227] <= 8'h10 ;
			data[8228] <= 8'h10 ;
			data[8229] <= 8'h10 ;
			data[8230] <= 8'h10 ;
			data[8231] <= 8'h10 ;
			data[8232] <= 8'h10 ;
			data[8233] <= 8'h10 ;
			data[8234] <= 8'h10 ;
			data[8235] <= 8'h10 ;
			data[8236] <= 8'h10 ;
			data[8237] <= 8'h10 ;
			data[8238] <= 8'h10 ;
			data[8239] <= 8'h10 ;
			data[8240] <= 8'h10 ;
			data[8241] <= 8'h10 ;
			data[8242] <= 8'h10 ;
			data[8243] <= 8'h10 ;
			data[8244] <= 8'h10 ;
			data[8245] <= 8'h10 ;
			data[8246] <= 8'h10 ;
			data[8247] <= 8'h10 ;
			data[8248] <= 8'h10 ;
			data[8249] <= 8'h10 ;
			data[8250] <= 8'h10 ;
			data[8251] <= 8'h10 ;
			data[8252] <= 8'h10 ;
			data[8253] <= 8'h10 ;
			data[8254] <= 8'h10 ;
			data[8255] <= 8'h10 ;
			data[8256] <= 8'h10 ;
			data[8257] <= 8'h10 ;
			data[8258] <= 8'h10 ;
			data[8259] <= 8'h10 ;
			data[8260] <= 8'h10 ;
			data[8261] <= 8'h10 ;
			data[8262] <= 8'h10 ;
			data[8263] <= 8'h10 ;
			data[8264] <= 8'h10 ;
			data[8265] <= 8'h10 ;
			data[8266] <= 8'h10 ;
			data[8267] <= 8'h10 ;
			data[8268] <= 8'h10 ;
			data[8269] <= 8'h10 ;
			data[8270] <= 8'h10 ;
			data[8271] <= 8'h10 ;
			data[8272] <= 8'h10 ;
			data[8273] <= 8'h10 ;
			data[8274] <= 8'h10 ;
			data[8275] <= 8'h10 ;
			data[8276] <= 8'h10 ;
			data[8277] <= 8'h10 ;
			data[8278] <= 8'h10 ;
			data[8279] <= 8'h10 ;
			data[8280] <= 8'h10 ;
			data[8281] <= 8'h10 ;
			data[8282] <= 8'h10 ;
			data[8283] <= 8'h10 ;
			data[8284] <= 8'h10 ;
			data[8285] <= 8'h10 ;
			data[8286] <= 8'h10 ;
			data[8287] <= 8'h10 ;
			data[8288] <= 8'h10 ;
			data[8289] <= 8'h10 ;
			data[8290] <= 8'h10 ;
			data[8291] <= 8'h10 ;
			data[8292] <= 8'h10 ;
			data[8293] <= 8'h10 ;
			data[8294] <= 8'h10 ;
			data[8295] <= 8'h10 ;
			data[8296] <= 8'h10 ;
			data[8297] <= 8'h10 ;
			data[8298] <= 8'h10 ;
			data[8299] <= 8'h10 ;
			data[8300] <= 8'h10 ;
			data[8301] <= 8'h10 ;
			data[8302] <= 8'h10 ;
			data[8303] <= 8'h10 ;
			data[8304] <= 8'h10 ;
			data[8305] <= 8'h10 ;
			data[8306] <= 8'h10 ;
			data[8307] <= 8'h10 ;
			data[8308] <= 8'h10 ;
			data[8309] <= 8'h10 ;
			data[8310] <= 8'h10 ;
			data[8311] <= 8'h10 ;
			data[8312] <= 8'h10 ;
			data[8313] <= 8'h10 ;
			data[8314] <= 8'h10 ;
			data[8315] <= 8'h10 ;
			data[8316] <= 8'h10 ;
			data[8317] <= 8'h10 ;
			data[8318] <= 8'h10 ;
			data[8319] <= 8'h10 ;
			data[8320] <= 8'h10 ;
			data[8321] <= 8'h10 ;
			data[8322] <= 8'h10 ;
			data[8323] <= 8'h10 ;
			data[8324] <= 8'h10 ;
			data[8325] <= 8'h10 ;
			data[8326] <= 8'h10 ;
			data[8327] <= 8'h10 ;
			data[8328] <= 8'h10 ;
			data[8329] <= 8'h10 ;
			data[8330] <= 8'h10 ;
			data[8331] <= 8'h10 ;
			data[8332] <= 8'h10 ;
			data[8333] <= 8'h10 ;
			data[8334] <= 8'h10 ;
			data[8335] <= 8'h10 ;
			data[8336] <= 8'h10 ;
			data[8337] <= 8'h10 ;
			data[8338] <= 8'h10 ;
			data[8339] <= 8'h10 ;
			data[8340] <= 8'h10 ;
			data[8341] <= 8'h10 ;
			data[8342] <= 8'h10 ;
			data[8343] <= 8'h10 ;
			data[8344] <= 8'h10 ;
			data[8345] <= 8'h10 ;
			data[8346] <= 8'h10 ;
			data[8347] <= 8'h10 ;
			data[8348] <= 8'h10 ;
			data[8349] <= 8'h10 ;
			data[8350] <= 8'h10 ;
			data[8351] <= 8'h10 ;
			data[8352] <= 8'h10 ;
			data[8353] <= 8'h10 ;
			data[8354] <= 8'h10 ;
			data[8355] <= 8'h10 ;
			data[8356] <= 8'h10 ;
			data[8357] <= 8'h10 ;
			data[8358] <= 8'h10 ;
			data[8359] <= 8'h10 ;
			data[8360] <= 8'h10 ;
			data[8361] <= 8'h10 ;
			data[8362] <= 8'h10 ;
			data[8363] <= 8'h10 ;
			data[8364] <= 8'h10 ;
			data[8365] <= 8'h10 ;
			data[8366] <= 8'h10 ;
			data[8367] <= 8'h10 ;
			data[8368] <= 8'h10 ;
			data[8369] <= 8'h10 ;
			data[8370] <= 8'h10 ;
			data[8371] <= 8'h10 ;
			data[8372] <= 8'h10 ;
			data[8373] <= 8'h10 ;
			data[8374] <= 8'h10 ;
			data[8375] <= 8'h10 ;
			data[8376] <= 8'h10 ;
			data[8377] <= 8'h10 ;
			data[8378] <= 8'h10 ;
			data[8379] <= 8'h10 ;
			data[8380] <= 8'h10 ;
			data[8381] <= 8'h10 ;
			data[8382] <= 8'h10 ;
			data[8383] <= 8'h10 ;
			data[8384] <= 8'h10 ;
			data[8385] <= 8'h10 ;
			data[8386] <= 8'h10 ;
			data[8387] <= 8'h10 ;
			data[8388] <= 8'h10 ;
			data[8389] <= 8'h10 ;
			data[8390] <= 8'h10 ;
			data[8391] <= 8'h10 ;
			data[8392] <= 8'h10 ;
			data[8393] <= 8'h10 ;
			data[8394] <= 8'h10 ;
			data[8395] <= 8'h10 ;
			data[8396] <= 8'h10 ;
			data[8397] <= 8'h10 ;
			data[8398] <= 8'h10 ;
			data[8399] <= 8'h10 ;
			data[8400] <= 8'h10 ;
			data[8401] <= 8'h10 ;
			data[8402] <= 8'h10 ;
			data[8403] <= 8'h10 ;
			data[8404] <= 8'h10 ;
			data[8405] <= 8'h10 ;
			data[8406] <= 8'h10 ;
			data[8407] <= 8'h10 ;
			data[8408] <= 8'h10 ;
			data[8409] <= 8'h10 ;
			data[8410] <= 8'h10 ;
			data[8411] <= 8'h10 ;
			data[8412] <= 8'h10 ;
			data[8413] <= 8'h10 ;
			data[8414] <= 8'h10 ;
			data[8415] <= 8'h10 ;
			data[8416] <= 8'h10 ;
			data[8417] <= 8'h10 ;
			data[8418] <= 8'h10 ;
			data[8419] <= 8'h10 ;
			data[8420] <= 8'h10 ;
			data[8421] <= 8'h10 ;
			data[8422] <= 8'h10 ;
			data[8423] <= 8'h10 ;
			data[8424] <= 8'h10 ;
			data[8425] <= 8'h10 ;
			data[8426] <= 8'h10 ;
			data[8427] <= 8'h10 ;
			data[8428] <= 8'h10 ;
			data[8429] <= 8'h10 ;
			data[8430] <= 8'h10 ;
			data[8431] <= 8'h10 ;
			data[8432] <= 8'h10 ;
			data[8433] <= 8'h10 ;
			data[8434] <= 8'h10 ;
			data[8435] <= 8'h10 ;
			data[8436] <= 8'h10 ;
			data[8437] <= 8'h10 ;
			data[8438] <= 8'h10 ;
			data[8439] <= 8'h10 ;
			data[8440] <= 8'h10 ;
			data[8441] <= 8'h10 ;
			data[8442] <= 8'h10 ;
			data[8443] <= 8'h10 ;
			data[8444] <= 8'h10 ;
			data[8445] <= 8'h10 ;
			data[8446] <= 8'h10 ;
			data[8447] <= 8'h10 ;
			data[8448] <= 8'h10 ;
			data[8449] <= 8'h10 ;
			data[8450] <= 8'h10 ;
			data[8451] <= 8'h10 ;
			data[8452] <= 8'h10 ;
			data[8453] <= 8'h10 ;
			data[8454] <= 8'h10 ;
			data[8455] <= 8'h10 ;
			data[8456] <= 8'h10 ;
			data[8457] <= 8'h10 ;
			data[8458] <= 8'h10 ;
			data[8459] <= 8'h10 ;
			data[8460] <= 8'h10 ;
			data[8461] <= 8'h10 ;
			data[8462] <= 8'h10 ;
			data[8463] <= 8'h10 ;
			data[8464] <= 8'h10 ;
			data[8465] <= 8'h10 ;
			data[8466] <= 8'h10 ;
			data[8467] <= 8'h10 ;
			data[8468] <= 8'h10 ;
			data[8469] <= 8'h10 ;
			data[8470] <= 8'h10 ;
			data[8471] <= 8'h10 ;
			data[8472] <= 8'h10 ;
			data[8473] <= 8'h10 ;
			data[8474] <= 8'h10 ;
			data[8475] <= 8'h10 ;
			data[8476] <= 8'h10 ;
			data[8477] <= 8'h10 ;
			data[8478] <= 8'h10 ;
			data[8479] <= 8'h10 ;
			data[8480] <= 8'h10 ;
			data[8481] <= 8'h10 ;
			data[8482] <= 8'h10 ;
			data[8483] <= 8'h10 ;
			data[8484] <= 8'h10 ;
			data[8485] <= 8'h10 ;
			data[8486] <= 8'h10 ;
			data[8487] <= 8'h10 ;
			data[8488] <= 8'h10 ;
			data[8489] <= 8'h10 ;
			data[8490] <= 8'h10 ;
			data[8491] <= 8'h10 ;
			data[8492] <= 8'h10 ;
			data[8493] <= 8'h10 ;
			data[8494] <= 8'h10 ;
			data[8495] <= 8'h10 ;
			data[8496] <= 8'h10 ;
			data[8497] <= 8'h10 ;
			data[8498] <= 8'h10 ;
			data[8499] <= 8'h10 ;
			data[8500] <= 8'h10 ;
			data[8501] <= 8'h10 ;
			data[8502] <= 8'h10 ;
			data[8503] <= 8'h10 ;
			data[8504] <= 8'h10 ;
			data[8505] <= 8'h10 ;
			data[8506] <= 8'h10 ;
			data[8507] <= 8'h10 ;
			data[8508] <= 8'h10 ;
			data[8509] <= 8'h10 ;
			data[8510] <= 8'h10 ;
			data[8511] <= 8'h10 ;
			data[8512] <= 8'h10 ;
			data[8513] <= 8'h10 ;
			data[8514] <= 8'h10 ;
			data[8515] <= 8'h10 ;
			data[8516] <= 8'h10 ;
			data[8517] <= 8'h10 ;
			data[8518] <= 8'h10 ;
			data[8519] <= 8'h10 ;
			data[8520] <= 8'h10 ;
			data[8521] <= 8'h10 ;
			data[8522] <= 8'h10 ;
			data[8523] <= 8'h10 ;
			data[8524] <= 8'h10 ;
			data[8525] <= 8'h10 ;
			data[8526] <= 8'h10 ;
			data[8527] <= 8'h10 ;
			data[8528] <= 8'h10 ;
			data[8529] <= 8'h10 ;
			data[8530] <= 8'h10 ;
			data[8531] <= 8'h10 ;
			data[8532] <= 8'h10 ;
			data[8533] <= 8'h10 ;
			data[8534] <= 8'h10 ;
			data[8535] <= 8'h10 ;
			data[8536] <= 8'h10 ;
			data[8537] <= 8'h10 ;
			data[8538] <= 8'h10 ;
			data[8539] <= 8'h10 ;
			data[8540] <= 8'h10 ;
			data[8541] <= 8'h10 ;
			data[8542] <= 8'h10 ;
			data[8543] <= 8'h10 ;
			data[8544] <= 8'h10 ;
			data[8545] <= 8'h10 ;
			data[8546] <= 8'h10 ;
			data[8547] <= 8'h10 ;
			data[8548] <= 8'h10 ;
			data[8549] <= 8'h10 ;
			data[8550] <= 8'h10 ;
			data[8551] <= 8'h10 ;
			data[8552] <= 8'h10 ;
			data[8553] <= 8'h10 ;
			data[8554] <= 8'h10 ;
			data[8555] <= 8'h10 ;
			data[8556] <= 8'h10 ;
			data[8557] <= 8'h10 ;
			data[8558] <= 8'h10 ;
			data[8559] <= 8'h10 ;
			data[8560] <= 8'h10 ;
			data[8561] <= 8'h10 ;
			data[8562] <= 8'h10 ;
			data[8563] <= 8'h10 ;
			data[8564] <= 8'h10 ;
			data[8565] <= 8'h10 ;
			data[8566] <= 8'h10 ;
			data[8567] <= 8'h10 ;
			data[8568] <= 8'h10 ;
			data[8569] <= 8'h10 ;
			data[8570] <= 8'h10 ;
			data[8571] <= 8'h10 ;
			data[8572] <= 8'h10 ;
			data[8573] <= 8'h10 ;
			data[8574] <= 8'h10 ;
			data[8575] <= 8'h10 ;
			data[8576] <= 8'h10 ;
			data[8577] <= 8'h10 ;
			data[8578] <= 8'h10 ;
			data[8579] <= 8'h10 ;
			data[8580] <= 8'h10 ;
			data[8581] <= 8'h10 ;
			data[8582] <= 8'h10 ;
			data[8583] <= 8'h10 ;
			data[8584] <= 8'h10 ;
			data[8585] <= 8'h10 ;
			data[8586] <= 8'h10 ;
			data[8587] <= 8'h10 ;
			data[8588] <= 8'h10 ;
			data[8589] <= 8'h10 ;
			data[8590] <= 8'h10 ;
			data[8591] <= 8'h10 ;
			data[8592] <= 8'h10 ;
			data[8593] <= 8'h10 ;
			data[8594] <= 8'h10 ;
			data[8595] <= 8'h10 ;
			data[8596] <= 8'h10 ;
			data[8597] <= 8'h10 ;
			data[8598] <= 8'h10 ;
			data[8599] <= 8'h10 ;
			data[8600] <= 8'h10 ;
			data[8601] <= 8'h10 ;
			data[8602] <= 8'h10 ;
			data[8603] <= 8'h10 ;
			data[8604] <= 8'h10 ;
			data[8605] <= 8'h10 ;
			data[8606] <= 8'h10 ;
			data[8607] <= 8'h10 ;
			data[8608] <= 8'h10 ;
			data[8609] <= 8'h10 ;
			data[8610] <= 8'h10 ;
			data[8611] <= 8'h10 ;
			data[8612] <= 8'h10 ;
			data[8613] <= 8'h10 ;
			data[8614] <= 8'h10 ;
			data[8615] <= 8'h10 ;
			data[8616] <= 8'h10 ;
			data[8617] <= 8'h10 ;
			data[8618] <= 8'h10 ;
			data[8619] <= 8'h10 ;
			data[8620] <= 8'h10 ;
			data[8621] <= 8'h10 ;
			data[8622] <= 8'h10 ;
			data[8623] <= 8'h10 ;
			data[8624] <= 8'h10 ;
			data[8625] <= 8'h10 ;
			data[8626] <= 8'h10 ;
			data[8627] <= 8'h10 ;
			data[8628] <= 8'h10 ;
			data[8629] <= 8'h10 ;
			data[8630] <= 8'h10 ;
			data[8631] <= 8'h10 ;
			data[8632] <= 8'h10 ;
			data[8633] <= 8'h10 ;
			data[8634] <= 8'h10 ;
			data[8635] <= 8'h10 ;
			data[8636] <= 8'h10 ;
			data[8637] <= 8'h10 ;
			data[8638] <= 8'h10 ;
			data[8639] <= 8'h10 ;
			data[8640] <= 8'h10 ;
			data[8641] <= 8'h10 ;
			data[8642] <= 8'h10 ;
			data[8643] <= 8'h10 ;
			data[8644] <= 8'h10 ;
			data[8645] <= 8'h10 ;
			data[8646] <= 8'h10 ;
			data[8647] <= 8'h10 ;
			data[8648] <= 8'h10 ;
			data[8649] <= 8'h10 ;
			data[8650] <= 8'h10 ;
			data[8651] <= 8'h10 ;
			data[8652] <= 8'h10 ;
			data[8653] <= 8'h10 ;
			data[8654] <= 8'h10 ;
			data[8655] <= 8'h10 ;
			data[8656] <= 8'h10 ;
			data[8657] <= 8'h10 ;
			data[8658] <= 8'h10 ;
			data[8659] <= 8'h10 ;
			data[8660] <= 8'h10 ;
			data[8661] <= 8'h10 ;
			data[8662] <= 8'h10 ;
			data[8663] <= 8'h10 ;
			data[8664] <= 8'h10 ;
			data[8665] <= 8'h10 ;
			data[8666] <= 8'h10 ;
			data[8667] <= 8'h10 ;
			data[8668] <= 8'h10 ;
			data[8669] <= 8'h10 ;
			data[8670] <= 8'h10 ;
			data[8671] <= 8'h10 ;
			data[8672] <= 8'h10 ;
			data[8673] <= 8'h10 ;
			data[8674] <= 8'h10 ;
			data[8675] <= 8'h10 ;
			data[8676] <= 8'h10 ;
			data[8677] <= 8'h10 ;
			data[8678] <= 8'h10 ;
			data[8679] <= 8'h10 ;
			data[8680] <= 8'h10 ;
			data[8681] <= 8'h10 ;
			data[8682] <= 8'h10 ;
			data[8683] <= 8'h10 ;
			data[8684] <= 8'h10 ;
			data[8685] <= 8'h10 ;
			data[8686] <= 8'h10 ;
			data[8687] <= 8'h10 ;
			data[8688] <= 8'h10 ;
			data[8689] <= 8'h10 ;
			data[8690] <= 8'h10 ;
			data[8691] <= 8'h10 ;
			data[8692] <= 8'h10 ;
			data[8693] <= 8'h10 ;
			data[8694] <= 8'h10 ;
			data[8695] <= 8'h10 ;
			data[8696] <= 8'h10 ;
			data[8697] <= 8'h10 ;
			data[8698] <= 8'h10 ;
			data[8699] <= 8'h10 ;
			data[8700] <= 8'h10 ;
			data[8701] <= 8'h10 ;
			data[8702] <= 8'h10 ;
			data[8703] <= 8'h10 ;
			data[8704] <= 8'h10 ;
			data[8705] <= 8'h10 ;
			data[8706] <= 8'h10 ;
			data[8707] <= 8'h10 ;
			data[8708] <= 8'h10 ;
			data[8709] <= 8'h10 ;
			data[8710] <= 8'h10 ;
			data[8711] <= 8'h10 ;
			data[8712] <= 8'h10 ;
			data[8713] <= 8'h10 ;
			data[8714] <= 8'h10 ;
			data[8715] <= 8'h10 ;
			data[8716] <= 8'h10 ;
			data[8717] <= 8'h10 ;
			data[8718] <= 8'h10 ;
			data[8719] <= 8'h10 ;
			data[8720] <= 8'h10 ;
			data[8721] <= 8'h10 ;
			data[8722] <= 8'h10 ;
			data[8723] <= 8'h10 ;
			data[8724] <= 8'h10 ;
			data[8725] <= 8'h10 ;
			data[8726] <= 8'h10 ;
			data[8727] <= 8'h10 ;
			data[8728] <= 8'h10 ;
			data[8729] <= 8'h10 ;
			data[8730] <= 8'h10 ;
			data[8731] <= 8'h10 ;
			data[8732] <= 8'h10 ;
			data[8733] <= 8'h10 ;
			data[8734] <= 8'h10 ;
			data[8735] <= 8'h10 ;
			data[8736] <= 8'h10 ;
			data[8737] <= 8'h10 ;
			data[8738] <= 8'h10 ;
			data[8739] <= 8'h10 ;
			data[8740] <= 8'h10 ;
			data[8741] <= 8'h10 ;
			data[8742] <= 8'h10 ;
			data[8743] <= 8'h10 ;
			data[8744] <= 8'h10 ;
			data[8745] <= 8'h10 ;
			data[8746] <= 8'h10 ;
			data[8747] <= 8'h10 ;
			data[8748] <= 8'h10 ;
			data[8749] <= 8'h10 ;
			data[8750] <= 8'h10 ;
			data[8751] <= 8'h10 ;
			data[8752] <= 8'h10 ;
			data[8753] <= 8'h10 ;
			data[8754] <= 8'h10 ;
			data[8755] <= 8'h10 ;
			data[8756] <= 8'h10 ;
			data[8757] <= 8'h10 ;
			data[8758] <= 8'h10 ;
			data[8759] <= 8'h10 ;
			data[8760] <= 8'h10 ;
			data[8761] <= 8'h10 ;
			data[8762] <= 8'h10 ;
			data[8763] <= 8'h10 ;
			data[8764] <= 8'h10 ;
			data[8765] <= 8'h10 ;
			data[8766] <= 8'h10 ;
			data[8767] <= 8'h10 ;
			data[8768] <= 8'h10 ;
			data[8769] <= 8'h10 ;
			data[8770] <= 8'h10 ;
			data[8771] <= 8'h10 ;
			data[8772] <= 8'h10 ;
			data[8773] <= 8'h10 ;
			data[8774] <= 8'h10 ;
			data[8775] <= 8'h10 ;
			data[8776] <= 8'h10 ;
			data[8777] <= 8'h10 ;
			data[8778] <= 8'h10 ;
			data[8779] <= 8'h10 ;
			data[8780] <= 8'h10 ;
			data[8781] <= 8'h10 ;
			data[8782] <= 8'h10 ;
			data[8783] <= 8'h10 ;
			data[8784] <= 8'h10 ;
			data[8785] <= 8'h10 ;
			data[8786] <= 8'h10 ;
			data[8787] <= 8'h10 ;
			data[8788] <= 8'h10 ;
			data[8789] <= 8'h10 ;
			data[8790] <= 8'h10 ;
			data[8791] <= 8'h10 ;
			data[8792] <= 8'h10 ;
			data[8793] <= 8'h10 ;
			data[8794] <= 8'h10 ;
			data[8795] <= 8'h10 ;
			data[8796] <= 8'h10 ;
			data[8797] <= 8'h10 ;
			data[8798] <= 8'h10 ;
			data[8799] <= 8'h10 ;
			data[8800] <= 8'h10 ;
			data[8801] <= 8'h10 ;
			data[8802] <= 8'h10 ;
			data[8803] <= 8'h10 ;
			data[8804] <= 8'h10 ;
			data[8805] <= 8'h10 ;
			data[8806] <= 8'h10 ;
			data[8807] <= 8'h10 ;
			data[8808] <= 8'h10 ;
			data[8809] <= 8'h10 ;
			data[8810] <= 8'h10 ;
			data[8811] <= 8'h10 ;
			data[8812] <= 8'h10 ;
			data[8813] <= 8'h10 ;
			data[8814] <= 8'h10 ;
			data[8815] <= 8'h10 ;
			data[8816] <= 8'h10 ;
			data[8817] <= 8'h10 ;
			data[8818] <= 8'h10 ;
			data[8819] <= 8'h10 ;
			data[8820] <= 8'h10 ;
			data[8821] <= 8'h10 ;
			data[8822] <= 8'h10 ;
			data[8823] <= 8'h10 ;
			data[8824] <= 8'h10 ;
			data[8825] <= 8'h10 ;
			data[8826] <= 8'h10 ;
			data[8827] <= 8'h10 ;
			data[8828] <= 8'h10 ;
			data[8829] <= 8'h10 ;
			data[8830] <= 8'h10 ;
			data[8831] <= 8'h10 ;
			data[8832] <= 8'h10 ;
			data[8833] <= 8'h10 ;
			data[8834] <= 8'h10 ;
			data[8835] <= 8'h10 ;
			data[8836] <= 8'h10 ;
			data[8837] <= 8'h10 ;
			data[8838] <= 8'h10 ;
			data[8839] <= 8'h10 ;
			data[8840] <= 8'h10 ;
			data[8841] <= 8'h10 ;
			data[8842] <= 8'h10 ;
			data[8843] <= 8'h10 ;
			data[8844] <= 8'h10 ;
			data[8845] <= 8'h10 ;
			data[8846] <= 8'h10 ;
			data[8847] <= 8'h10 ;
			data[8848] <= 8'h10 ;
			data[8849] <= 8'h10 ;
			data[8850] <= 8'h10 ;
			data[8851] <= 8'h10 ;
			data[8852] <= 8'h10 ;
			data[8853] <= 8'h10 ;
			data[8854] <= 8'h10 ;
			data[8855] <= 8'h10 ;
			data[8856] <= 8'h10 ;
			data[8857] <= 8'h10 ;
			data[8858] <= 8'h10 ;
			data[8859] <= 8'h10 ;
			data[8860] <= 8'h10 ;
			data[8861] <= 8'h10 ;
			data[8862] <= 8'h10 ;
			data[8863] <= 8'h10 ;
			data[8864] <= 8'h10 ;
			data[8865] <= 8'h10 ;
			data[8866] <= 8'h10 ;
			data[8867] <= 8'h10 ;
			data[8868] <= 8'h10 ;
			data[8869] <= 8'h10 ;
			data[8870] <= 8'h10 ;
			data[8871] <= 8'h10 ;
			data[8872] <= 8'h10 ;
			data[8873] <= 8'h10 ;
			data[8874] <= 8'h10 ;
			data[8875] <= 8'h10 ;
			data[8876] <= 8'h10 ;
			data[8877] <= 8'h10 ;
			data[8878] <= 8'h10 ;
			data[8879] <= 8'h10 ;
			data[8880] <= 8'h10 ;
			data[8881] <= 8'h10 ;
			data[8882] <= 8'h10 ;
			data[8883] <= 8'h10 ;
			data[8884] <= 8'h10 ;
			data[8885] <= 8'h10 ;
			data[8886] <= 8'h10 ;
			data[8887] <= 8'h10 ;
			data[8888] <= 8'h10 ;
			data[8889] <= 8'h10 ;
			data[8890] <= 8'h10 ;
			data[8891] <= 8'h10 ;
			data[8892] <= 8'h10 ;
			data[8893] <= 8'h10 ;
			data[8894] <= 8'h10 ;
			data[8895] <= 8'h10 ;
			data[8896] <= 8'h10 ;
			data[8897] <= 8'h10 ;
			data[8898] <= 8'h10 ;
			data[8899] <= 8'h10 ;
			data[8900] <= 8'h10 ;
			data[8901] <= 8'h10 ;
			data[8902] <= 8'h10 ;
			data[8903] <= 8'h10 ;
			data[8904] <= 8'h10 ;
			data[8905] <= 8'h10 ;
			data[8906] <= 8'h10 ;
			data[8907] <= 8'h10 ;
			data[8908] <= 8'h10 ;
			data[8909] <= 8'h10 ;
			data[8910] <= 8'h10 ;
			data[8911] <= 8'h10 ;
			data[8912] <= 8'h10 ;
			data[8913] <= 8'h10 ;
			data[8914] <= 8'h10 ;
			data[8915] <= 8'h10 ;
			data[8916] <= 8'h10 ;
			data[8917] <= 8'h10 ;
			data[8918] <= 8'h10 ;
			data[8919] <= 8'h10 ;
			data[8920] <= 8'h10 ;
			data[8921] <= 8'h10 ;
			data[8922] <= 8'h10 ;
			data[8923] <= 8'h10 ;
			data[8924] <= 8'h10 ;
			data[8925] <= 8'h10 ;
			data[8926] <= 8'h10 ;
			data[8927] <= 8'h10 ;
			data[8928] <= 8'h10 ;
			data[8929] <= 8'h10 ;
			data[8930] <= 8'h10 ;
			data[8931] <= 8'h10 ;
			data[8932] <= 8'h10 ;
			data[8933] <= 8'h10 ;
			data[8934] <= 8'h10 ;
			data[8935] <= 8'h10 ;
			data[8936] <= 8'h10 ;
			data[8937] <= 8'h10 ;
			data[8938] <= 8'h10 ;
			data[8939] <= 8'h10 ;
			data[8940] <= 8'h10 ;
			data[8941] <= 8'h10 ;
			data[8942] <= 8'h10 ;
			data[8943] <= 8'h10 ;
			data[8944] <= 8'h10 ;
			data[8945] <= 8'h10 ;
			data[8946] <= 8'h10 ;
			data[8947] <= 8'h10 ;
			data[8948] <= 8'h10 ;
			data[8949] <= 8'h10 ;
			data[8950] <= 8'h10 ;
			data[8951] <= 8'h10 ;
			data[8952] <= 8'h10 ;
			data[8953] <= 8'h10 ;
			data[8954] <= 8'h10 ;
			data[8955] <= 8'h10 ;
			data[8956] <= 8'h10 ;
			data[8957] <= 8'h10 ;
			data[8958] <= 8'h10 ;
			data[8959] <= 8'h10 ;
			data[8960] <= 8'h10 ;
			data[8961] <= 8'h10 ;
			data[8962] <= 8'h10 ;
			data[8963] <= 8'h10 ;
			data[8964] <= 8'h10 ;
			data[8965] <= 8'h10 ;
			data[8966] <= 8'h10 ;
			data[8967] <= 8'h10 ;
			data[8968] <= 8'h10 ;
			data[8969] <= 8'h10 ;
			data[8970] <= 8'h10 ;
			data[8971] <= 8'h10 ;
			data[8972] <= 8'h10 ;
			data[8973] <= 8'h10 ;
			data[8974] <= 8'h10 ;
			data[8975] <= 8'h10 ;
			data[8976] <= 8'h10 ;
			data[8977] <= 8'h10 ;
			data[8978] <= 8'h10 ;
			data[8979] <= 8'h10 ;
			data[8980] <= 8'h10 ;
			data[8981] <= 8'h10 ;
			data[8982] <= 8'h10 ;
			data[8983] <= 8'h10 ;
			data[8984] <= 8'h10 ;
			data[8985] <= 8'h10 ;
			data[8986] <= 8'h10 ;
			data[8987] <= 8'h10 ;
			data[8988] <= 8'h10 ;
			data[8989] <= 8'h10 ;
			data[8990] <= 8'h10 ;
			data[8991] <= 8'h10 ;
			data[8992] <= 8'h10 ;
			data[8993] <= 8'h10 ;
			data[8994] <= 8'h10 ;
			data[8995] <= 8'h10 ;
			data[8996] <= 8'h10 ;
			data[8997] <= 8'h10 ;
			data[8998] <= 8'h10 ;
			data[8999] <= 8'h10 ;
			data[9000] <= 8'h10 ;
			data[9001] <= 8'h10 ;
			data[9002] <= 8'h10 ;
			data[9003] <= 8'h10 ;
			data[9004] <= 8'h10 ;
			data[9005] <= 8'h10 ;
			data[9006] <= 8'h10 ;
			data[9007] <= 8'h10 ;
			data[9008] <= 8'h10 ;
			data[9009] <= 8'h10 ;
			data[9010] <= 8'h10 ;
			data[9011] <= 8'h10 ;
			data[9012] <= 8'h10 ;
			data[9013] <= 8'h10 ;
			data[9014] <= 8'h10 ;
			data[9015] <= 8'h10 ;
			data[9016] <= 8'h10 ;
			data[9017] <= 8'h10 ;
			data[9018] <= 8'h10 ;
			data[9019] <= 8'h10 ;
			data[9020] <= 8'h10 ;
			data[9021] <= 8'h10 ;
			data[9022] <= 8'h10 ;
			data[9023] <= 8'h10 ;
			data[9024] <= 8'h10 ;
			data[9025] <= 8'h10 ;
			data[9026] <= 8'h10 ;
			data[9027] <= 8'h10 ;
			data[9028] <= 8'h10 ;
			data[9029] <= 8'h10 ;
			data[9030] <= 8'h10 ;
			data[9031] <= 8'h10 ;
			data[9032] <= 8'h10 ;
			data[9033] <= 8'h10 ;
			data[9034] <= 8'h10 ;
			data[9035] <= 8'h10 ;
			data[9036] <= 8'h10 ;
			data[9037] <= 8'h10 ;
			data[9038] <= 8'h10 ;
			data[9039] <= 8'h10 ;
			data[9040] <= 8'h10 ;
			data[9041] <= 8'h10 ;
			data[9042] <= 8'h10 ;
			data[9043] <= 8'h10 ;
			data[9044] <= 8'h10 ;
			data[9045] <= 8'h10 ;
			data[9046] <= 8'h10 ;
			data[9047] <= 8'h10 ;
			data[9048] <= 8'h10 ;
			data[9049] <= 8'h10 ;
			data[9050] <= 8'h10 ;
			data[9051] <= 8'h10 ;
			data[9052] <= 8'h10 ;
			data[9053] <= 8'h10 ;
			data[9054] <= 8'h10 ;
			data[9055] <= 8'h10 ;
			data[9056] <= 8'h10 ;
			data[9057] <= 8'h10 ;
			data[9058] <= 8'h10 ;
			data[9059] <= 8'h10 ;
			data[9060] <= 8'h10 ;
			data[9061] <= 8'h10 ;
			data[9062] <= 8'h10 ;
			data[9063] <= 8'h10 ;
			data[9064] <= 8'h10 ;
			data[9065] <= 8'h10 ;
			data[9066] <= 8'h10 ;
			data[9067] <= 8'h10 ;
			data[9068] <= 8'h10 ;
			data[9069] <= 8'h10 ;
			data[9070] <= 8'h10 ;
			data[9071] <= 8'h10 ;
			data[9072] <= 8'h10 ;
			data[9073] <= 8'h10 ;
			data[9074] <= 8'h10 ;
			data[9075] <= 8'h10 ;
			data[9076] <= 8'h10 ;
			data[9077] <= 8'h10 ;
			data[9078] <= 8'h10 ;
			data[9079] <= 8'h10 ;
			data[9080] <= 8'h10 ;
			data[9081] <= 8'h10 ;
			data[9082] <= 8'h10 ;
			data[9083] <= 8'h10 ;
			data[9084] <= 8'h10 ;
			data[9085] <= 8'h10 ;
			data[9086] <= 8'h10 ;
			data[9087] <= 8'h10 ;
			data[9088] <= 8'h10 ;
			data[9089] <= 8'h10 ;
			data[9090] <= 8'h10 ;
			data[9091] <= 8'h10 ;
			data[9092] <= 8'h10 ;
			data[9093] <= 8'h10 ;
			data[9094] <= 8'h10 ;
			data[9095] <= 8'h10 ;
			data[9096] <= 8'h10 ;
			data[9097] <= 8'h10 ;
			data[9098] <= 8'h10 ;
			data[9099] <= 8'h10 ;
			data[9100] <= 8'h10 ;
			data[9101] <= 8'h10 ;
			data[9102] <= 8'h10 ;
			data[9103] <= 8'h10 ;
			data[9104] <= 8'h10 ;
			data[9105] <= 8'h10 ;
			data[9106] <= 8'h10 ;
			data[9107] <= 8'h10 ;
			data[9108] <= 8'h10 ;
			data[9109] <= 8'h10 ;
			data[9110] <= 8'h10 ;
			data[9111] <= 8'h10 ;
			data[9112] <= 8'h10 ;
			data[9113] <= 8'h10 ;
			data[9114] <= 8'h10 ;
			data[9115] <= 8'h10 ;
			data[9116] <= 8'h10 ;
			data[9117] <= 8'h10 ;
			data[9118] <= 8'h10 ;
			data[9119] <= 8'h10 ;
			data[9120] <= 8'h10 ;
			data[9121] <= 8'h10 ;
			data[9122] <= 8'h10 ;
			data[9123] <= 8'h10 ;
			data[9124] <= 8'h10 ;
			data[9125] <= 8'h10 ;
			data[9126] <= 8'h10 ;
			data[9127] <= 8'h10 ;
			data[9128] <= 8'h10 ;
			data[9129] <= 8'h10 ;
			data[9130] <= 8'h10 ;
			data[9131] <= 8'h10 ;
			data[9132] <= 8'h10 ;
			data[9133] <= 8'h10 ;
			data[9134] <= 8'h10 ;
			data[9135] <= 8'h10 ;
			data[9136] <= 8'h10 ;
			data[9137] <= 8'h10 ;
			data[9138] <= 8'h10 ;
			data[9139] <= 8'h10 ;
			data[9140] <= 8'h10 ;
			data[9141] <= 8'h10 ;
			data[9142] <= 8'h10 ;
			data[9143] <= 8'h10 ;
			data[9144] <= 8'h10 ;
			data[9145] <= 8'h10 ;
			data[9146] <= 8'h10 ;
			data[9147] <= 8'h10 ;
			data[9148] <= 8'h10 ;
			data[9149] <= 8'h10 ;
			data[9150] <= 8'h10 ;
			data[9151] <= 8'h10 ;
			data[9152] <= 8'h10 ;
			data[9153] <= 8'h10 ;
			data[9154] <= 8'h10 ;
			data[9155] <= 8'h10 ;
			data[9156] <= 8'h10 ;
			data[9157] <= 8'h10 ;
			data[9158] <= 8'h10 ;
			data[9159] <= 8'h10 ;
			data[9160] <= 8'h10 ;
			data[9161] <= 8'h10 ;
			data[9162] <= 8'h10 ;
			data[9163] <= 8'h10 ;
			data[9164] <= 8'h10 ;
			data[9165] <= 8'h10 ;
			data[9166] <= 8'h10 ;
			data[9167] <= 8'h10 ;
			data[9168] <= 8'h10 ;
			data[9169] <= 8'h10 ;
			data[9170] <= 8'h10 ;
			data[9171] <= 8'h10 ;
			data[9172] <= 8'h10 ;
			data[9173] <= 8'h10 ;
			data[9174] <= 8'h10 ;
			data[9175] <= 8'h10 ;
			data[9176] <= 8'h10 ;
			data[9177] <= 8'h10 ;
			data[9178] <= 8'h10 ;
			data[9179] <= 8'h10 ;
			data[9180] <= 8'h10 ;
			data[9181] <= 8'h10 ;
			data[9182] <= 8'h10 ;
			data[9183] <= 8'h10 ;
			data[9184] <= 8'h10 ;
			data[9185] <= 8'h10 ;
			data[9186] <= 8'h10 ;
			data[9187] <= 8'h10 ;
			data[9188] <= 8'h10 ;
			data[9189] <= 8'h10 ;
			data[9190] <= 8'h10 ;
			data[9191] <= 8'h10 ;
			data[9192] <= 8'h10 ;
			data[9193] <= 8'h10 ;
			data[9194] <= 8'h10 ;
			data[9195] <= 8'h10 ;
			data[9196] <= 8'h10 ;
			data[9197] <= 8'h10 ;
			data[9198] <= 8'h10 ;
			data[9199] <= 8'h10 ;
			data[9200] <= 8'h10 ;
			data[9201] <= 8'h10 ;
			data[9202] <= 8'h10 ;
			data[9203] <= 8'h10 ;
			data[9204] <= 8'h10 ;
			data[9205] <= 8'h10 ;
			data[9206] <= 8'h10 ;
			data[9207] <= 8'h10 ;
			data[9208] <= 8'h10 ;
			data[9209] <= 8'h10 ;
			data[9210] <= 8'h10 ;
			data[9211] <= 8'h10 ;
			data[9212] <= 8'h10 ;
			data[9213] <= 8'h10 ;
			data[9214] <= 8'h10 ;
			data[9215] <= 8'h10 ;
			data[9216] <= 8'h10 ;
			data[9217] <= 8'h10 ;
			data[9218] <= 8'h10 ;
			data[9219] <= 8'h10 ;
			data[9220] <= 8'h10 ;
			data[9221] <= 8'h10 ;
			data[9222] <= 8'h10 ;
			data[9223] <= 8'h10 ;
			data[9224] <= 8'h10 ;
			data[9225] <= 8'h10 ;
			data[9226] <= 8'h10 ;
			data[9227] <= 8'h10 ;
			data[9228] <= 8'h10 ;
			data[9229] <= 8'h10 ;
			data[9230] <= 8'h10 ;
			data[9231] <= 8'h10 ;
			data[9232] <= 8'h10 ;
			data[9233] <= 8'h10 ;
			data[9234] <= 8'h10 ;
			data[9235] <= 8'h10 ;
			data[9236] <= 8'h10 ;
			data[9237] <= 8'h10 ;
			data[9238] <= 8'h10 ;
			data[9239] <= 8'h10 ;
			data[9240] <= 8'h10 ;
			data[9241] <= 8'h10 ;
			data[9242] <= 8'h10 ;
			data[9243] <= 8'h10 ;
			data[9244] <= 8'h10 ;
			data[9245] <= 8'h10 ;
			data[9246] <= 8'h10 ;
			data[9247] <= 8'h10 ;
			data[9248] <= 8'h10 ;
			data[9249] <= 8'h10 ;
			data[9250] <= 8'h10 ;
			data[9251] <= 8'h10 ;
			data[9252] <= 8'h10 ;
			data[9253] <= 8'h10 ;
			data[9254] <= 8'h10 ;
			data[9255] <= 8'h10 ;
			data[9256] <= 8'h10 ;
			data[9257] <= 8'h10 ;
			data[9258] <= 8'h10 ;
			data[9259] <= 8'h10 ;
			data[9260] <= 8'h10 ;
			data[9261] <= 8'h10 ;
			data[9262] <= 8'h10 ;
			data[9263] <= 8'h10 ;
			data[9264] <= 8'h10 ;
			data[9265] <= 8'h10 ;
			data[9266] <= 8'h10 ;
			data[9267] <= 8'h10 ;
			data[9268] <= 8'h10 ;
			data[9269] <= 8'h10 ;
			data[9270] <= 8'h10 ;
			data[9271] <= 8'h10 ;
			data[9272] <= 8'h10 ;
			data[9273] <= 8'h10 ;
			data[9274] <= 8'h10 ;
			data[9275] <= 8'h10 ;
			data[9276] <= 8'h10 ;
			data[9277] <= 8'h10 ;
			data[9278] <= 8'h10 ;
			data[9279] <= 8'h10 ;
			data[9280] <= 8'h10 ;
			data[9281] <= 8'h10 ;
			data[9282] <= 8'h10 ;
			data[9283] <= 8'h10 ;
			data[9284] <= 8'h10 ;
			data[9285] <= 8'h10 ;
			data[9286] <= 8'h10 ;
			data[9287] <= 8'h10 ;
			data[9288] <= 8'h10 ;
			data[9289] <= 8'h10 ;
			data[9290] <= 8'h10 ;
			data[9291] <= 8'h10 ;
			data[9292] <= 8'h10 ;
			data[9293] <= 8'h10 ;
			data[9294] <= 8'h10 ;
			data[9295] <= 8'h10 ;
			data[9296] <= 8'h10 ;
			data[9297] <= 8'h10 ;
			data[9298] <= 8'h10 ;
			data[9299] <= 8'h10 ;
			data[9300] <= 8'h10 ;
			data[9301] <= 8'h10 ;
			data[9302] <= 8'h10 ;
			data[9303] <= 8'h10 ;
			data[9304] <= 8'h10 ;
			data[9305] <= 8'h10 ;
			data[9306] <= 8'h10 ;
			data[9307] <= 8'h10 ;
			data[9308] <= 8'h10 ;
			data[9309] <= 8'h10 ;
			data[9310] <= 8'h10 ;
			data[9311] <= 8'h10 ;
			data[9312] <= 8'h10 ;
			data[9313] <= 8'h10 ;
			data[9314] <= 8'h10 ;
			data[9315] <= 8'h10 ;
			data[9316] <= 8'h10 ;
			data[9317] <= 8'h10 ;
			data[9318] <= 8'h10 ;
			data[9319] <= 8'h10 ;
			data[9320] <= 8'h10 ;
			data[9321] <= 8'h10 ;
			data[9322] <= 8'h10 ;
			data[9323] <= 8'h10 ;
			data[9324] <= 8'h10 ;
			data[9325] <= 8'h10 ;
			data[9326] <= 8'h10 ;
			data[9327] <= 8'h10 ;
			data[9328] <= 8'h10 ;
			data[9329] <= 8'h10 ;
			data[9330] <= 8'h10 ;
			data[9331] <= 8'h10 ;
			data[9332] <= 8'h10 ;
			data[9333] <= 8'h10 ;
			data[9334] <= 8'h10 ;
			data[9335] <= 8'h10 ;
			data[9336] <= 8'h10 ;
			data[9337] <= 8'h10 ;
			data[9338] <= 8'h10 ;
			data[9339] <= 8'h10 ;
			data[9340] <= 8'h10 ;
			data[9341] <= 8'h10 ;
			data[9342] <= 8'h10 ;
			data[9343] <= 8'h10 ;
			data[9344] <= 8'h10 ;
			data[9345] <= 8'h10 ;
			data[9346] <= 8'h10 ;
			data[9347] <= 8'h10 ;
			data[9348] <= 8'h10 ;
			data[9349] <= 8'h10 ;
			data[9350] <= 8'h10 ;
			data[9351] <= 8'h10 ;
			data[9352] <= 8'h10 ;
			data[9353] <= 8'h10 ;
			data[9354] <= 8'h10 ;
			data[9355] <= 8'h10 ;
			data[9356] <= 8'h10 ;
			data[9357] <= 8'h10 ;
			data[9358] <= 8'h10 ;
			data[9359] <= 8'h10 ;
			data[9360] <= 8'h10 ;
			data[9361] <= 8'h10 ;
			data[9362] <= 8'h10 ;
			data[9363] <= 8'h10 ;
			data[9364] <= 8'h10 ;
			data[9365] <= 8'h10 ;
			data[9366] <= 8'h10 ;
			data[9367] <= 8'h10 ;
			data[9368] <= 8'h10 ;
			data[9369] <= 8'h10 ;
			data[9370] <= 8'h10 ;
			data[9371] <= 8'h10 ;
			data[9372] <= 8'h10 ;
			data[9373] <= 8'h10 ;
			data[9374] <= 8'h10 ;
			data[9375] <= 8'h10 ;
			data[9376] <= 8'h10 ;
			data[9377] <= 8'h10 ;
			data[9378] <= 8'h10 ;
			data[9379] <= 8'h10 ;
			data[9380] <= 8'h10 ;
			data[9381] <= 8'h10 ;
			data[9382] <= 8'h10 ;
			data[9383] <= 8'h10 ;
			data[9384] <= 8'h10 ;
			data[9385] <= 8'h10 ;
			data[9386] <= 8'h10 ;
			data[9387] <= 8'h10 ;
			data[9388] <= 8'h10 ;
			data[9389] <= 8'h10 ;
			data[9390] <= 8'h10 ;
			data[9391] <= 8'h10 ;
			data[9392] <= 8'h10 ;
			data[9393] <= 8'h10 ;
			data[9394] <= 8'h10 ;
			data[9395] <= 8'h10 ;
			data[9396] <= 8'h10 ;
			data[9397] <= 8'h10 ;
			data[9398] <= 8'h10 ;
			data[9399] <= 8'h10 ;
			data[9400] <= 8'h10 ;
			data[9401] <= 8'h10 ;
			data[9402] <= 8'h10 ;
			data[9403] <= 8'h10 ;
			data[9404] <= 8'h10 ;
			data[9405] <= 8'h10 ;
			data[9406] <= 8'h10 ;
			data[9407] <= 8'h10 ;
			data[9408] <= 8'h10 ;
			data[9409] <= 8'h10 ;
			data[9410] <= 8'h10 ;
			data[9411] <= 8'h10 ;
			data[9412] <= 8'h10 ;
			data[9413] <= 8'h10 ;
			data[9414] <= 8'h10 ;
			data[9415] <= 8'h10 ;
			data[9416] <= 8'h10 ;
			data[9417] <= 8'h10 ;
			data[9418] <= 8'h10 ;
			data[9419] <= 8'h10 ;
			data[9420] <= 8'h10 ;
			data[9421] <= 8'h10 ;
			data[9422] <= 8'h10 ;
			data[9423] <= 8'h10 ;
			data[9424] <= 8'h10 ;
			data[9425] <= 8'h10 ;
			data[9426] <= 8'h10 ;
			data[9427] <= 8'h10 ;
			data[9428] <= 8'h10 ;
			data[9429] <= 8'h10 ;
			data[9430] <= 8'h10 ;
			data[9431] <= 8'h10 ;
			data[9432] <= 8'h10 ;
			data[9433] <= 8'h10 ;
			data[9434] <= 8'h10 ;
			data[9435] <= 8'h10 ;
			data[9436] <= 8'h10 ;
			data[9437] <= 8'h10 ;
			data[9438] <= 8'h10 ;
			data[9439] <= 8'h10 ;
			data[9440] <= 8'h10 ;
			data[9441] <= 8'h10 ;
			data[9442] <= 8'h10 ;
			data[9443] <= 8'h10 ;
			data[9444] <= 8'h10 ;
			data[9445] <= 8'h10 ;
			data[9446] <= 8'h10 ;
			data[9447] <= 8'h10 ;
			data[9448] <= 8'h10 ;
			data[9449] <= 8'h10 ;
			data[9450] <= 8'h10 ;
			data[9451] <= 8'h10 ;
			data[9452] <= 8'h10 ;
			data[9453] <= 8'h10 ;
			data[9454] <= 8'h10 ;
			data[9455] <= 8'h10 ;
			data[9456] <= 8'h10 ;
			data[9457] <= 8'h10 ;
			data[9458] <= 8'h10 ;
			data[9459] <= 8'h10 ;
			data[9460] <= 8'h10 ;
			data[9461] <= 8'h10 ;
			data[9462] <= 8'h10 ;
			data[9463] <= 8'h10 ;
			data[9464] <= 8'h10 ;
			data[9465] <= 8'h10 ;
			data[9466] <= 8'h10 ;
			data[9467] <= 8'h10 ;
			data[9468] <= 8'h10 ;
			data[9469] <= 8'h10 ;
			data[9470] <= 8'h10 ;
			data[9471] <= 8'h10 ;
			data[9472] <= 8'h10 ;
			data[9473] <= 8'h10 ;
			data[9474] <= 8'h10 ;
			data[9475] <= 8'h10 ;
			data[9476] <= 8'h10 ;
			data[9477] <= 8'h10 ;
			data[9478] <= 8'h10 ;
			data[9479] <= 8'h10 ;
			data[9480] <= 8'h10 ;
			data[9481] <= 8'h10 ;
			data[9482] <= 8'h10 ;
			data[9483] <= 8'h10 ;
			data[9484] <= 8'h10 ;
			data[9485] <= 8'h10 ;
			data[9486] <= 8'h10 ;
			data[9487] <= 8'h10 ;
			data[9488] <= 8'h10 ;
			data[9489] <= 8'h10 ;
			data[9490] <= 8'h10 ;
			data[9491] <= 8'h10 ;
			data[9492] <= 8'h10 ;
			data[9493] <= 8'h10 ;
			data[9494] <= 8'h10 ;
			data[9495] <= 8'h10 ;
			data[9496] <= 8'h10 ;
			data[9497] <= 8'h10 ;
			data[9498] <= 8'h10 ;
			data[9499] <= 8'h10 ;
			data[9500] <= 8'h10 ;
			data[9501] <= 8'h10 ;
			data[9502] <= 8'h10 ;
			data[9503] <= 8'h10 ;
			data[9504] <= 8'h10 ;
			data[9505] <= 8'h10 ;
			data[9506] <= 8'h10 ;
			data[9507] <= 8'h10 ;
			data[9508] <= 8'h10 ;
			data[9509] <= 8'h10 ;
			data[9510] <= 8'h10 ;
			data[9511] <= 8'h10 ;
			data[9512] <= 8'h10 ;
			data[9513] <= 8'h10 ;
			data[9514] <= 8'h10 ;
			data[9515] <= 8'h10 ;
			data[9516] <= 8'h10 ;
			data[9517] <= 8'h10 ;
			data[9518] <= 8'h10 ;
			data[9519] <= 8'h10 ;
			data[9520] <= 8'h10 ;
			data[9521] <= 8'h10 ;
			data[9522] <= 8'h10 ;
			data[9523] <= 8'h10 ;
			data[9524] <= 8'h10 ;
			data[9525] <= 8'h10 ;
			data[9526] <= 8'h10 ;
			data[9527] <= 8'h10 ;
			data[9528] <= 8'h10 ;
			data[9529] <= 8'h10 ;
			data[9530] <= 8'h10 ;
			data[9531] <= 8'h10 ;
			data[9532] <= 8'h10 ;
			data[9533] <= 8'h10 ;
			data[9534] <= 8'h10 ;
			data[9535] <= 8'h10 ;
			data[9536] <= 8'h10 ;
			data[9537] <= 8'h10 ;
			data[9538] <= 8'h10 ;
			data[9539] <= 8'h10 ;
			data[9540] <= 8'h10 ;
			data[9541] <= 8'h10 ;
			data[9542] <= 8'h10 ;
			data[9543] <= 8'h10 ;
			data[9544] <= 8'h10 ;
			data[9545] <= 8'h10 ;
			data[9546] <= 8'h10 ;
			data[9547] <= 8'h10 ;
			data[9548] <= 8'h10 ;
			data[9549] <= 8'h10 ;
			data[9550] <= 8'h10 ;
			data[9551] <= 8'h10 ;
			data[9552] <= 8'h10 ;
			data[9553] <= 8'h10 ;
			data[9554] <= 8'h10 ;
			data[9555] <= 8'h10 ;
			data[9556] <= 8'h10 ;
			data[9557] <= 8'h10 ;
			data[9558] <= 8'h10 ;
			data[9559] <= 8'h10 ;
			data[9560] <= 8'h10 ;
			data[9561] <= 8'h10 ;
			data[9562] <= 8'h10 ;
			data[9563] <= 8'h10 ;
			data[9564] <= 8'h10 ;
			data[9565] <= 8'h10 ;
			data[9566] <= 8'h10 ;
			data[9567] <= 8'h10 ;
			data[9568] <= 8'h10 ;
			data[9569] <= 8'h10 ;
			data[9570] <= 8'h10 ;
			data[9571] <= 8'h10 ;
			data[9572] <= 8'h10 ;
			data[9573] <= 8'h10 ;
			data[9574] <= 8'h10 ;
			data[9575] <= 8'h10 ;
			data[9576] <= 8'h10 ;
			data[9577] <= 8'h10 ;
			data[9578] <= 8'h10 ;
			data[9579] <= 8'h10 ;
			data[9580] <= 8'h10 ;
			data[9581] <= 8'h10 ;
			data[9582] <= 8'h10 ;
			data[9583] <= 8'h10 ;
			data[9584] <= 8'h10 ;
			data[9585] <= 8'h10 ;
			data[9586] <= 8'h10 ;
			data[9587] <= 8'h10 ;
			data[9588] <= 8'h10 ;
			data[9589] <= 8'h10 ;
			data[9590] <= 8'h10 ;
			data[9591] <= 8'h10 ;
			data[9592] <= 8'h10 ;
			data[9593] <= 8'h10 ;
			data[9594] <= 8'h10 ;
			data[9595] <= 8'h10 ;
			data[9596] <= 8'h10 ;
			data[9597] <= 8'h10 ;
			data[9598] <= 8'h10 ;
			data[9599] <= 8'h10 ;
			data[9600] <= 8'h10 ;
			data[9601] <= 8'h10 ;
			data[9602] <= 8'h10 ;
			data[9603] <= 8'h10 ;
			data[9604] <= 8'h10 ;
			data[9605] <= 8'h10 ;
			data[9606] <= 8'h10 ;
			data[9607] <= 8'h10 ;
			data[9608] <= 8'h10 ;
			data[9609] <= 8'h10 ;
			data[9610] <= 8'h10 ;
			data[9611] <= 8'h10 ;
			data[9612] <= 8'h10 ;
			data[9613] <= 8'h10 ;
			data[9614] <= 8'h10 ;
			data[9615] <= 8'h10 ;
			data[9616] <= 8'h10 ;
			data[9617] <= 8'h10 ;
			data[9618] <= 8'h10 ;
			data[9619] <= 8'h10 ;
			data[9620] <= 8'h10 ;
			data[9621] <= 8'h10 ;
			data[9622] <= 8'h10 ;
			data[9623] <= 8'h10 ;
			data[9624] <= 8'h10 ;
			data[9625] <= 8'h10 ;
			data[9626] <= 8'h10 ;
			data[9627] <= 8'h10 ;
			data[9628] <= 8'h10 ;
			data[9629] <= 8'h10 ;
			data[9630] <= 8'h10 ;
			data[9631] <= 8'h10 ;
			data[9632] <= 8'h10 ;
			data[9633] <= 8'h10 ;
			data[9634] <= 8'h10 ;
			data[9635] <= 8'h10 ;
			data[9636] <= 8'h10 ;
			data[9637] <= 8'h10 ;
			data[9638] <= 8'h10 ;
			data[9639] <= 8'h10 ;
			data[9640] <= 8'h10 ;
			data[9641] <= 8'h10 ;
			data[9642] <= 8'h10 ;
			data[9643] <= 8'h10 ;
			data[9644] <= 8'h10 ;
			data[9645] <= 8'h10 ;
			data[9646] <= 8'h10 ;
			data[9647] <= 8'h10 ;
			data[9648] <= 8'h10 ;
			data[9649] <= 8'h10 ;
			data[9650] <= 8'h10 ;
			data[9651] <= 8'h10 ;
			data[9652] <= 8'h10 ;
			data[9653] <= 8'h10 ;
			data[9654] <= 8'h10 ;
			data[9655] <= 8'h10 ;
			data[9656] <= 8'h10 ;
			data[9657] <= 8'h10 ;
			data[9658] <= 8'h10 ;
			data[9659] <= 8'h10 ;
			data[9660] <= 8'h10 ;
			data[9661] <= 8'h10 ;
			data[9662] <= 8'h10 ;
			data[9663] <= 8'h10 ;
			data[9664] <= 8'h10 ;
			data[9665] <= 8'h10 ;
			data[9666] <= 8'h10 ;
			data[9667] <= 8'h10 ;
			data[9668] <= 8'h10 ;
			data[9669] <= 8'h10 ;
			data[9670] <= 8'h10 ;
			data[9671] <= 8'h10 ;
			data[9672] <= 8'h10 ;
			data[9673] <= 8'h10 ;
			data[9674] <= 8'h10 ;
			data[9675] <= 8'h10 ;
			data[9676] <= 8'h10 ;
			data[9677] <= 8'h10 ;
			data[9678] <= 8'h10 ;
			data[9679] <= 8'h10 ;
			data[9680] <= 8'h10 ;
			data[9681] <= 8'h10 ;
			data[9682] <= 8'h10 ;
			data[9683] <= 8'h10 ;
			data[9684] <= 8'h10 ;
			data[9685] <= 8'h10 ;
			data[9686] <= 8'h10 ;
			data[9687] <= 8'h10 ;
			data[9688] <= 8'h10 ;
			data[9689] <= 8'h10 ;
			data[9690] <= 8'h10 ;
			data[9691] <= 8'h10 ;
			data[9692] <= 8'h10 ;
			data[9693] <= 8'h10 ;
			data[9694] <= 8'h10 ;
			data[9695] <= 8'h10 ;
			data[9696] <= 8'h10 ;
			data[9697] <= 8'h10 ;
			data[9698] <= 8'h10 ;
			data[9699] <= 8'h10 ;
			data[9700] <= 8'h10 ;
			data[9701] <= 8'h10 ;
			data[9702] <= 8'h10 ;
			data[9703] <= 8'h10 ;
			data[9704] <= 8'h10 ;
			data[9705] <= 8'h10 ;
			data[9706] <= 8'h10 ;
			data[9707] <= 8'h10 ;
			data[9708] <= 8'h10 ;
			data[9709] <= 8'h10 ;
			data[9710] <= 8'h10 ;
			data[9711] <= 8'h10 ;
			data[9712] <= 8'h10 ;
			data[9713] <= 8'h10 ;
			data[9714] <= 8'h10 ;
			data[9715] <= 8'h10 ;
			data[9716] <= 8'h10 ;
			data[9717] <= 8'h10 ;
			data[9718] <= 8'h10 ;
			data[9719] <= 8'h10 ;
			data[9720] <= 8'h10 ;
			data[9721] <= 8'h10 ;
			data[9722] <= 8'h10 ;
			data[9723] <= 8'h10 ;
			data[9724] <= 8'h10 ;
			data[9725] <= 8'h10 ;
			data[9726] <= 8'h10 ;
			data[9727] <= 8'h10 ;
			data[9728] <= 8'h10 ;
			data[9729] <= 8'h10 ;
			data[9730] <= 8'h10 ;
			data[9731] <= 8'h10 ;
			data[9732] <= 8'h10 ;
			data[9733] <= 8'h10 ;
			data[9734] <= 8'h10 ;
			data[9735] <= 8'h10 ;
			data[9736] <= 8'h10 ;
			data[9737] <= 8'h10 ;
			data[9738] <= 8'h10 ;
			data[9739] <= 8'h10 ;
			data[9740] <= 8'h10 ;
			data[9741] <= 8'h10 ;
			data[9742] <= 8'h10 ;
			data[9743] <= 8'h10 ;
			data[9744] <= 8'h10 ;
			data[9745] <= 8'h10 ;
			data[9746] <= 8'h10 ;
			data[9747] <= 8'h10 ;
			data[9748] <= 8'h10 ;
			data[9749] <= 8'h10 ;
			data[9750] <= 8'h10 ;
			data[9751] <= 8'h10 ;
			data[9752] <= 8'h10 ;
			data[9753] <= 8'h10 ;
			data[9754] <= 8'h10 ;
			data[9755] <= 8'h10 ;
			data[9756] <= 8'h10 ;
			data[9757] <= 8'h10 ;
			data[9758] <= 8'h10 ;
			data[9759] <= 8'h10 ;
			data[9760] <= 8'h10 ;
			data[9761] <= 8'h10 ;
			data[9762] <= 8'h10 ;
			data[9763] <= 8'h10 ;
			data[9764] <= 8'h10 ;
			data[9765] <= 8'h10 ;
			data[9766] <= 8'h10 ;
			data[9767] <= 8'h10 ;
			data[9768] <= 8'h10 ;
			data[9769] <= 8'h10 ;
			data[9770] <= 8'h10 ;
			data[9771] <= 8'h10 ;
			data[9772] <= 8'h10 ;
			data[9773] <= 8'h10 ;
			data[9774] <= 8'h10 ;
			data[9775] <= 8'h10 ;
			data[9776] <= 8'h10 ;
			data[9777] <= 8'h10 ;
			data[9778] <= 8'h10 ;
			data[9779] <= 8'h10 ;
			data[9780] <= 8'h10 ;
			data[9781] <= 8'h10 ;
			data[9782] <= 8'h10 ;
			data[9783] <= 8'h10 ;
			data[9784] <= 8'h10 ;
			data[9785] <= 8'h10 ;
			data[9786] <= 8'h10 ;
			data[9787] <= 8'h10 ;
			data[9788] <= 8'h10 ;
			data[9789] <= 8'h10 ;
			data[9790] <= 8'h10 ;
			data[9791] <= 8'h10 ;
			data[9792] <= 8'h10 ;
			data[9793] <= 8'h10 ;
			data[9794] <= 8'h10 ;
			data[9795] <= 8'h10 ;
			data[9796] <= 8'h10 ;
			data[9797] <= 8'h10 ;
			data[9798] <= 8'h10 ;
			data[9799] <= 8'h10 ;
			data[9800] <= 8'h10 ;
			data[9801] <= 8'h10 ;
			data[9802] <= 8'h10 ;
			data[9803] <= 8'h10 ;
			data[9804] <= 8'h10 ;
			data[9805] <= 8'h10 ;
			data[9806] <= 8'h10 ;
			data[9807] <= 8'h10 ;
			data[9808] <= 8'h10 ;
			data[9809] <= 8'h10 ;
			data[9810] <= 8'h10 ;
			data[9811] <= 8'h10 ;
			data[9812] <= 8'h10 ;
			data[9813] <= 8'h10 ;
			data[9814] <= 8'h10 ;
			data[9815] <= 8'h10 ;
			data[9816] <= 8'h10 ;
			data[9817] <= 8'h10 ;
			data[9818] <= 8'h10 ;
			data[9819] <= 8'h10 ;
			data[9820] <= 8'h10 ;
			data[9821] <= 8'h10 ;
			data[9822] <= 8'h10 ;
			data[9823] <= 8'h10 ;
			data[9824] <= 8'h10 ;
			data[9825] <= 8'h10 ;
			data[9826] <= 8'h10 ;
			data[9827] <= 8'h10 ;
			data[9828] <= 8'h10 ;
			data[9829] <= 8'h10 ;
			data[9830] <= 8'h10 ;
			data[9831] <= 8'h10 ;
			data[9832] <= 8'h10 ;
			data[9833] <= 8'h10 ;
			data[9834] <= 8'h10 ;
			data[9835] <= 8'h10 ;
			data[9836] <= 8'h10 ;
			data[9837] <= 8'h10 ;
			data[9838] <= 8'h10 ;
			data[9839] <= 8'h10 ;
			data[9840] <= 8'h10 ;
			data[9841] <= 8'h10 ;
			data[9842] <= 8'h10 ;
			data[9843] <= 8'h10 ;
			data[9844] <= 8'h10 ;
			data[9845] <= 8'h10 ;
			data[9846] <= 8'h10 ;
			data[9847] <= 8'h10 ;
			data[9848] <= 8'h10 ;
			data[9849] <= 8'h10 ;
			data[9850] <= 8'h10 ;
			data[9851] <= 8'h10 ;
			data[9852] <= 8'h10 ;
			data[9853] <= 8'h10 ;
			data[9854] <= 8'h10 ;
			data[9855] <= 8'h10 ;
			data[9856] <= 8'h10 ;
			data[9857] <= 8'h10 ;
			data[9858] <= 8'h10 ;
			data[9859] <= 8'h10 ;
			data[9860] <= 8'h10 ;
			data[9861] <= 8'h10 ;
			data[9862] <= 8'h10 ;
			data[9863] <= 8'h10 ;
			data[9864] <= 8'h10 ;
			data[9865] <= 8'h10 ;
			data[9866] <= 8'h10 ;
			data[9867] <= 8'h10 ;
			data[9868] <= 8'h10 ;
			data[9869] <= 8'h10 ;
			data[9870] <= 8'h10 ;
			data[9871] <= 8'h10 ;
			data[9872] <= 8'h10 ;
			data[9873] <= 8'h10 ;
			data[9874] <= 8'h10 ;
			data[9875] <= 8'h10 ;
			data[9876] <= 8'h10 ;
			data[9877] <= 8'h10 ;
			data[9878] <= 8'h10 ;
			data[9879] <= 8'h10 ;
			data[9880] <= 8'h10 ;
			data[9881] <= 8'h10 ;
			data[9882] <= 8'h10 ;
			data[9883] <= 8'h10 ;
			data[9884] <= 8'h10 ;
			data[9885] <= 8'h10 ;
			data[9886] <= 8'h10 ;
			data[9887] <= 8'h10 ;
			data[9888] <= 8'h10 ;
			data[9889] <= 8'h10 ;
			data[9890] <= 8'h10 ;
			data[9891] <= 8'h10 ;
			data[9892] <= 8'h10 ;
			data[9893] <= 8'h10 ;
			data[9894] <= 8'h10 ;
			data[9895] <= 8'h10 ;
			data[9896] <= 8'h10 ;
			data[9897] <= 8'h10 ;
			data[9898] <= 8'h10 ;
			data[9899] <= 8'h10 ;
			data[9900] <= 8'h10 ;
			data[9901] <= 8'h10 ;
			data[9902] <= 8'h10 ;
			data[9903] <= 8'h10 ;
			data[9904] <= 8'h10 ;
			data[9905] <= 8'h10 ;
			data[9906] <= 8'h10 ;
			data[9907] <= 8'h10 ;
			data[9908] <= 8'h10 ;
			data[9909] <= 8'h10 ;
			data[9910] <= 8'h10 ;
			data[9911] <= 8'h10 ;
			data[9912] <= 8'h10 ;
			data[9913] <= 8'h10 ;
			data[9914] <= 8'h10 ;
			data[9915] <= 8'h10 ;
			data[9916] <= 8'h10 ;
			data[9917] <= 8'h10 ;
			data[9918] <= 8'h10 ;
			data[9919] <= 8'h10 ;
			data[9920] <= 8'h10 ;
			data[9921] <= 8'h10 ;
			data[9922] <= 8'h10 ;
			data[9923] <= 8'h10 ;
			data[9924] <= 8'h10 ;
			data[9925] <= 8'h10 ;
			data[9926] <= 8'h10 ;
			data[9927] <= 8'h10 ;
			data[9928] <= 8'h10 ;
			data[9929] <= 8'h10 ;
			data[9930] <= 8'h10 ;
			data[9931] <= 8'h10 ;
			data[9932] <= 8'h10 ;
			data[9933] <= 8'h10 ;
			data[9934] <= 8'h10 ;
			data[9935] <= 8'h10 ;
			data[9936] <= 8'h10 ;
			data[9937] <= 8'h10 ;
			data[9938] <= 8'h10 ;
			data[9939] <= 8'h10 ;
			data[9940] <= 8'h10 ;
			data[9941] <= 8'h10 ;
			data[9942] <= 8'h10 ;
			data[9943] <= 8'h10 ;
			data[9944] <= 8'h10 ;
			data[9945] <= 8'h10 ;
			data[9946] <= 8'h10 ;
			data[9947] <= 8'h10 ;
			data[9948] <= 8'h10 ;
			data[9949] <= 8'h10 ;
			data[9950] <= 8'h10 ;
			data[9951] <= 8'h10 ;
			data[9952] <= 8'h10 ;
			data[9953] <= 8'h10 ;
			data[9954] <= 8'h10 ;
			data[9955] <= 8'h10 ;
			data[9956] <= 8'h10 ;
			data[9957] <= 8'h10 ;
			data[9958] <= 8'h10 ;
			data[9959] <= 8'h10 ;
			data[9960] <= 8'h10 ;
			data[9961] <= 8'h10 ;
			data[9962] <= 8'h10 ;
			data[9963] <= 8'h10 ;
			data[9964] <= 8'h10 ;
			data[9965] <= 8'h10 ;
			data[9966] <= 8'h10 ;
			data[9967] <= 8'h10 ;
			data[9968] <= 8'h10 ;
			data[9969] <= 8'h10 ;
			data[9970] <= 8'h10 ;
			data[9971] <= 8'h10 ;
			data[9972] <= 8'h10 ;
			data[9973] <= 8'h10 ;
			data[9974] <= 8'h10 ;
			data[9975] <= 8'h10 ;
			data[9976] <= 8'h10 ;
			data[9977] <= 8'h10 ;
			data[9978] <= 8'h10 ;
			data[9979] <= 8'h10 ;
			data[9980] <= 8'h10 ;
			data[9981] <= 8'h10 ;
			data[9982] <= 8'h10 ;
			data[9983] <= 8'h10 ;
			data[9984] <= 8'h10 ;
			data[9985] <= 8'h10 ;
			data[9986] <= 8'h10 ;
			data[9987] <= 8'h10 ;
			data[9988] <= 8'h10 ;
			data[9989] <= 8'h10 ;
			data[9990] <= 8'h10 ;
			data[9991] <= 8'h10 ;
			data[9992] <= 8'h10 ;
			data[9993] <= 8'h10 ;
			data[9994] <= 8'h10 ;
			data[9995] <= 8'h10 ;
			data[9996] <= 8'h10 ;
			data[9997] <= 8'h10 ;
			data[9998] <= 8'h10 ;
			data[9999] <= 8'h10 ;
			data[10000] <= 8'h10 ;
			data[10001] <= 8'h10 ;
			data[10002] <= 8'h10 ;
			data[10003] <= 8'h10 ;
			data[10004] <= 8'h10 ;
			data[10005] <= 8'h10 ;
			data[10006] <= 8'h10 ;
			data[10007] <= 8'h10 ;
			data[10008] <= 8'h10 ;
			data[10009] <= 8'h10 ;
			data[10010] <= 8'h10 ;
			data[10011] <= 8'h10 ;
			data[10012] <= 8'h10 ;
			data[10013] <= 8'h10 ;
			data[10014] <= 8'h10 ;
			data[10015] <= 8'h10 ;
			data[10016] <= 8'h10 ;
			data[10017] <= 8'h10 ;
			data[10018] <= 8'h10 ;
			data[10019] <= 8'h10 ;
			data[10020] <= 8'h10 ;
			data[10021] <= 8'h10 ;
			data[10022] <= 8'h10 ;
			data[10023] <= 8'h10 ;
			data[10024] <= 8'h10 ;
			data[10025] <= 8'h10 ;
			data[10026] <= 8'h10 ;
			data[10027] <= 8'h10 ;
			data[10028] <= 8'h10 ;
			data[10029] <= 8'h10 ;
			data[10030] <= 8'h10 ;
			data[10031] <= 8'h10 ;
			data[10032] <= 8'h10 ;
			data[10033] <= 8'h10 ;
			data[10034] <= 8'h10 ;
			data[10035] <= 8'h10 ;
			data[10036] <= 8'h10 ;
			data[10037] <= 8'h10 ;
			data[10038] <= 8'h10 ;
			data[10039] <= 8'h10 ;
			data[10040] <= 8'h10 ;
			data[10041] <= 8'h10 ;
			data[10042] <= 8'h10 ;
			data[10043] <= 8'h10 ;
			data[10044] <= 8'h10 ;
			data[10045] <= 8'h10 ;
			data[10046] <= 8'h10 ;
			data[10047] <= 8'h10 ;
			data[10048] <= 8'h10 ;
			data[10049] <= 8'h10 ;
			data[10050] <= 8'h10 ;
			data[10051] <= 8'h10 ;
			data[10052] <= 8'h10 ;
			data[10053] <= 8'h10 ;
			data[10054] <= 8'h10 ;
			data[10055] <= 8'h10 ;
			data[10056] <= 8'h10 ;
			data[10057] <= 8'h10 ;
			data[10058] <= 8'h10 ;
			data[10059] <= 8'h10 ;
			data[10060] <= 8'h10 ;
			data[10061] <= 8'h10 ;
			data[10062] <= 8'h10 ;
			data[10063] <= 8'h10 ;
			data[10064] <= 8'h10 ;
			data[10065] <= 8'h10 ;
			data[10066] <= 8'h10 ;
			data[10067] <= 8'h10 ;
			data[10068] <= 8'h10 ;
			data[10069] <= 8'h10 ;
			data[10070] <= 8'h10 ;
			data[10071] <= 8'h10 ;
			data[10072] <= 8'h10 ;
			data[10073] <= 8'h10 ;
			data[10074] <= 8'h10 ;
			data[10075] <= 8'h10 ;
			data[10076] <= 8'h10 ;
			data[10077] <= 8'h10 ;
			data[10078] <= 8'h10 ;
			data[10079] <= 8'h10 ;
			data[10080] <= 8'h10 ;
			data[10081] <= 8'h10 ;
			data[10082] <= 8'h10 ;
			data[10083] <= 8'h10 ;
			data[10084] <= 8'h10 ;
			data[10085] <= 8'h10 ;
			data[10086] <= 8'h10 ;
			data[10087] <= 8'h10 ;
			data[10088] <= 8'h10 ;
			data[10089] <= 8'h10 ;
			data[10090] <= 8'h10 ;
			data[10091] <= 8'h10 ;
			data[10092] <= 8'h10 ;
			data[10093] <= 8'h10 ;
			data[10094] <= 8'h10 ;
			data[10095] <= 8'h10 ;
			data[10096] <= 8'h10 ;
			data[10097] <= 8'h10 ;
			data[10098] <= 8'h10 ;
			data[10099] <= 8'h10 ;
			data[10100] <= 8'h10 ;
			data[10101] <= 8'h10 ;
			data[10102] <= 8'h10 ;
			data[10103] <= 8'h10 ;
			data[10104] <= 8'h10 ;
			data[10105] <= 8'h10 ;
			data[10106] <= 8'h10 ;
			data[10107] <= 8'h10 ;
			data[10108] <= 8'h10 ;
			data[10109] <= 8'h10 ;
			data[10110] <= 8'h10 ;
			data[10111] <= 8'h10 ;
			data[10112] <= 8'h10 ;
			data[10113] <= 8'h10 ;
			data[10114] <= 8'h10 ;
			data[10115] <= 8'h10 ;
			data[10116] <= 8'h10 ;
			data[10117] <= 8'h10 ;
			data[10118] <= 8'h10 ;
			data[10119] <= 8'h10 ;
			data[10120] <= 8'h10 ;
			data[10121] <= 8'h10 ;
			data[10122] <= 8'h10 ;
			data[10123] <= 8'h10 ;
			data[10124] <= 8'h10 ;
			data[10125] <= 8'h10 ;
			data[10126] <= 8'h10 ;
			data[10127] <= 8'h10 ;
			data[10128] <= 8'h10 ;
			data[10129] <= 8'h10 ;
			data[10130] <= 8'h10 ;
			data[10131] <= 8'h10 ;
			data[10132] <= 8'h10 ;
			data[10133] <= 8'h10 ;
			data[10134] <= 8'h10 ;
			data[10135] <= 8'h10 ;
			data[10136] <= 8'h10 ;
			data[10137] <= 8'h10 ;
			data[10138] <= 8'h10 ;
			data[10139] <= 8'h10 ;
			data[10140] <= 8'h10 ;
			data[10141] <= 8'h10 ;
			data[10142] <= 8'h10 ;
			data[10143] <= 8'h10 ;
			data[10144] <= 8'h10 ;
			data[10145] <= 8'h10 ;
			data[10146] <= 8'h10 ;
			data[10147] <= 8'h10 ;
			data[10148] <= 8'h10 ;
			data[10149] <= 8'h10 ;
			data[10150] <= 8'h10 ;
			data[10151] <= 8'h10 ;
			data[10152] <= 8'h10 ;
			data[10153] <= 8'h10 ;
			data[10154] <= 8'h10 ;
			data[10155] <= 8'h10 ;
			data[10156] <= 8'h10 ;
			data[10157] <= 8'h10 ;
			data[10158] <= 8'h10 ;
			data[10159] <= 8'h10 ;
			data[10160] <= 8'h10 ;
			data[10161] <= 8'h10 ;
			data[10162] <= 8'h10 ;
			data[10163] <= 8'h10 ;
			data[10164] <= 8'h10 ;
			data[10165] <= 8'h10 ;
			data[10166] <= 8'h10 ;
			data[10167] <= 8'h10 ;
			data[10168] <= 8'h10 ;
			data[10169] <= 8'h10 ;
			data[10170] <= 8'h10 ;
			data[10171] <= 8'h10 ;
			data[10172] <= 8'h10 ;
			data[10173] <= 8'h10 ;
			data[10174] <= 8'h10 ;
			data[10175] <= 8'h10 ;
			data[10176] <= 8'h10 ;
			data[10177] <= 8'h10 ;
			data[10178] <= 8'h10 ;
			data[10179] <= 8'h10 ;
			data[10180] <= 8'h10 ;
			data[10181] <= 8'h10 ;
			data[10182] <= 8'h10 ;
			data[10183] <= 8'h10 ;
			data[10184] <= 8'h10 ;
			data[10185] <= 8'h10 ;
			data[10186] <= 8'h10 ;
			data[10187] <= 8'h10 ;
			data[10188] <= 8'h10 ;
			data[10189] <= 8'h10 ;
			data[10190] <= 8'h10 ;
			data[10191] <= 8'h10 ;
			data[10192] <= 8'h10 ;
			data[10193] <= 8'h10 ;
			data[10194] <= 8'h10 ;
			data[10195] <= 8'h10 ;
			data[10196] <= 8'h10 ;
			data[10197] <= 8'h10 ;
			data[10198] <= 8'h10 ;
			data[10199] <= 8'h10 ;
			data[10200] <= 8'h10 ;
			data[10201] <= 8'h10 ;
			data[10202] <= 8'h10 ;
			data[10203] <= 8'h10 ;
			data[10204] <= 8'h10 ;
			data[10205] <= 8'h10 ;
			data[10206] <= 8'h10 ;
			data[10207] <= 8'h10 ;
			data[10208] <= 8'h10 ;
			data[10209] <= 8'h10 ;
			data[10210] <= 8'h10 ;
			data[10211] <= 8'h10 ;
			data[10212] <= 8'h10 ;
			data[10213] <= 8'h10 ;
			data[10214] <= 8'h10 ;
			data[10215] <= 8'h10 ;
			data[10216] <= 8'h10 ;
			data[10217] <= 8'h10 ;
			data[10218] <= 8'h10 ;
			data[10219] <= 8'h10 ;
			data[10220] <= 8'h10 ;
			data[10221] <= 8'h10 ;
			data[10222] <= 8'h10 ;
			data[10223] <= 8'h10 ;
			data[10224] <= 8'h10 ;
			data[10225] <= 8'h10 ;
			data[10226] <= 8'h10 ;
			data[10227] <= 8'h10 ;
			data[10228] <= 8'h10 ;
			data[10229] <= 8'h10 ;
			data[10230] <= 8'h10 ;
			data[10231] <= 8'h10 ;
			data[10232] <= 8'h10 ;
			data[10233] <= 8'h10 ;
			data[10234] <= 8'h10 ;
			data[10235] <= 8'h10 ;
			data[10236] <= 8'h10 ;
			data[10237] <= 8'h10 ;
			data[10238] <= 8'h10 ;
			data[10239] <= 8'h10 ;
			data[10240] <= 8'h10 ;
			data[10241] <= 8'h10 ;
			data[10242] <= 8'h10 ;
			data[10243] <= 8'h10 ;
			data[10244] <= 8'h10 ;
			data[10245] <= 8'h10 ;
			data[10246] <= 8'h10 ;
			data[10247] <= 8'h10 ;
			data[10248] <= 8'h10 ;
			data[10249] <= 8'h10 ;
			data[10250] <= 8'h10 ;
			data[10251] <= 8'h10 ;
			data[10252] <= 8'h10 ;
			data[10253] <= 8'h10 ;
			data[10254] <= 8'h10 ;
			data[10255] <= 8'h10 ;
			data[10256] <= 8'h10 ;
			data[10257] <= 8'h10 ;
			data[10258] <= 8'h10 ;
			data[10259] <= 8'h10 ;
			data[10260] <= 8'h10 ;
			data[10261] <= 8'h10 ;
			data[10262] <= 8'h10 ;
			data[10263] <= 8'h10 ;
			data[10264] <= 8'h10 ;
			data[10265] <= 8'h10 ;
			data[10266] <= 8'h10 ;
			data[10267] <= 8'h10 ;
			data[10268] <= 8'h10 ;
			data[10269] <= 8'h10 ;
			data[10270] <= 8'h10 ;
			data[10271] <= 8'h10 ;
			data[10272] <= 8'h10 ;
			data[10273] <= 8'h10 ;
			data[10274] <= 8'h10 ;
			data[10275] <= 8'h10 ;
			data[10276] <= 8'h10 ;
			data[10277] <= 8'h10 ;
			data[10278] <= 8'h10 ;
			data[10279] <= 8'h10 ;
			data[10280] <= 8'h10 ;
			data[10281] <= 8'h10 ;
			data[10282] <= 8'h10 ;
			data[10283] <= 8'h10 ;
			data[10284] <= 8'h10 ;
			data[10285] <= 8'h10 ;
			data[10286] <= 8'h10 ;
			data[10287] <= 8'h10 ;
			data[10288] <= 8'h10 ;
			data[10289] <= 8'h10 ;
			data[10290] <= 8'h10 ;
			data[10291] <= 8'h10 ;
			data[10292] <= 8'h10 ;
			data[10293] <= 8'h10 ;
			data[10294] <= 8'h10 ;
			data[10295] <= 8'h10 ;
			data[10296] <= 8'h10 ;
			data[10297] <= 8'h10 ;
			data[10298] <= 8'h10 ;
			data[10299] <= 8'h10 ;
			data[10300] <= 8'h10 ;
			data[10301] <= 8'h10 ;
			data[10302] <= 8'h10 ;
			data[10303] <= 8'h10 ;
			data[10304] <= 8'h10 ;
			data[10305] <= 8'h10 ;
			data[10306] <= 8'h10 ;
			data[10307] <= 8'h10 ;
			data[10308] <= 8'h10 ;
			data[10309] <= 8'h10 ;
			data[10310] <= 8'h10 ;
			data[10311] <= 8'h10 ;
			data[10312] <= 8'h10 ;
			data[10313] <= 8'h10 ;
			data[10314] <= 8'h10 ;
			data[10315] <= 8'h10 ;
			data[10316] <= 8'h10 ;
			data[10317] <= 8'h10 ;
			data[10318] <= 8'h10 ;
			data[10319] <= 8'h10 ;
			data[10320] <= 8'h10 ;
			data[10321] <= 8'h10 ;
			data[10322] <= 8'h10 ;
			data[10323] <= 8'h10 ;
			data[10324] <= 8'h10 ;
			data[10325] <= 8'h10 ;
			data[10326] <= 8'h10 ;
			data[10327] <= 8'h10 ;
			data[10328] <= 8'h10 ;
			data[10329] <= 8'h10 ;
			data[10330] <= 8'h10 ;
			data[10331] <= 8'h10 ;
			data[10332] <= 8'h10 ;
			data[10333] <= 8'h10 ;
			data[10334] <= 8'h10 ;
			data[10335] <= 8'h10 ;
			data[10336] <= 8'h10 ;
			data[10337] <= 8'h10 ;
			data[10338] <= 8'h10 ;
			data[10339] <= 8'h10 ;
			data[10340] <= 8'h10 ;
			data[10341] <= 8'h10 ;
			data[10342] <= 8'h10 ;
			data[10343] <= 8'h10 ;
			data[10344] <= 8'h10 ;
			data[10345] <= 8'h10 ;
			data[10346] <= 8'h10 ;
			data[10347] <= 8'h10 ;
			data[10348] <= 8'h10 ;
			data[10349] <= 8'h10 ;
			data[10350] <= 8'h10 ;
			data[10351] <= 8'h10 ;
			data[10352] <= 8'h10 ;
			data[10353] <= 8'h10 ;
			data[10354] <= 8'h10 ;
			data[10355] <= 8'h10 ;
			data[10356] <= 8'h10 ;
			data[10357] <= 8'h10 ;
			data[10358] <= 8'h10 ;
			data[10359] <= 8'h10 ;
			data[10360] <= 8'h10 ;
			data[10361] <= 8'h10 ;
			data[10362] <= 8'h10 ;
			data[10363] <= 8'h10 ;
			data[10364] <= 8'h10 ;
			data[10365] <= 8'h10 ;
			data[10366] <= 8'h10 ;
			data[10367] <= 8'h10 ;
			data[10368] <= 8'h10 ;
			data[10369] <= 8'h10 ;
			data[10370] <= 8'h10 ;
			data[10371] <= 8'h10 ;
			data[10372] <= 8'h10 ;
			data[10373] <= 8'h10 ;
			data[10374] <= 8'h10 ;
			data[10375] <= 8'h10 ;
			data[10376] <= 8'h10 ;
			data[10377] <= 8'h10 ;
			data[10378] <= 8'h10 ;
			data[10379] <= 8'h10 ;
			data[10380] <= 8'h10 ;
			data[10381] <= 8'h10 ;
			data[10382] <= 8'h10 ;
			data[10383] <= 8'h10 ;
			data[10384] <= 8'h10 ;
			data[10385] <= 8'h10 ;
			data[10386] <= 8'h10 ;
			data[10387] <= 8'h10 ;
			data[10388] <= 8'h10 ;
			data[10389] <= 8'h10 ;
			data[10390] <= 8'h10 ;
			data[10391] <= 8'h10 ;
			data[10392] <= 8'h10 ;
			data[10393] <= 8'h10 ;
			data[10394] <= 8'h10 ;
			data[10395] <= 8'h10 ;
			data[10396] <= 8'h10 ;
			data[10397] <= 8'h10 ;
			data[10398] <= 8'h10 ;
			data[10399] <= 8'h10 ;
			data[10400] <= 8'h10 ;
			data[10401] <= 8'h10 ;
			data[10402] <= 8'h10 ;
			data[10403] <= 8'h10 ;
			data[10404] <= 8'h10 ;
			data[10405] <= 8'h10 ;
			data[10406] <= 8'h10 ;
			data[10407] <= 8'h10 ;
			data[10408] <= 8'h10 ;
			data[10409] <= 8'h10 ;
			data[10410] <= 8'h10 ;
			data[10411] <= 8'h10 ;
			data[10412] <= 8'h10 ;
			data[10413] <= 8'h10 ;
			data[10414] <= 8'h10 ;
			data[10415] <= 8'h10 ;
			data[10416] <= 8'h10 ;
			data[10417] <= 8'h10 ;
			data[10418] <= 8'h10 ;
			data[10419] <= 8'h10 ;
			data[10420] <= 8'h10 ;
			data[10421] <= 8'h10 ;
			data[10422] <= 8'h10 ;
			data[10423] <= 8'h10 ;
			data[10424] <= 8'h10 ;
			data[10425] <= 8'h10 ;
			data[10426] <= 8'h10 ;
			data[10427] <= 8'h10 ;
			data[10428] <= 8'h10 ;
			data[10429] <= 8'h10 ;
			data[10430] <= 8'h10 ;
			data[10431] <= 8'h10 ;
			data[10432] <= 8'h10 ;
			data[10433] <= 8'h10 ;
			data[10434] <= 8'h10 ;
			data[10435] <= 8'h10 ;
			data[10436] <= 8'h10 ;
			data[10437] <= 8'h10 ;
			data[10438] <= 8'h10 ;
			data[10439] <= 8'h10 ;
			data[10440] <= 8'h10 ;
			data[10441] <= 8'h10 ;
			data[10442] <= 8'h10 ;
			data[10443] <= 8'h10 ;
			data[10444] <= 8'h10 ;
			data[10445] <= 8'h10 ;
			data[10446] <= 8'h10 ;
			data[10447] <= 8'h10 ;
			data[10448] <= 8'h10 ;
			data[10449] <= 8'h10 ;
			data[10450] <= 8'h10 ;
			data[10451] <= 8'h10 ;
			data[10452] <= 8'h10 ;
			data[10453] <= 8'h10 ;
			data[10454] <= 8'h10 ;
			data[10455] <= 8'h10 ;
			data[10456] <= 8'h10 ;
			data[10457] <= 8'h10 ;
			data[10458] <= 8'h10 ;
			data[10459] <= 8'h10 ;
			data[10460] <= 8'h10 ;
			data[10461] <= 8'h10 ;
			data[10462] <= 8'h10 ;
			data[10463] <= 8'h10 ;
			data[10464] <= 8'h10 ;
			data[10465] <= 8'h10 ;
			data[10466] <= 8'h10 ;
			data[10467] <= 8'h10 ;
			data[10468] <= 8'h10 ;
			data[10469] <= 8'h10 ;
			data[10470] <= 8'h10 ;
			data[10471] <= 8'h10 ;
			data[10472] <= 8'h10 ;
			data[10473] <= 8'h10 ;
			data[10474] <= 8'h10 ;
			data[10475] <= 8'h10 ;
			data[10476] <= 8'h10 ;
			data[10477] <= 8'h10 ;
			data[10478] <= 8'h10 ;
			data[10479] <= 8'h10 ;
			data[10480] <= 8'h10 ;
			data[10481] <= 8'h10 ;
			data[10482] <= 8'h10 ;
			data[10483] <= 8'h10 ;
			data[10484] <= 8'h10 ;
			data[10485] <= 8'h10 ;
			data[10486] <= 8'h10 ;
			data[10487] <= 8'h10 ;
			data[10488] <= 8'h10 ;
			data[10489] <= 8'h10 ;
			data[10490] <= 8'h10 ;
			data[10491] <= 8'h10 ;
			data[10492] <= 8'h10 ;
			data[10493] <= 8'h10 ;
			data[10494] <= 8'h10 ;
			data[10495] <= 8'h10 ;
			data[10496] <= 8'h10 ;
			data[10497] <= 8'h10 ;
			data[10498] <= 8'h10 ;
			data[10499] <= 8'h10 ;
			data[10500] <= 8'h10 ;
			data[10501] <= 8'h10 ;
			data[10502] <= 8'h10 ;
			data[10503] <= 8'h10 ;
			data[10504] <= 8'h10 ;
			data[10505] <= 8'h10 ;
			data[10506] <= 8'h10 ;
			data[10507] <= 8'h10 ;
			data[10508] <= 8'h10 ;
			data[10509] <= 8'h10 ;
			data[10510] <= 8'h10 ;
			data[10511] <= 8'h10 ;
			data[10512] <= 8'h10 ;
			data[10513] <= 8'h10 ;
			data[10514] <= 8'h10 ;
			data[10515] <= 8'h10 ;
			data[10516] <= 8'h10 ;
			data[10517] <= 8'h10 ;
			data[10518] <= 8'h10 ;
			data[10519] <= 8'h10 ;
			data[10520] <= 8'h10 ;
			data[10521] <= 8'h10 ;
			data[10522] <= 8'h10 ;
			data[10523] <= 8'h10 ;
			data[10524] <= 8'h10 ;
			data[10525] <= 8'h10 ;
			data[10526] <= 8'h10 ;
			data[10527] <= 8'h10 ;
			data[10528] <= 8'h10 ;
			data[10529] <= 8'h10 ;
			data[10530] <= 8'h10 ;
			data[10531] <= 8'h10 ;
			data[10532] <= 8'h10 ;
			data[10533] <= 8'h10 ;
			data[10534] <= 8'h10 ;
			data[10535] <= 8'h10 ;
			data[10536] <= 8'h10 ;
			data[10537] <= 8'h10 ;
			data[10538] <= 8'h10 ;
			data[10539] <= 8'h10 ;
			data[10540] <= 8'h10 ;
			data[10541] <= 8'h10 ;
			data[10542] <= 8'h10 ;
			data[10543] <= 8'h10 ;
			data[10544] <= 8'h10 ;
			data[10545] <= 8'h10 ;
			data[10546] <= 8'h10 ;
			data[10547] <= 8'h10 ;
			data[10548] <= 8'h10 ;
			data[10549] <= 8'h10 ;
			data[10550] <= 8'h10 ;
			data[10551] <= 8'h10 ;
			data[10552] <= 8'h10 ;
			data[10553] <= 8'h10 ;
			data[10554] <= 8'h10 ;
			data[10555] <= 8'h10 ;
			data[10556] <= 8'h10 ;
			data[10557] <= 8'h10 ;
			data[10558] <= 8'h10 ;
			data[10559] <= 8'h10 ;
			data[10560] <= 8'h10 ;
			data[10561] <= 8'h10 ;
			data[10562] <= 8'h10 ;
			data[10563] <= 8'h10 ;
			data[10564] <= 8'h10 ;
			data[10565] <= 8'h10 ;
			data[10566] <= 8'h10 ;
			data[10567] <= 8'h10 ;
			data[10568] <= 8'h10 ;
			data[10569] <= 8'h10 ;
			data[10570] <= 8'h10 ;
			data[10571] <= 8'h10 ;
			data[10572] <= 8'h10 ;
			data[10573] <= 8'h10 ;
			data[10574] <= 8'h10 ;
			data[10575] <= 8'h10 ;
			data[10576] <= 8'h10 ;
			data[10577] <= 8'h10 ;
			data[10578] <= 8'h10 ;
			data[10579] <= 8'h10 ;
			data[10580] <= 8'h10 ;
			data[10581] <= 8'h10 ;
			data[10582] <= 8'h10 ;
			data[10583] <= 8'h10 ;
			data[10584] <= 8'h10 ;
			data[10585] <= 8'h10 ;
			data[10586] <= 8'h10 ;
			data[10587] <= 8'h10 ;
			data[10588] <= 8'h10 ;
			data[10589] <= 8'h10 ;
			data[10590] <= 8'h10 ;
			data[10591] <= 8'h10 ;
			data[10592] <= 8'h10 ;
			data[10593] <= 8'h10 ;
			data[10594] <= 8'h10 ;
			data[10595] <= 8'h10 ;
			data[10596] <= 8'h10 ;
			data[10597] <= 8'h10 ;
			data[10598] <= 8'h10 ;
			data[10599] <= 8'h10 ;
			data[10600] <= 8'h10 ;
			data[10601] <= 8'h10 ;
			data[10602] <= 8'h10 ;
			data[10603] <= 8'h10 ;
			data[10604] <= 8'h10 ;
			data[10605] <= 8'h10 ;
			data[10606] <= 8'h10 ;
			data[10607] <= 8'h10 ;
			data[10608] <= 8'h10 ;
			data[10609] <= 8'h10 ;
			data[10610] <= 8'h10 ;
			data[10611] <= 8'h10 ;
			data[10612] <= 8'h10 ;
			data[10613] <= 8'h10 ;
			data[10614] <= 8'h10 ;
			data[10615] <= 8'h10 ;
			data[10616] <= 8'h10 ;
			data[10617] <= 8'h10 ;
			data[10618] <= 8'h10 ;
			data[10619] <= 8'h10 ;
			data[10620] <= 8'h10 ;
			data[10621] <= 8'h10 ;
			data[10622] <= 8'h10 ;
			data[10623] <= 8'h10 ;
			data[10624] <= 8'h10 ;
			data[10625] <= 8'h10 ;
			data[10626] <= 8'h10 ;
			data[10627] <= 8'h10 ;
			data[10628] <= 8'h10 ;
			data[10629] <= 8'h10 ;
			data[10630] <= 8'h10 ;
			data[10631] <= 8'h10 ;
			data[10632] <= 8'h10 ;
			data[10633] <= 8'h10 ;
			data[10634] <= 8'h10 ;
			data[10635] <= 8'h10 ;
			data[10636] <= 8'h10 ;
			data[10637] <= 8'h10 ;
			data[10638] <= 8'h10 ;
			data[10639] <= 8'h10 ;
			data[10640] <= 8'h10 ;
			data[10641] <= 8'h10 ;
			data[10642] <= 8'h10 ;
			data[10643] <= 8'h10 ;
			data[10644] <= 8'h10 ;
			data[10645] <= 8'h10 ;
			data[10646] <= 8'h10 ;
			data[10647] <= 8'h10 ;
			data[10648] <= 8'h10 ;
			data[10649] <= 8'h10 ;
			data[10650] <= 8'h10 ;
			data[10651] <= 8'h10 ;
			data[10652] <= 8'h10 ;
			data[10653] <= 8'h10 ;
			data[10654] <= 8'h10 ;
			data[10655] <= 8'h10 ;
			data[10656] <= 8'h10 ;
			data[10657] <= 8'h10 ;
			data[10658] <= 8'h10 ;
			data[10659] <= 8'h10 ;
			data[10660] <= 8'h10 ;
			data[10661] <= 8'h10 ;
			data[10662] <= 8'h10 ;
			data[10663] <= 8'h10 ;
			data[10664] <= 8'h10 ;
			data[10665] <= 8'h10 ;
			data[10666] <= 8'h10 ;
			data[10667] <= 8'h10 ;
			data[10668] <= 8'h10 ;
			data[10669] <= 8'h10 ;
			data[10670] <= 8'h10 ;
			data[10671] <= 8'h10 ;
			data[10672] <= 8'h10 ;
			data[10673] <= 8'h10 ;
			data[10674] <= 8'h10 ;
			data[10675] <= 8'h10 ;
			data[10676] <= 8'h10 ;
			data[10677] <= 8'h10 ;
			data[10678] <= 8'h10 ;
			data[10679] <= 8'h10 ;
			data[10680] <= 8'h10 ;
			data[10681] <= 8'h10 ;
			data[10682] <= 8'h10 ;
			data[10683] <= 8'h10 ;
			data[10684] <= 8'h10 ;
			data[10685] <= 8'h10 ;
			data[10686] <= 8'h10 ;
			data[10687] <= 8'h10 ;
			data[10688] <= 8'h10 ;
			data[10689] <= 8'h10 ;
			data[10690] <= 8'h10 ;
			data[10691] <= 8'h10 ;
			data[10692] <= 8'h10 ;
			data[10693] <= 8'h10 ;
			data[10694] <= 8'h10 ;
			data[10695] <= 8'h10 ;
			data[10696] <= 8'h10 ;
			data[10697] <= 8'h10 ;
			data[10698] <= 8'h10 ;
			data[10699] <= 8'h10 ;
			data[10700] <= 8'h10 ;
			data[10701] <= 8'h10 ;
			data[10702] <= 8'h10 ;
			data[10703] <= 8'h10 ;
			data[10704] <= 8'h10 ;
			data[10705] <= 8'h10 ;
			data[10706] <= 8'h10 ;
			data[10707] <= 8'h10 ;
			data[10708] <= 8'h10 ;
			data[10709] <= 8'h10 ;
			data[10710] <= 8'h10 ;
			data[10711] <= 8'h10 ;
			data[10712] <= 8'h10 ;
			data[10713] <= 8'h10 ;
			data[10714] <= 8'h10 ;
			data[10715] <= 8'h10 ;
			data[10716] <= 8'h10 ;
			data[10717] <= 8'h10 ;
			data[10718] <= 8'h10 ;
			data[10719] <= 8'h10 ;
			data[10720] <= 8'h10 ;
			data[10721] <= 8'h10 ;
			data[10722] <= 8'h10 ;
			data[10723] <= 8'h10 ;
			data[10724] <= 8'h10 ;
			data[10725] <= 8'h10 ;
			data[10726] <= 8'h10 ;
			data[10727] <= 8'h10 ;
			data[10728] <= 8'h10 ;
			data[10729] <= 8'h10 ;
			data[10730] <= 8'h10 ;
			data[10731] <= 8'h10 ;
			data[10732] <= 8'h10 ;
			data[10733] <= 8'h10 ;
			data[10734] <= 8'h10 ;
			data[10735] <= 8'h10 ;
			data[10736] <= 8'h10 ;
			data[10737] <= 8'h10 ;
			data[10738] <= 8'h10 ;
			data[10739] <= 8'h10 ;
			data[10740] <= 8'h10 ;
			data[10741] <= 8'h10 ;
			data[10742] <= 8'h10 ;
			data[10743] <= 8'h10 ;
			data[10744] <= 8'h10 ;
			data[10745] <= 8'h10 ;
			data[10746] <= 8'h10 ;
			data[10747] <= 8'h10 ;
			data[10748] <= 8'h10 ;
			data[10749] <= 8'h10 ;
			data[10750] <= 8'h10 ;
			data[10751] <= 8'h10 ;
			data[10752] <= 8'h10 ;
			data[10753] <= 8'h10 ;
			data[10754] <= 8'h10 ;
			data[10755] <= 8'h10 ;
			data[10756] <= 8'h10 ;
			data[10757] <= 8'h10 ;
			data[10758] <= 8'h10 ;
			data[10759] <= 8'h10 ;
			data[10760] <= 8'h10 ;
			data[10761] <= 8'h10 ;
			data[10762] <= 8'h10 ;
			data[10763] <= 8'h10 ;
			data[10764] <= 8'h10 ;
			data[10765] <= 8'h10 ;
			data[10766] <= 8'h10 ;
			data[10767] <= 8'h10 ;
			data[10768] <= 8'h10 ;
			data[10769] <= 8'h10 ;
			data[10770] <= 8'h10 ;
			data[10771] <= 8'h10 ;
			data[10772] <= 8'h10 ;
			data[10773] <= 8'h10 ;
			data[10774] <= 8'h10 ;
			data[10775] <= 8'h10 ;
			data[10776] <= 8'h10 ;
			data[10777] <= 8'h10 ;
			data[10778] <= 8'h10 ;
			data[10779] <= 8'h10 ;
			data[10780] <= 8'h10 ;
			data[10781] <= 8'h10 ;
			data[10782] <= 8'h10 ;
			data[10783] <= 8'h10 ;
			data[10784] <= 8'h10 ;
			data[10785] <= 8'h10 ;
			data[10786] <= 8'h10 ;
			data[10787] <= 8'h10 ;
			data[10788] <= 8'h10 ;
			data[10789] <= 8'h10 ;
			data[10790] <= 8'h10 ;
			data[10791] <= 8'h10 ;
			data[10792] <= 8'h10 ;
			data[10793] <= 8'h10 ;
			data[10794] <= 8'h10 ;
			data[10795] <= 8'h10 ;
			data[10796] <= 8'h10 ;
			data[10797] <= 8'h10 ;
			data[10798] <= 8'h10 ;
			data[10799] <= 8'h10 ;
			data[10800] <= 8'h10 ;
			data[10801] <= 8'h10 ;
			data[10802] <= 8'h10 ;
			data[10803] <= 8'h10 ;
			data[10804] <= 8'h10 ;
			data[10805] <= 8'h10 ;
			data[10806] <= 8'h10 ;
			data[10807] <= 8'h10 ;
			data[10808] <= 8'h10 ;
			data[10809] <= 8'h10 ;
			data[10810] <= 8'h10 ;
			data[10811] <= 8'h10 ;
			data[10812] <= 8'h10 ;
			data[10813] <= 8'h10 ;
			data[10814] <= 8'h10 ;
			data[10815] <= 8'h10 ;
			data[10816] <= 8'h10 ;
			data[10817] <= 8'h10 ;
			data[10818] <= 8'h10 ;
			data[10819] <= 8'h10 ;
			data[10820] <= 8'h10 ;
			data[10821] <= 8'h10 ;
			data[10822] <= 8'h10 ;
			data[10823] <= 8'h10 ;
			data[10824] <= 8'h10 ;
			data[10825] <= 8'h10 ;
			data[10826] <= 8'h10 ;
			data[10827] <= 8'h10 ;
			data[10828] <= 8'h10 ;
			data[10829] <= 8'h10 ;
			data[10830] <= 8'h10 ;
			data[10831] <= 8'h10 ;
			data[10832] <= 8'h10 ;
			data[10833] <= 8'h10 ;
			data[10834] <= 8'h10 ;
			data[10835] <= 8'h10 ;
			data[10836] <= 8'h10 ;
			data[10837] <= 8'h10 ;
			data[10838] <= 8'h10 ;
			data[10839] <= 8'h10 ;
			data[10840] <= 8'h10 ;
			data[10841] <= 8'h10 ;
			data[10842] <= 8'h10 ;
			data[10843] <= 8'h10 ;
			data[10844] <= 8'h10 ;
			data[10845] <= 8'h10 ;
			data[10846] <= 8'h10 ;
			data[10847] <= 8'h10 ;
			data[10848] <= 8'h10 ;
			data[10849] <= 8'h10 ;
			data[10850] <= 8'h10 ;
			data[10851] <= 8'h10 ;
			data[10852] <= 8'h10 ;
			data[10853] <= 8'h10 ;
			data[10854] <= 8'h10 ;
			data[10855] <= 8'h10 ;
			data[10856] <= 8'h10 ;
			data[10857] <= 8'h10 ;
			data[10858] <= 8'h10 ;
			data[10859] <= 8'h10 ;
			data[10860] <= 8'h10 ;
			data[10861] <= 8'h10 ;
			data[10862] <= 8'h10 ;
			data[10863] <= 8'h10 ;
			data[10864] <= 8'h10 ;
			data[10865] <= 8'h10 ;
			data[10866] <= 8'h10 ;
			data[10867] <= 8'h10 ;
			data[10868] <= 8'h10 ;
			data[10869] <= 8'h10 ;
			data[10870] <= 8'h10 ;
			data[10871] <= 8'h10 ;
			data[10872] <= 8'h10 ;
			data[10873] <= 8'h10 ;
			data[10874] <= 8'h10 ;
			data[10875] <= 8'h10 ;
			data[10876] <= 8'h10 ;
			data[10877] <= 8'h10 ;
			data[10878] <= 8'h10 ;
			data[10879] <= 8'h10 ;
			data[10880] <= 8'h10 ;
			data[10881] <= 8'h10 ;
			data[10882] <= 8'h10 ;
			data[10883] <= 8'h10 ;
			data[10884] <= 8'h10 ;
			data[10885] <= 8'h10 ;
			data[10886] <= 8'h10 ;
			data[10887] <= 8'h10 ;
			data[10888] <= 8'h10 ;
			data[10889] <= 8'h10 ;
			data[10890] <= 8'h10 ;
			data[10891] <= 8'h10 ;
			data[10892] <= 8'h10 ;
			data[10893] <= 8'h10 ;
			data[10894] <= 8'h10 ;
			data[10895] <= 8'h10 ;
			data[10896] <= 8'h10 ;
			data[10897] <= 8'h10 ;
			data[10898] <= 8'h10 ;
			data[10899] <= 8'h10 ;
			data[10900] <= 8'h10 ;
			data[10901] <= 8'h10 ;
			data[10902] <= 8'h10 ;
			data[10903] <= 8'h10 ;
			data[10904] <= 8'h10 ;
			data[10905] <= 8'h10 ;
			data[10906] <= 8'h10 ;
			data[10907] <= 8'h10 ;
			data[10908] <= 8'h10 ;
			data[10909] <= 8'h10 ;
			data[10910] <= 8'h10 ;
			data[10911] <= 8'h10 ;
			data[10912] <= 8'h10 ;
			data[10913] <= 8'h10 ;
			data[10914] <= 8'h10 ;
			data[10915] <= 8'h10 ;
			data[10916] <= 8'h10 ;
			data[10917] <= 8'h10 ;
			data[10918] <= 8'h10 ;
			data[10919] <= 8'h10 ;
			data[10920] <= 8'h10 ;
			data[10921] <= 8'h10 ;
			data[10922] <= 8'h10 ;
			data[10923] <= 8'h10 ;
			data[10924] <= 8'h10 ;
			data[10925] <= 8'h10 ;
			data[10926] <= 8'h10 ;
			data[10927] <= 8'h10 ;
			data[10928] <= 8'h10 ;
			data[10929] <= 8'h10 ;
			data[10930] <= 8'h10 ;
			data[10931] <= 8'h10 ;
			data[10932] <= 8'h10 ;
			data[10933] <= 8'h10 ;
			data[10934] <= 8'h10 ;
			data[10935] <= 8'h10 ;
			data[10936] <= 8'h10 ;
			data[10937] <= 8'h10 ;
			data[10938] <= 8'h10 ;
			data[10939] <= 8'h10 ;
			data[10940] <= 8'h10 ;
			data[10941] <= 8'h10 ;
			data[10942] <= 8'h10 ;
			data[10943] <= 8'h10 ;
			data[10944] <= 8'h10 ;
			data[10945] <= 8'h10 ;
			data[10946] <= 8'h10 ;
			data[10947] <= 8'h10 ;
			data[10948] <= 8'h10 ;
			data[10949] <= 8'h10 ;
			data[10950] <= 8'h10 ;
			data[10951] <= 8'h10 ;
			data[10952] <= 8'h10 ;
			data[10953] <= 8'h10 ;
			data[10954] <= 8'h10 ;
			data[10955] <= 8'h10 ;
			data[10956] <= 8'h10 ;
			data[10957] <= 8'h10 ;
			data[10958] <= 8'h10 ;
			data[10959] <= 8'h10 ;
			data[10960] <= 8'h10 ;
			data[10961] <= 8'h10 ;
			data[10962] <= 8'h10 ;
			data[10963] <= 8'h10 ;
			data[10964] <= 8'h10 ;
			data[10965] <= 8'h10 ;
			data[10966] <= 8'h10 ;
			data[10967] <= 8'h10 ;
			data[10968] <= 8'h10 ;
			data[10969] <= 8'h10 ;
			data[10970] <= 8'h10 ;
			data[10971] <= 8'h10 ;
			data[10972] <= 8'h10 ;
			data[10973] <= 8'h10 ;
			data[10974] <= 8'h10 ;
			data[10975] <= 8'h10 ;
			data[10976] <= 8'h10 ;
			data[10977] <= 8'h10 ;
			data[10978] <= 8'h10 ;
			data[10979] <= 8'h10 ;
			data[10980] <= 8'h10 ;
			data[10981] <= 8'h10 ;
			data[10982] <= 8'h10 ;
			data[10983] <= 8'h10 ;
			data[10984] <= 8'h10 ;
			data[10985] <= 8'h10 ;
			data[10986] <= 8'h10 ;
			data[10987] <= 8'h10 ;
			data[10988] <= 8'h10 ;
			data[10989] <= 8'h10 ;
			data[10990] <= 8'h10 ;
			data[10991] <= 8'h10 ;
			data[10992] <= 8'h10 ;
			data[10993] <= 8'h10 ;
			data[10994] <= 8'h10 ;
			data[10995] <= 8'h10 ;
			data[10996] <= 8'h10 ;
			data[10997] <= 8'h10 ;
			data[10998] <= 8'h10 ;
			data[10999] <= 8'h10 ;
			data[11000] <= 8'h10 ;
			data[11001] <= 8'h10 ;
			data[11002] <= 8'h10 ;
			data[11003] <= 8'h10 ;
			data[11004] <= 8'h10 ;
			data[11005] <= 8'h10 ;
			data[11006] <= 8'h10 ;
			data[11007] <= 8'h10 ;
			data[11008] <= 8'h10 ;
			data[11009] <= 8'h10 ;
			data[11010] <= 8'h10 ;
			data[11011] <= 8'h10 ;
			data[11012] <= 8'h10 ;
			data[11013] <= 8'h10 ;
			data[11014] <= 8'h10 ;
			data[11015] <= 8'h10 ;
			data[11016] <= 8'h10 ;
			data[11017] <= 8'h10 ;
			data[11018] <= 8'h10 ;
			data[11019] <= 8'h10 ;
			data[11020] <= 8'h10 ;
			data[11021] <= 8'h10 ;
			data[11022] <= 8'h10 ;
			data[11023] <= 8'h10 ;
			data[11024] <= 8'h10 ;
			data[11025] <= 8'h10 ;
			data[11026] <= 8'h10 ;
			data[11027] <= 8'h10 ;
			data[11028] <= 8'h10 ;
			data[11029] <= 8'h10 ;
			data[11030] <= 8'h10 ;
			data[11031] <= 8'h10 ;
			data[11032] <= 8'h10 ;
			data[11033] <= 8'h10 ;
			data[11034] <= 8'h10 ;
			data[11035] <= 8'h10 ;
			data[11036] <= 8'h10 ;
			data[11037] <= 8'h10 ;
			data[11038] <= 8'h10 ;
			data[11039] <= 8'h10 ;
			data[11040] <= 8'h10 ;
			data[11041] <= 8'h10 ;
			data[11042] <= 8'h10 ;
			data[11043] <= 8'h10 ;
			data[11044] <= 8'h10 ;
			data[11045] <= 8'h10 ;
			data[11046] <= 8'h10 ;
			data[11047] <= 8'h10 ;
			data[11048] <= 8'h10 ;
			data[11049] <= 8'h10 ;
			data[11050] <= 8'h10 ;
			data[11051] <= 8'h10 ;
			data[11052] <= 8'h10 ;
			data[11053] <= 8'h10 ;
			data[11054] <= 8'h10 ;
			data[11055] <= 8'h10 ;
			data[11056] <= 8'h10 ;
			data[11057] <= 8'h10 ;
			data[11058] <= 8'h10 ;
			data[11059] <= 8'h10 ;
			data[11060] <= 8'h10 ;
			data[11061] <= 8'h10 ;
			data[11062] <= 8'h10 ;
			data[11063] <= 8'h10 ;
			data[11064] <= 8'h10 ;
			data[11065] <= 8'h10 ;
			data[11066] <= 8'h10 ;
			data[11067] <= 8'h10 ;
			data[11068] <= 8'h10 ;
			data[11069] <= 8'h10 ;
			data[11070] <= 8'h10 ;
			data[11071] <= 8'h10 ;
			data[11072] <= 8'h10 ;
			data[11073] <= 8'h10 ;
			data[11074] <= 8'h10 ;
			data[11075] <= 8'h10 ;
			data[11076] <= 8'h10 ;
			data[11077] <= 8'h10 ;
			data[11078] <= 8'h10 ;
			data[11079] <= 8'h10 ;
			data[11080] <= 8'h10 ;
			data[11081] <= 8'h10 ;
			data[11082] <= 8'h10 ;
			data[11083] <= 8'h10 ;
			data[11084] <= 8'h10 ;
			data[11085] <= 8'h10 ;
			data[11086] <= 8'h10 ;
			data[11087] <= 8'h10 ;
			data[11088] <= 8'h10 ;
			data[11089] <= 8'h10 ;
			data[11090] <= 8'h10 ;
			data[11091] <= 8'h10 ;
			data[11092] <= 8'h10 ;
			data[11093] <= 8'h10 ;
			data[11094] <= 8'h10 ;
			data[11095] <= 8'h10 ;
			data[11096] <= 8'h10 ;
			data[11097] <= 8'h10 ;
			data[11098] <= 8'h10 ;
			data[11099] <= 8'h10 ;
			data[11100] <= 8'h10 ;
			data[11101] <= 8'h10 ;
			data[11102] <= 8'h10 ;
			data[11103] <= 8'h10 ;
			data[11104] <= 8'h10 ;
			data[11105] <= 8'h10 ;
			data[11106] <= 8'h10 ;
			data[11107] <= 8'h10 ;
			data[11108] <= 8'h10 ;
			data[11109] <= 8'h10 ;
			data[11110] <= 8'h10 ;
			data[11111] <= 8'h10 ;
			data[11112] <= 8'h10 ;
			data[11113] <= 8'h10 ;
			data[11114] <= 8'h10 ;
			data[11115] <= 8'h10 ;
			data[11116] <= 8'h10 ;
			data[11117] <= 8'h10 ;
			data[11118] <= 8'h10 ;
			data[11119] <= 8'h10 ;
			data[11120] <= 8'h10 ;
			data[11121] <= 8'h10 ;
			data[11122] <= 8'h10 ;
			data[11123] <= 8'h10 ;
			data[11124] <= 8'h10 ;
			data[11125] <= 8'h10 ;
			data[11126] <= 8'h10 ;
			data[11127] <= 8'h10 ;
			data[11128] <= 8'h10 ;
			data[11129] <= 8'h10 ;
			data[11130] <= 8'h10 ;
			data[11131] <= 8'h10 ;
			data[11132] <= 8'h10 ;
			data[11133] <= 8'h10 ;
			data[11134] <= 8'h10 ;
			data[11135] <= 8'h10 ;
			data[11136] <= 8'h10 ;
			data[11137] <= 8'h10 ;
			data[11138] <= 8'h10 ;
			data[11139] <= 8'h10 ;
			data[11140] <= 8'h10 ;
			data[11141] <= 8'h10 ;
			data[11142] <= 8'h10 ;
			data[11143] <= 8'h10 ;
			data[11144] <= 8'h10 ;
			data[11145] <= 8'h10 ;
			data[11146] <= 8'h10 ;
			data[11147] <= 8'h10 ;
			data[11148] <= 8'h10 ;
			data[11149] <= 8'h10 ;
			data[11150] <= 8'h10 ;
			data[11151] <= 8'h10 ;
			data[11152] <= 8'h10 ;
			data[11153] <= 8'h10 ;
			data[11154] <= 8'h10 ;
			data[11155] <= 8'h10 ;
			data[11156] <= 8'h10 ;
			data[11157] <= 8'h10 ;
			data[11158] <= 8'h10 ;
			data[11159] <= 8'h10 ;
			data[11160] <= 8'h10 ;
			data[11161] <= 8'h10 ;
			data[11162] <= 8'h10 ;
			data[11163] <= 8'h10 ;
			data[11164] <= 8'h10 ;
			data[11165] <= 8'h10 ;
			data[11166] <= 8'h10 ;
			data[11167] <= 8'h10 ;
			data[11168] <= 8'h10 ;
			data[11169] <= 8'h10 ;
			data[11170] <= 8'h10 ;
			data[11171] <= 8'h10 ;
			data[11172] <= 8'h10 ;
			data[11173] <= 8'h10 ;
			data[11174] <= 8'h10 ;
			data[11175] <= 8'h10 ;
			data[11176] <= 8'h10 ;
			data[11177] <= 8'h10 ;
			data[11178] <= 8'h10 ;
			data[11179] <= 8'h10 ;
			data[11180] <= 8'h10 ;
			data[11181] <= 8'h10 ;
			data[11182] <= 8'h10 ;
			data[11183] <= 8'h10 ;
			data[11184] <= 8'h10 ;
			data[11185] <= 8'h10 ;
			data[11186] <= 8'h10 ;
			data[11187] <= 8'h10 ;
			data[11188] <= 8'h10 ;
			data[11189] <= 8'h10 ;
			data[11190] <= 8'h10 ;
			data[11191] <= 8'h10 ;
			data[11192] <= 8'h10 ;
			data[11193] <= 8'h10 ;
			data[11194] <= 8'h10 ;
			data[11195] <= 8'h10 ;
			data[11196] <= 8'h10 ;
			data[11197] <= 8'h10 ;
			data[11198] <= 8'h10 ;
			data[11199] <= 8'h10 ;
			data[11200] <= 8'h10 ;
			data[11201] <= 8'h10 ;
			data[11202] <= 8'h10 ;
			data[11203] <= 8'h10 ;
			data[11204] <= 8'h10 ;
			data[11205] <= 8'h10 ;
			data[11206] <= 8'h10 ;
			data[11207] <= 8'h10 ;
			data[11208] <= 8'h10 ;
			data[11209] <= 8'h10 ;
			data[11210] <= 8'h10 ;
			data[11211] <= 8'h10 ;
			data[11212] <= 8'h10 ;
			data[11213] <= 8'h10 ;
			data[11214] <= 8'h10 ;
			data[11215] <= 8'h10 ;
			data[11216] <= 8'h10 ;
			data[11217] <= 8'h10 ;
			data[11218] <= 8'h10 ;
			data[11219] <= 8'h10 ;
			data[11220] <= 8'h10 ;
			data[11221] <= 8'h10 ;
			data[11222] <= 8'h10 ;
			data[11223] <= 8'h10 ;
			data[11224] <= 8'h10 ;
			data[11225] <= 8'h10 ;
			data[11226] <= 8'h10 ;
			data[11227] <= 8'h10 ;
			data[11228] <= 8'h10 ;
			data[11229] <= 8'h10 ;
			data[11230] <= 8'h10 ;
			data[11231] <= 8'h10 ;
			data[11232] <= 8'h10 ;
			data[11233] <= 8'h10 ;
			data[11234] <= 8'h10 ;
			data[11235] <= 8'h10 ;
			data[11236] <= 8'h10 ;
			data[11237] <= 8'h10 ;
			data[11238] <= 8'h10 ;
			data[11239] <= 8'h10 ;
			data[11240] <= 8'h10 ;
			data[11241] <= 8'h10 ;
			data[11242] <= 8'h10 ;
			data[11243] <= 8'h10 ;
			data[11244] <= 8'h10 ;
			data[11245] <= 8'h10 ;
			data[11246] <= 8'h10 ;
			data[11247] <= 8'h10 ;
			data[11248] <= 8'h10 ;
			data[11249] <= 8'h10 ;
			data[11250] <= 8'h10 ;
			data[11251] <= 8'h10 ;
			data[11252] <= 8'h10 ;
			data[11253] <= 8'h10 ;
			data[11254] <= 8'h10 ;
			data[11255] <= 8'h10 ;
			data[11256] <= 8'h10 ;
			data[11257] <= 8'h10 ;
			data[11258] <= 8'h10 ;
			data[11259] <= 8'h10 ;
			data[11260] <= 8'h10 ;
			data[11261] <= 8'h10 ;
			data[11262] <= 8'h10 ;
			data[11263] <= 8'h10 ;
			data[11264] <= 8'h10 ;
			data[11265] <= 8'h10 ;
			data[11266] <= 8'h10 ;
			data[11267] <= 8'h10 ;
			data[11268] <= 8'h10 ;
			data[11269] <= 8'h10 ;
			data[11270] <= 8'h10 ;
			data[11271] <= 8'h10 ;
			data[11272] <= 8'h10 ;
			data[11273] <= 8'h10 ;
			data[11274] <= 8'h10 ;
			data[11275] <= 8'h10 ;
			data[11276] <= 8'h10 ;
			data[11277] <= 8'h10 ;
			data[11278] <= 8'h10 ;
			data[11279] <= 8'h10 ;
			data[11280] <= 8'h10 ;
			data[11281] <= 8'h10 ;
			data[11282] <= 8'h10 ;
			data[11283] <= 8'h10 ;
			data[11284] <= 8'h10 ;
			data[11285] <= 8'h10 ;
			data[11286] <= 8'h10 ;
			data[11287] <= 8'h10 ;
			data[11288] <= 8'h10 ;
			data[11289] <= 8'h10 ;
			data[11290] <= 8'h10 ;
			data[11291] <= 8'h10 ;
			data[11292] <= 8'h10 ;
			data[11293] <= 8'h10 ;
			data[11294] <= 8'h10 ;
			data[11295] <= 8'h10 ;
			data[11296] <= 8'h10 ;
			data[11297] <= 8'h10 ;
			data[11298] <= 8'h10 ;
			data[11299] <= 8'h10 ;
			data[11300] <= 8'h10 ;
			data[11301] <= 8'h10 ;
			data[11302] <= 8'h10 ;
			data[11303] <= 8'h10 ;
			data[11304] <= 8'h10 ;
			data[11305] <= 8'h10 ;
			data[11306] <= 8'h10 ;
			data[11307] <= 8'h10 ;
			data[11308] <= 8'h10 ;
			data[11309] <= 8'h10 ;
			data[11310] <= 8'h10 ;
			data[11311] <= 8'h10 ;
			data[11312] <= 8'h10 ;
			data[11313] <= 8'h10 ;
			data[11314] <= 8'h10 ;
			data[11315] <= 8'h10 ;
			data[11316] <= 8'h10 ;
			data[11317] <= 8'h10 ;
			data[11318] <= 8'h10 ;
			data[11319] <= 8'h10 ;
			data[11320] <= 8'h10 ;
			data[11321] <= 8'h10 ;
			data[11322] <= 8'h10 ;
			data[11323] <= 8'h10 ;
			data[11324] <= 8'h10 ;
			data[11325] <= 8'h10 ;
			data[11326] <= 8'h10 ;
			data[11327] <= 8'h10 ;
			data[11328] <= 8'h10 ;
			data[11329] <= 8'h10 ;
			data[11330] <= 8'h10 ;
			data[11331] <= 8'h10 ;
			data[11332] <= 8'h10 ;
			data[11333] <= 8'h10 ;
			data[11334] <= 8'h10 ;
			data[11335] <= 8'h10 ;
			data[11336] <= 8'h10 ;
			data[11337] <= 8'h10 ;
			data[11338] <= 8'h10 ;
			data[11339] <= 8'h10 ;
			data[11340] <= 8'h10 ;
			data[11341] <= 8'h10 ;
			data[11342] <= 8'h10 ;
			data[11343] <= 8'h10 ;
			data[11344] <= 8'h10 ;
			data[11345] <= 8'h10 ;
			data[11346] <= 8'h10 ;
			data[11347] <= 8'h10 ;
			data[11348] <= 8'h10 ;
			data[11349] <= 8'h10 ;
			data[11350] <= 8'h10 ;
			data[11351] <= 8'h10 ;
			data[11352] <= 8'h10 ;
			data[11353] <= 8'h10 ;
			data[11354] <= 8'h10 ;
			data[11355] <= 8'h10 ;
			data[11356] <= 8'h10 ;
			data[11357] <= 8'h10 ;
			data[11358] <= 8'h10 ;
			data[11359] <= 8'h10 ;
			data[11360] <= 8'h10 ;
			data[11361] <= 8'h10 ;
			data[11362] <= 8'h10 ;
			data[11363] <= 8'h10 ;
			data[11364] <= 8'h10 ;
			data[11365] <= 8'h10 ;
			data[11366] <= 8'h10 ;
			data[11367] <= 8'h10 ;
			data[11368] <= 8'h10 ;
			data[11369] <= 8'h10 ;
			data[11370] <= 8'h10 ;
			data[11371] <= 8'h10 ;
			data[11372] <= 8'h10 ;
			data[11373] <= 8'h10 ;
			data[11374] <= 8'h10 ;
			data[11375] <= 8'h10 ;
			data[11376] <= 8'h10 ;
			data[11377] <= 8'h10 ;
			data[11378] <= 8'h10 ;
			data[11379] <= 8'h10 ;
			data[11380] <= 8'h10 ;
			data[11381] <= 8'h10 ;
			data[11382] <= 8'h10 ;
			data[11383] <= 8'h10 ;
			data[11384] <= 8'h10 ;
			data[11385] <= 8'h10 ;
			data[11386] <= 8'h10 ;
			data[11387] <= 8'h10 ;
			data[11388] <= 8'h10 ;
			data[11389] <= 8'h10 ;
			data[11390] <= 8'h10 ;
			data[11391] <= 8'h10 ;
			data[11392] <= 8'h10 ;
			data[11393] <= 8'h10 ;
			data[11394] <= 8'h10 ;
			data[11395] <= 8'h10 ;
			data[11396] <= 8'h10 ;
			data[11397] <= 8'h10 ;
			data[11398] <= 8'h10 ;
			data[11399] <= 8'h10 ;
			data[11400] <= 8'h10 ;
			data[11401] <= 8'h10 ;
			data[11402] <= 8'h10 ;
			data[11403] <= 8'h10 ;
			data[11404] <= 8'h10 ;
			data[11405] <= 8'h10 ;
			data[11406] <= 8'h10 ;
			data[11407] <= 8'h10 ;
			data[11408] <= 8'h10 ;
			data[11409] <= 8'h10 ;
			data[11410] <= 8'h10 ;
			data[11411] <= 8'h10 ;
			data[11412] <= 8'h10 ;
			data[11413] <= 8'h10 ;
			data[11414] <= 8'h10 ;
			data[11415] <= 8'h10 ;
			data[11416] <= 8'h10 ;
			data[11417] <= 8'h10 ;
			data[11418] <= 8'h10 ;
			data[11419] <= 8'h10 ;
			data[11420] <= 8'h10 ;
			data[11421] <= 8'h10 ;
			data[11422] <= 8'h10 ;
			data[11423] <= 8'h10 ;
			data[11424] <= 8'h10 ;
			data[11425] <= 8'h10 ;
			data[11426] <= 8'h10 ;
			data[11427] <= 8'h10 ;
			data[11428] <= 8'h10 ;
			data[11429] <= 8'h10 ;
			data[11430] <= 8'h10 ;
			data[11431] <= 8'h10 ;
			data[11432] <= 8'h10 ;
			data[11433] <= 8'h10 ;
			data[11434] <= 8'h10 ;
			data[11435] <= 8'h10 ;
			data[11436] <= 8'h10 ;
			data[11437] <= 8'h10 ;
			data[11438] <= 8'h10 ;
			data[11439] <= 8'h10 ;
			data[11440] <= 8'h10 ;
			data[11441] <= 8'h10 ;
			data[11442] <= 8'h10 ;
			data[11443] <= 8'h10 ;
			data[11444] <= 8'h10 ;
			data[11445] <= 8'h10 ;
			data[11446] <= 8'h10 ;
			data[11447] <= 8'h10 ;
			data[11448] <= 8'h10 ;
			data[11449] <= 8'h10 ;
			data[11450] <= 8'h10 ;
			data[11451] <= 8'h10 ;
			data[11452] <= 8'h10 ;
			data[11453] <= 8'h10 ;
			data[11454] <= 8'h10 ;
			data[11455] <= 8'h10 ;
			data[11456] <= 8'h10 ;
			data[11457] <= 8'h10 ;
			data[11458] <= 8'h10 ;
			data[11459] <= 8'h10 ;
			data[11460] <= 8'h10 ;
			data[11461] <= 8'h10 ;
			data[11462] <= 8'h10 ;
			data[11463] <= 8'h10 ;
			data[11464] <= 8'h10 ;
			data[11465] <= 8'h10 ;
			data[11466] <= 8'h10 ;
			data[11467] <= 8'h10 ;
			data[11468] <= 8'h10 ;
			data[11469] <= 8'h10 ;
			data[11470] <= 8'h10 ;
			data[11471] <= 8'h10 ;
			data[11472] <= 8'h10 ;
			data[11473] <= 8'h10 ;
			data[11474] <= 8'h10 ;
			data[11475] <= 8'h10 ;
			data[11476] <= 8'h10 ;
			data[11477] <= 8'h10 ;
			data[11478] <= 8'h10 ;
			data[11479] <= 8'h10 ;
			data[11480] <= 8'h10 ;
			data[11481] <= 8'h10 ;
			data[11482] <= 8'h10 ;
			data[11483] <= 8'h10 ;
			data[11484] <= 8'h10 ;
			data[11485] <= 8'h10 ;
			data[11486] <= 8'h10 ;
			data[11487] <= 8'h10 ;
			data[11488] <= 8'h10 ;
			data[11489] <= 8'h10 ;
			data[11490] <= 8'h10 ;
			data[11491] <= 8'h10 ;
			data[11492] <= 8'h10 ;
			data[11493] <= 8'h10 ;
			data[11494] <= 8'h10 ;
			data[11495] <= 8'h10 ;
			data[11496] <= 8'h10 ;
			data[11497] <= 8'h10 ;
			data[11498] <= 8'h10 ;
			data[11499] <= 8'h10 ;
			data[11500] <= 8'h10 ;
			data[11501] <= 8'h10 ;
			data[11502] <= 8'h10 ;
			data[11503] <= 8'h10 ;
			data[11504] <= 8'h10 ;
			data[11505] <= 8'h10 ;
			data[11506] <= 8'h10 ;
			data[11507] <= 8'h10 ;
			data[11508] <= 8'h10 ;
			data[11509] <= 8'h10 ;
			data[11510] <= 8'h10 ;
			data[11511] <= 8'h10 ;
			data[11512] <= 8'h10 ;
			data[11513] <= 8'h10 ;
			data[11514] <= 8'h10 ;
			data[11515] <= 8'h10 ;
			data[11516] <= 8'h10 ;
			data[11517] <= 8'h10 ;
			data[11518] <= 8'h10 ;
			data[11519] <= 8'h10 ;
			data[11520] <= 8'h10 ;
			data[11521] <= 8'h10 ;
			data[11522] <= 8'h10 ;
			data[11523] <= 8'h10 ;
			data[11524] <= 8'h10 ;
			data[11525] <= 8'h10 ;
			data[11526] <= 8'h10 ;
			data[11527] <= 8'h10 ;
			data[11528] <= 8'h10 ;
			data[11529] <= 8'h10 ;
			data[11530] <= 8'h10 ;
			data[11531] <= 8'h10 ;
			data[11532] <= 8'h10 ;
			data[11533] <= 8'h10 ;
			data[11534] <= 8'h10 ;
			data[11535] <= 8'h10 ;
			data[11536] <= 8'h10 ;
			data[11537] <= 8'h10 ;
			data[11538] <= 8'h10 ;
			data[11539] <= 8'h10 ;
			data[11540] <= 8'h10 ;
			data[11541] <= 8'h10 ;
			data[11542] <= 8'h10 ;
			data[11543] <= 8'h10 ;
			data[11544] <= 8'h10 ;
			data[11545] <= 8'h10 ;
			data[11546] <= 8'h10 ;
			data[11547] <= 8'h10 ;
			data[11548] <= 8'h10 ;
			data[11549] <= 8'h10 ;
			data[11550] <= 8'h10 ;
			data[11551] <= 8'h10 ;
			data[11552] <= 8'h10 ;
			data[11553] <= 8'h10 ;
			data[11554] <= 8'h10 ;
			data[11555] <= 8'h10 ;
			data[11556] <= 8'h10 ;
			data[11557] <= 8'h10 ;
			data[11558] <= 8'h10 ;
			data[11559] <= 8'h10 ;
			data[11560] <= 8'h10 ;
			data[11561] <= 8'h10 ;
			data[11562] <= 8'h10 ;
			data[11563] <= 8'h10 ;
			data[11564] <= 8'h10 ;
			data[11565] <= 8'h10 ;
			data[11566] <= 8'h10 ;
			data[11567] <= 8'h10 ;
			data[11568] <= 8'h10 ;
			data[11569] <= 8'h10 ;
			data[11570] <= 8'h10 ;
			data[11571] <= 8'h10 ;
			data[11572] <= 8'h10 ;
			data[11573] <= 8'h10 ;
			data[11574] <= 8'h10 ;
			data[11575] <= 8'h10 ;
			data[11576] <= 8'h10 ;
			data[11577] <= 8'h10 ;
			data[11578] <= 8'h10 ;
			data[11579] <= 8'h10 ;
			data[11580] <= 8'h10 ;
			data[11581] <= 8'h10 ;
			data[11582] <= 8'h10 ;
			data[11583] <= 8'h10 ;
			data[11584] <= 8'h10 ;
			data[11585] <= 8'h10 ;
			data[11586] <= 8'h10 ;
			data[11587] <= 8'h10 ;
			data[11588] <= 8'h10 ;
			data[11589] <= 8'h10 ;
			data[11590] <= 8'h10 ;
			data[11591] <= 8'h10 ;
			data[11592] <= 8'h10 ;
			data[11593] <= 8'h10 ;
			data[11594] <= 8'h10 ;
			data[11595] <= 8'h10 ;
			data[11596] <= 8'h10 ;
			data[11597] <= 8'h10 ;
			data[11598] <= 8'h10 ;
			data[11599] <= 8'h10 ;
			data[11600] <= 8'h10 ;
			data[11601] <= 8'h10 ;
			data[11602] <= 8'h10 ;
			data[11603] <= 8'h10 ;
			data[11604] <= 8'h10 ;
			data[11605] <= 8'h10 ;
			data[11606] <= 8'h10 ;
			data[11607] <= 8'h10 ;
			data[11608] <= 8'h10 ;
			data[11609] <= 8'h10 ;
			data[11610] <= 8'h10 ;
			data[11611] <= 8'h10 ;
			data[11612] <= 8'h10 ;
			data[11613] <= 8'h10 ;
			data[11614] <= 8'h10 ;
			data[11615] <= 8'h10 ;
			data[11616] <= 8'h10 ;
			data[11617] <= 8'h10 ;
			data[11618] <= 8'h10 ;
			data[11619] <= 8'h10 ;
			data[11620] <= 8'h10 ;
			data[11621] <= 8'h10 ;
			data[11622] <= 8'h10 ;
			data[11623] <= 8'h10 ;
			data[11624] <= 8'h10 ;
			data[11625] <= 8'h10 ;
			data[11626] <= 8'h10 ;
			data[11627] <= 8'h10 ;
			data[11628] <= 8'h10 ;
			data[11629] <= 8'h10 ;
			data[11630] <= 8'h10 ;
			data[11631] <= 8'h10 ;
			data[11632] <= 8'h10 ;
			data[11633] <= 8'h10 ;
			data[11634] <= 8'h10 ;
			data[11635] <= 8'h10 ;
			data[11636] <= 8'h10 ;
			data[11637] <= 8'h10 ;
			data[11638] <= 8'h10 ;
			data[11639] <= 8'h10 ;
			data[11640] <= 8'h10 ;
			data[11641] <= 8'h10 ;
			data[11642] <= 8'h10 ;
			data[11643] <= 8'h10 ;
			data[11644] <= 8'h10 ;
			data[11645] <= 8'h10 ;
			data[11646] <= 8'h10 ;
			data[11647] <= 8'h10 ;
			data[11648] <= 8'h10 ;
			data[11649] <= 8'h10 ;
			data[11650] <= 8'h10 ;
			data[11651] <= 8'h10 ;
			data[11652] <= 8'h10 ;
			data[11653] <= 8'h10 ;
			data[11654] <= 8'h10 ;
			data[11655] <= 8'h10 ;
			data[11656] <= 8'h10 ;
			data[11657] <= 8'h10 ;
			data[11658] <= 8'h10 ;
			data[11659] <= 8'h10 ;
			data[11660] <= 8'h10 ;
			data[11661] <= 8'h10 ;
			data[11662] <= 8'h10 ;
			data[11663] <= 8'h10 ;
			data[11664] <= 8'h10 ;
			data[11665] <= 8'h10 ;
			data[11666] <= 8'h10 ;
			data[11667] <= 8'h10 ;
			data[11668] <= 8'h10 ;
			data[11669] <= 8'h10 ;
			data[11670] <= 8'h10 ;
			data[11671] <= 8'h10 ;
			data[11672] <= 8'h10 ;
			data[11673] <= 8'h10 ;
			data[11674] <= 8'h10 ;
			data[11675] <= 8'h10 ;
			data[11676] <= 8'h10 ;
			data[11677] <= 8'h10 ;
			data[11678] <= 8'h10 ;
			data[11679] <= 8'h10 ;
			data[11680] <= 8'h10 ;
			data[11681] <= 8'h10 ;
			data[11682] <= 8'h10 ;
			data[11683] <= 8'h10 ;
			data[11684] <= 8'h10 ;
			data[11685] <= 8'h10 ;
			data[11686] <= 8'h10 ;
			data[11687] <= 8'h10 ;
			data[11688] <= 8'h10 ;
			data[11689] <= 8'h10 ;
			data[11690] <= 8'h10 ;
			data[11691] <= 8'h10 ;
			data[11692] <= 8'h10 ;
			data[11693] <= 8'h10 ;
			data[11694] <= 8'h10 ;
			data[11695] <= 8'h10 ;
			data[11696] <= 8'h10 ;
			data[11697] <= 8'h10 ;
			data[11698] <= 8'h10 ;
			data[11699] <= 8'h10 ;
			data[11700] <= 8'h10 ;
			data[11701] <= 8'h10 ;
			data[11702] <= 8'h10 ;
			data[11703] <= 8'h10 ;
			data[11704] <= 8'h10 ;
			data[11705] <= 8'h10 ;
			data[11706] <= 8'h10 ;
			data[11707] <= 8'h10 ;
			data[11708] <= 8'h10 ;
			data[11709] <= 8'h10 ;
			data[11710] <= 8'h10 ;
			data[11711] <= 8'h10 ;
			data[11712] <= 8'h10 ;
			data[11713] <= 8'h10 ;
			data[11714] <= 8'h10 ;
			data[11715] <= 8'h10 ;
			data[11716] <= 8'h10 ;
			data[11717] <= 8'h10 ;
			data[11718] <= 8'h10 ;
			data[11719] <= 8'h10 ;
			data[11720] <= 8'h10 ;
			data[11721] <= 8'h10 ;
			data[11722] <= 8'h10 ;
			data[11723] <= 8'h10 ;
			data[11724] <= 8'h10 ;
			data[11725] <= 8'h10 ;
			data[11726] <= 8'h10 ;
			data[11727] <= 8'h10 ;
			data[11728] <= 8'h10 ;
			data[11729] <= 8'h10 ;
			data[11730] <= 8'h10 ;
			data[11731] <= 8'h10 ;
			data[11732] <= 8'h10 ;
			data[11733] <= 8'h10 ;
			data[11734] <= 8'h10 ;
			data[11735] <= 8'h10 ;
			data[11736] <= 8'h10 ;
			data[11737] <= 8'h10 ;
			data[11738] <= 8'h10 ;
			data[11739] <= 8'h10 ;
			data[11740] <= 8'h10 ;
			data[11741] <= 8'h10 ;
			data[11742] <= 8'h10 ;
			data[11743] <= 8'h10 ;
			data[11744] <= 8'h10 ;
			data[11745] <= 8'h10 ;
			data[11746] <= 8'h10 ;
			data[11747] <= 8'h10 ;
			data[11748] <= 8'h10 ;
			data[11749] <= 8'h10 ;
			data[11750] <= 8'h10 ;
			data[11751] <= 8'h10 ;
			data[11752] <= 8'h10 ;
			data[11753] <= 8'h10 ;
			data[11754] <= 8'h10 ;
			data[11755] <= 8'h10 ;
			data[11756] <= 8'h10 ;
			data[11757] <= 8'h10 ;
			data[11758] <= 8'h10 ;
			data[11759] <= 8'h10 ;
			data[11760] <= 8'h10 ;
			data[11761] <= 8'h10 ;
			data[11762] <= 8'h10 ;
			data[11763] <= 8'h10 ;
			data[11764] <= 8'h10 ;
			data[11765] <= 8'h10 ;
			data[11766] <= 8'h10 ;
			data[11767] <= 8'h10 ;
			data[11768] <= 8'h10 ;
			data[11769] <= 8'h10 ;
			data[11770] <= 8'h10 ;
			data[11771] <= 8'h10 ;
			data[11772] <= 8'h10 ;
			data[11773] <= 8'h10 ;
			data[11774] <= 8'h10 ;
			data[11775] <= 8'h10 ;
			data[11776] <= 8'h10 ;
			data[11777] <= 8'h10 ;
			data[11778] <= 8'h10 ;
			data[11779] <= 8'h10 ;
			data[11780] <= 8'h10 ;
			data[11781] <= 8'h10 ;
			data[11782] <= 8'h10 ;
			data[11783] <= 8'h10 ;
			data[11784] <= 8'h10 ;
			data[11785] <= 8'h10 ;
			data[11786] <= 8'h10 ;
			data[11787] <= 8'h10 ;
			data[11788] <= 8'h10 ;
			data[11789] <= 8'h10 ;
			data[11790] <= 8'h10 ;
			data[11791] <= 8'h10 ;
			data[11792] <= 8'h10 ;
			data[11793] <= 8'h10 ;
			data[11794] <= 8'h10 ;
			data[11795] <= 8'h10 ;
			data[11796] <= 8'h10 ;
			data[11797] <= 8'h10 ;
			data[11798] <= 8'h10 ;
			data[11799] <= 8'h10 ;
			data[11800] <= 8'h10 ;
			data[11801] <= 8'h10 ;
			data[11802] <= 8'h10 ;
			data[11803] <= 8'h10 ;
			data[11804] <= 8'h10 ;
			data[11805] <= 8'h10 ;
			data[11806] <= 8'h10 ;
			data[11807] <= 8'h10 ;
			data[11808] <= 8'h10 ;
			data[11809] <= 8'h10 ;
			data[11810] <= 8'h10 ;
			data[11811] <= 8'h10 ;
			data[11812] <= 8'h10 ;
			data[11813] <= 8'h10 ;
			data[11814] <= 8'h10 ;
			data[11815] <= 8'h10 ;
			data[11816] <= 8'h10 ;
			data[11817] <= 8'h10 ;
			data[11818] <= 8'h10 ;
			data[11819] <= 8'h10 ;
			data[11820] <= 8'h10 ;
			data[11821] <= 8'h10 ;
			data[11822] <= 8'h10 ;
			data[11823] <= 8'h10 ;
			data[11824] <= 8'h10 ;
			data[11825] <= 8'h10 ;
			data[11826] <= 8'h10 ;
			data[11827] <= 8'h10 ;
			data[11828] <= 8'h10 ;
			data[11829] <= 8'h10 ;
			data[11830] <= 8'h10 ;
			data[11831] <= 8'h10 ;
			data[11832] <= 8'h10 ;
			data[11833] <= 8'h10 ;
			data[11834] <= 8'h10 ;
			data[11835] <= 8'h10 ;
			data[11836] <= 8'h10 ;
			data[11837] <= 8'h10 ;
			data[11838] <= 8'h10 ;
			data[11839] <= 8'h10 ;
			data[11840] <= 8'h10 ;
			data[11841] <= 8'h10 ;
			data[11842] <= 8'h10 ;
			data[11843] <= 8'h10 ;
			data[11844] <= 8'h10 ;
			data[11845] <= 8'h10 ;
			data[11846] <= 8'h10 ;
			data[11847] <= 8'h10 ;
			data[11848] <= 8'h10 ;
			data[11849] <= 8'h10 ;
			data[11850] <= 8'h10 ;
			data[11851] <= 8'h10 ;
			data[11852] <= 8'h10 ;
			data[11853] <= 8'h10 ;
			data[11854] <= 8'h10 ;
			data[11855] <= 8'h10 ;
			data[11856] <= 8'h10 ;
			data[11857] <= 8'h10 ;
			data[11858] <= 8'h10 ;
			data[11859] <= 8'h10 ;
			data[11860] <= 8'h10 ;
			data[11861] <= 8'h10 ;
			data[11862] <= 8'h10 ;
			data[11863] <= 8'h10 ;
			data[11864] <= 8'h10 ;
			data[11865] <= 8'h10 ;
			data[11866] <= 8'h10 ;
			data[11867] <= 8'h10 ;
			data[11868] <= 8'h10 ;
			data[11869] <= 8'h10 ;
			data[11870] <= 8'h10 ;
			data[11871] <= 8'h10 ;
			data[11872] <= 8'h10 ;
			data[11873] <= 8'h10 ;
			data[11874] <= 8'h10 ;
			data[11875] <= 8'h10 ;
			data[11876] <= 8'h10 ;
			data[11877] <= 8'h10 ;
			data[11878] <= 8'h10 ;
			data[11879] <= 8'h10 ;
			data[11880] <= 8'h10 ;
			data[11881] <= 8'h10 ;
			data[11882] <= 8'h10 ;
			data[11883] <= 8'h10 ;
			data[11884] <= 8'h10 ;
			data[11885] <= 8'h10 ;
			data[11886] <= 8'h10 ;
			data[11887] <= 8'h10 ;
			data[11888] <= 8'h10 ;
			data[11889] <= 8'h10 ;
			data[11890] <= 8'h10 ;
			data[11891] <= 8'h10 ;
			data[11892] <= 8'h10 ;
			data[11893] <= 8'h10 ;
			data[11894] <= 8'h10 ;
			data[11895] <= 8'h10 ;
			data[11896] <= 8'h10 ;
			data[11897] <= 8'h10 ;
			data[11898] <= 8'h10 ;
			data[11899] <= 8'h10 ;
			data[11900] <= 8'h10 ;
			data[11901] <= 8'h10 ;
			data[11902] <= 8'h10 ;
			data[11903] <= 8'h10 ;
			data[11904] <= 8'h10 ;
			data[11905] <= 8'h10 ;
			data[11906] <= 8'h10 ;
			data[11907] <= 8'h10 ;
			data[11908] <= 8'h10 ;
			data[11909] <= 8'h10 ;
			data[11910] <= 8'h10 ;
			data[11911] <= 8'h10 ;
			data[11912] <= 8'h10 ;
			data[11913] <= 8'h10 ;
			data[11914] <= 8'h10 ;
			data[11915] <= 8'h10 ;
			data[11916] <= 8'h10 ;
			data[11917] <= 8'h10 ;
			data[11918] <= 8'h10 ;
			data[11919] <= 8'h10 ;
			data[11920] <= 8'h10 ;
			data[11921] <= 8'h10 ;
			data[11922] <= 8'h10 ;
			data[11923] <= 8'h10 ;
			data[11924] <= 8'h10 ;
			data[11925] <= 8'h10 ;
			data[11926] <= 8'h10 ;
			data[11927] <= 8'h10 ;
			data[11928] <= 8'h10 ;
			data[11929] <= 8'h10 ;
			data[11930] <= 8'h10 ;
			data[11931] <= 8'h10 ;
			data[11932] <= 8'h10 ;
			data[11933] <= 8'h10 ;
			data[11934] <= 8'h10 ;
			data[11935] <= 8'h10 ;
			data[11936] <= 8'h10 ;
			data[11937] <= 8'h10 ;
			data[11938] <= 8'h10 ;
			data[11939] <= 8'h10 ;
			data[11940] <= 8'h10 ;
			data[11941] <= 8'h10 ;
			data[11942] <= 8'h10 ;
			data[11943] <= 8'h10 ;
			data[11944] <= 8'h10 ;
			data[11945] <= 8'h10 ;
			data[11946] <= 8'h10 ;
			data[11947] <= 8'h10 ;
			data[11948] <= 8'h10 ;
			data[11949] <= 8'h10 ;
			data[11950] <= 8'h10 ;
			data[11951] <= 8'h10 ;
			data[11952] <= 8'h10 ;
			data[11953] <= 8'h10 ;
			data[11954] <= 8'h10 ;
			data[11955] <= 8'h10 ;
			data[11956] <= 8'h10 ;
			data[11957] <= 8'h10 ;
			data[11958] <= 8'h10 ;
			data[11959] <= 8'h10 ;
			data[11960] <= 8'h10 ;
			data[11961] <= 8'h10 ;
			data[11962] <= 8'h10 ;
			data[11963] <= 8'h10 ;
			data[11964] <= 8'h10 ;
			data[11965] <= 8'h10 ;
			data[11966] <= 8'h10 ;
			data[11967] <= 8'h10 ;
			data[11968] <= 8'h10 ;
			data[11969] <= 8'h10 ;
			data[11970] <= 8'h10 ;
			data[11971] <= 8'h10 ;
			data[11972] <= 8'h10 ;
			data[11973] <= 8'h10 ;
			data[11974] <= 8'h10 ;
			data[11975] <= 8'h10 ;
			data[11976] <= 8'h10 ;
			data[11977] <= 8'h10 ;
			data[11978] <= 8'h10 ;
			data[11979] <= 8'h10 ;
			data[11980] <= 8'h10 ;
			data[11981] <= 8'h10 ;
			data[11982] <= 8'h10 ;
			data[11983] <= 8'h10 ;
			data[11984] <= 8'h10 ;
			data[11985] <= 8'h10 ;
			data[11986] <= 8'h10 ;
			data[11987] <= 8'h10 ;
			data[11988] <= 8'h10 ;
			data[11989] <= 8'h10 ;
			data[11990] <= 8'h10 ;
			data[11991] <= 8'h10 ;
			data[11992] <= 8'h10 ;
			data[11993] <= 8'h10 ;
			data[11994] <= 8'h10 ;
			data[11995] <= 8'h10 ;
			data[11996] <= 8'h10 ;
			data[11997] <= 8'h10 ;
			data[11998] <= 8'h10 ;
			data[11999] <= 8'h10 ;
			data[12000] <= 8'h10 ;
			data[12001] <= 8'h10 ;
			data[12002] <= 8'h10 ;
			data[12003] <= 8'h10 ;
			data[12004] <= 8'h10 ;
			data[12005] <= 8'h10 ;
			data[12006] <= 8'h10 ;
			data[12007] <= 8'h10 ;
			data[12008] <= 8'h10 ;
			data[12009] <= 8'h10 ;
			data[12010] <= 8'h10 ;
			data[12011] <= 8'h10 ;
			data[12012] <= 8'h10 ;
			data[12013] <= 8'h10 ;
			data[12014] <= 8'h10 ;
			data[12015] <= 8'h10 ;
			data[12016] <= 8'h10 ;
			data[12017] <= 8'h10 ;
			data[12018] <= 8'h10 ;
			data[12019] <= 8'h10 ;
			data[12020] <= 8'h10 ;
			data[12021] <= 8'h10 ;
			data[12022] <= 8'h10 ;
			data[12023] <= 8'h10 ;
			data[12024] <= 8'h10 ;
			data[12025] <= 8'h10 ;
			data[12026] <= 8'h10 ;
			data[12027] <= 8'h10 ;
			data[12028] <= 8'h10 ;
			data[12029] <= 8'h10 ;
			data[12030] <= 8'h10 ;
			data[12031] <= 8'h10 ;
			data[12032] <= 8'h10 ;
			data[12033] <= 8'h10 ;
			data[12034] <= 8'h10 ;
			data[12035] <= 8'h10 ;
			data[12036] <= 8'h10 ;
			data[12037] <= 8'h10 ;
			data[12038] <= 8'h10 ;
			data[12039] <= 8'h10 ;
			data[12040] <= 8'h10 ;
			data[12041] <= 8'h10 ;
			data[12042] <= 8'h10 ;
			data[12043] <= 8'h10 ;
			data[12044] <= 8'h10 ;
			data[12045] <= 8'h10 ;
			data[12046] <= 8'h10 ;
			data[12047] <= 8'h10 ;
			data[12048] <= 8'h10 ;
			data[12049] <= 8'h10 ;
			data[12050] <= 8'h10 ;
			data[12051] <= 8'h10 ;
			data[12052] <= 8'h10 ;
			data[12053] <= 8'h10 ;
			data[12054] <= 8'h10 ;
			data[12055] <= 8'h10 ;
			data[12056] <= 8'h10 ;
			data[12057] <= 8'h10 ;
			data[12058] <= 8'h10 ;
			data[12059] <= 8'h10 ;
			data[12060] <= 8'h10 ;
			data[12061] <= 8'h10 ;
			data[12062] <= 8'h10 ;
			data[12063] <= 8'h10 ;
			data[12064] <= 8'h10 ;
			data[12065] <= 8'h10 ;
			data[12066] <= 8'h10 ;
			data[12067] <= 8'h10 ;
			data[12068] <= 8'h10 ;
			data[12069] <= 8'h10 ;
			data[12070] <= 8'h10 ;
			data[12071] <= 8'h10 ;
			data[12072] <= 8'h10 ;
			data[12073] <= 8'h10 ;
			data[12074] <= 8'h10 ;
			data[12075] <= 8'h10 ;
			data[12076] <= 8'h10 ;
			data[12077] <= 8'h10 ;
			data[12078] <= 8'h10 ;
			data[12079] <= 8'h10 ;
			data[12080] <= 8'h10 ;
			data[12081] <= 8'h10 ;
			data[12082] <= 8'h10 ;
			data[12083] <= 8'h10 ;
			data[12084] <= 8'h10 ;
			data[12085] <= 8'h10 ;
			data[12086] <= 8'h10 ;
			data[12087] <= 8'h10 ;
			data[12088] <= 8'h10 ;
			data[12089] <= 8'h10 ;
			data[12090] <= 8'h10 ;
			data[12091] <= 8'h10 ;
			data[12092] <= 8'h10 ;
			data[12093] <= 8'h10 ;
			data[12094] <= 8'h10 ;
			data[12095] <= 8'h10 ;
			data[12096] <= 8'h10 ;
			data[12097] <= 8'h10 ;
			data[12098] <= 8'h10 ;
			data[12099] <= 8'h10 ;
			data[12100] <= 8'h10 ;
			data[12101] <= 8'h10 ;
			data[12102] <= 8'h10 ;
			data[12103] <= 8'h10 ;
			data[12104] <= 8'h10 ;
			data[12105] <= 8'h10 ;
			data[12106] <= 8'h10 ;
			data[12107] <= 8'h10 ;
			data[12108] <= 8'h10 ;
			data[12109] <= 8'h10 ;
			data[12110] <= 8'h10 ;
			data[12111] <= 8'h10 ;
			data[12112] <= 8'h10 ;
			data[12113] <= 8'h10 ;
			data[12114] <= 8'h10 ;
			data[12115] <= 8'h10 ;
			data[12116] <= 8'h10 ;
			data[12117] <= 8'h10 ;
			data[12118] <= 8'h10 ;
			data[12119] <= 8'h10 ;
			data[12120] <= 8'h10 ;
			data[12121] <= 8'h10 ;
			data[12122] <= 8'h10 ;
			data[12123] <= 8'h10 ;
			data[12124] <= 8'h10 ;
			data[12125] <= 8'h10 ;
			data[12126] <= 8'h10 ;
			data[12127] <= 8'h10 ;
			data[12128] <= 8'h10 ;
			data[12129] <= 8'h10 ;
			data[12130] <= 8'h10 ;
			data[12131] <= 8'h10 ;
			data[12132] <= 8'h10 ;
			data[12133] <= 8'h10 ;
			data[12134] <= 8'h10 ;
			data[12135] <= 8'h10 ;
			data[12136] <= 8'h10 ;
			data[12137] <= 8'h10 ;
			data[12138] <= 8'h10 ;
			data[12139] <= 8'h10 ;
			data[12140] <= 8'h10 ;
			data[12141] <= 8'h10 ;
			data[12142] <= 8'h10 ;
			data[12143] <= 8'h10 ;
			data[12144] <= 8'h10 ;
			data[12145] <= 8'h10 ;
			data[12146] <= 8'h10 ;
			data[12147] <= 8'h10 ;
			data[12148] <= 8'h10 ;
			data[12149] <= 8'h10 ;
			data[12150] <= 8'h10 ;
			data[12151] <= 8'h10 ;
			data[12152] <= 8'h10 ;
			data[12153] <= 8'h10 ;
			data[12154] <= 8'h10 ;
			data[12155] <= 8'h10 ;
			data[12156] <= 8'h10 ;
			data[12157] <= 8'h10 ;
			data[12158] <= 8'h10 ;
			data[12159] <= 8'h10 ;
			data[12160] <= 8'h10 ;
			data[12161] <= 8'h10 ;
			data[12162] <= 8'h10 ;
			data[12163] <= 8'h10 ;
			data[12164] <= 8'h10 ;
			data[12165] <= 8'h10 ;
			data[12166] <= 8'h10 ;
			data[12167] <= 8'h10 ;
			data[12168] <= 8'h10 ;
			data[12169] <= 8'h10 ;
			data[12170] <= 8'h10 ;
			data[12171] <= 8'h10 ;
			data[12172] <= 8'h10 ;
			data[12173] <= 8'h10 ;
			data[12174] <= 8'h10 ;
			data[12175] <= 8'h10 ;
			data[12176] <= 8'h10 ;
			data[12177] <= 8'h10 ;
			data[12178] <= 8'h10 ;
			data[12179] <= 8'h10 ;
			data[12180] <= 8'h10 ;
			data[12181] <= 8'h10 ;
			data[12182] <= 8'h10 ;
			data[12183] <= 8'h10 ;
			data[12184] <= 8'h10 ;
			data[12185] <= 8'h10 ;
			data[12186] <= 8'h10 ;
			data[12187] <= 8'h10 ;
			data[12188] <= 8'h10 ;
			data[12189] <= 8'h10 ;
			data[12190] <= 8'h10 ;
			data[12191] <= 8'h10 ;
			data[12192] <= 8'h10 ;
			data[12193] <= 8'h10 ;
			data[12194] <= 8'h10 ;
			data[12195] <= 8'h10 ;
			data[12196] <= 8'h10 ;
			data[12197] <= 8'h10 ;
			data[12198] <= 8'h10 ;
			data[12199] <= 8'h10 ;
			data[12200] <= 8'h10 ;
			data[12201] <= 8'h10 ;
			data[12202] <= 8'h10 ;
			data[12203] <= 8'h10 ;
			data[12204] <= 8'h10 ;
			data[12205] <= 8'h10 ;
			data[12206] <= 8'h10 ;
			data[12207] <= 8'h10 ;
			data[12208] <= 8'h10 ;
			data[12209] <= 8'h10 ;
			data[12210] <= 8'h10 ;
			data[12211] <= 8'h10 ;
			data[12212] <= 8'h10 ;
			data[12213] <= 8'h10 ;
			data[12214] <= 8'h10 ;
			data[12215] <= 8'h10 ;
			data[12216] <= 8'h10 ;
			data[12217] <= 8'h10 ;
			data[12218] <= 8'h10 ;
			data[12219] <= 8'h10 ;
			data[12220] <= 8'h10 ;
			data[12221] <= 8'h10 ;
			data[12222] <= 8'h10 ;
			data[12223] <= 8'h10 ;
			data[12224] <= 8'h10 ;
			data[12225] <= 8'h10 ;
			data[12226] <= 8'h10 ;
			data[12227] <= 8'h10 ;
			data[12228] <= 8'h10 ;
			data[12229] <= 8'h10 ;
			data[12230] <= 8'h10 ;
			data[12231] <= 8'h10 ;
			data[12232] <= 8'h10 ;
			data[12233] <= 8'h10 ;
			data[12234] <= 8'h10 ;
			data[12235] <= 8'h10 ;
			data[12236] <= 8'h10 ;
			data[12237] <= 8'h10 ;
			data[12238] <= 8'h10 ;
			data[12239] <= 8'h10 ;
			data[12240] <= 8'h10 ;
			data[12241] <= 8'h10 ;
			data[12242] <= 8'h10 ;
			data[12243] <= 8'h10 ;
			data[12244] <= 8'h10 ;
			data[12245] <= 8'h10 ;
			data[12246] <= 8'h10 ;
			data[12247] <= 8'h10 ;
			data[12248] <= 8'h10 ;
			data[12249] <= 8'h10 ;
			data[12250] <= 8'h10 ;
			data[12251] <= 8'h10 ;
			data[12252] <= 8'h10 ;
			data[12253] <= 8'h10 ;
			data[12254] <= 8'h10 ;
			data[12255] <= 8'h10 ;
			data[12256] <= 8'h10 ;
			data[12257] <= 8'h10 ;
			data[12258] <= 8'h10 ;
			data[12259] <= 8'h10 ;
			data[12260] <= 8'h10 ;
			data[12261] <= 8'h10 ;
			data[12262] <= 8'h10 ;
			data[12263] <= 8'h10 ;
			data[12264] <= 8'h10 ;
			data[12265] <= 8'h10 ;
			data[12266] <= 8'h10 ;
			data[12267] <= 8'h10 ;
			data[12268] <= 8'h10 ;
			data[12269] <= 8'h10 ;
			data[12270] <= 8'h10 ;
			data[12271] <= 8'h10 ;
			data[12272] <= 8'h10 ;
			data[12273] <= 8'h10 ;
			data[12274] <= 8'h10 ;
			data[12275] <= 8'h10 ;
			data[12276] <= 8'h10 ;
			data[12277] <= 8'h10 ;
			data[12278] <= 8'h10 ;
			data[12279] <= 8'h10 ;
			data[12280] <= 8'h10 ;
			data[12281] <= 8'h10 ;
			data[12282] <= 8'h10 ;
			data[12283] <= 8'h10 ;
			data[12284] <= 8'h10 ;
			data[12285] <= 8'h10 ;
			data[12286] <= 8'h10 ;
			data[12287] <= 8'h10 ;
			data[12288] <= 8'h10 ;
			data[12289] <= 8'h10 ;
			data[12290] <= 8'h10 ;
			data[12291] <= 8'h10 ;
			data[12292] <= 8'h10 ;
			data[12293] <= 8'h10 ;
			data[12294] <= 8'h10 ;
			data[12295] <= 8'h10 ;
			data[12296] <= 8'h10 ;
			data[12297] <= 8'h10 ;
			data[12298] <= 8'h10 ;
			data[12299] <= 8'h10 ;
			data[12300] <= 8'h10 ;
			data[12301] <= 8'h10 ;
			data[12302] <= 8'h10 ;
			data[12303] <= 8'h10 ;
			data[12304] <= 8'h10 ;
			data[12305] <= 8'h10 ;
			data[12306] <= 8'h10 ;
			data[12307] <= 8'h10 ;
			data[12308] <= 8'h10 ;
			data[12309] <= 8'h10 ;
			data[12310] <= 8'h10 ;
			data[12311] <= 8'h10 ;
			data[12312] <= 8'h10 ;
			data[12313] <= 8'h10 ;
			data[12314] <= 8'h10 ;
			data[12315] <= 8'h10 ;
			data[12316] <= 8'h10 ;
			data[12317] <= 8'h10 ;
			data[12318] <= 8'h10 ;
			data[12319] <= 8'h10 ;
			data[12320] <= 8'h10 ;
			data[12321] <= 8'h10 ;
			data[12322] <= 8'h10 ;
			data[12323] <= 8'h10 ;
			data[12324] <= 8'h10 ;
			data[12325] <= 8'h10 ;
			data[12326] <= 8'h10 ;
			data[12327] <= 8'h10 ;
			data[12328] <= 8'h10 ;
			data[12329] <= 8'h10 ;
			data[12330] <= 8'h10 ;
			data[12331] <= 8'h10 ;
			data[12332] <= 8'h10 ;
			data[12333] <= 8'h10 ;
			data[12334] <= 8'h10 ;
			data[12335] <= 8'h10 ;
			data[12336] <= 8'h10 ;
			data[12337] <= 8'h10 ;
			data[12338] <= 8'h10 ;
			data[12339] <= 8'h10 ;
			data[12340] <= 8'h10 ;
			data[12341] <= 8'h10 ;
			data[12342] <= 8'h10 ;
			data[12343] <= 8'h10 ;
			data[12344] <= 8'h10 ;
			data[12345] <= 8'h10 ;
			data[12346] <= 8'h10 ;
			data[12347] <= 8'h10 ;
			data[12348] <= 8'h10 ;
			data[12349] <= 8'h10 ;
			data[12350] <= 8'h10 ;
			data[12351] <= 8'h10 ;
			data[12352] <= 8'h10 ;
			data[12353] <= 8'h10 ;
			data[12354] <= 8'h10 ;
			data[12355] <= 8'h10 ;
			data[12356] <= 8'h10 ;
			data[12357] <= 8'h10 ;
			data[12358] <= 8'h10 ;
			data[12359] <= 8'h10 ;
			data[12360] <= 8'h10 ;
			data[12361] <= 8'h10 ;
			data[12362] <= 8'h10 ;
			data[12363] <= 8'h10 ;
			data[12364] <= 8'h10 ;
			data[12365] <= 8'h10 ;
			data[12366] <= 8'h10 ;
			data[12367] <= 8'h10 ;
			data[12368] <= 8'h10 ;
			data[12369] <= 8'h10 ;
			data[12370] <= 8'h10 ;
			data[12371] <= 8'h10 ;
			data[12372] <= 8'h10 ;
			data[12373] <= 8'h10 ;
			data[12374] <= 8'h10 ;
			data[12375] <= 8'h10 ;
			data[12376] <= 8'h10 ;
			data[12377] <= 8'h10 ;
			data[12378] <= 8'h10 ;
			data[12379] <= 8'h10 ;
			data[12380] <= 8'h10 ;
			data[12381] <= 8'h10 ;
			data[12382] <= 8'h10 ;
			data[12383] <= 8'h10 ;
			data[12384] <= 8'h10 ;
			data[12385] <= 8'h10 ;
			data[12386] <= 8'h10 ;
			data[12387] <= 8'h10 ;
			data[12388] <= 8'h10 ;
			data[12389] <= 8'h10 ;
			data[12390] <= 8'h10 ;
			data[12391] <= 8'h10 ;
			data[12392] <= 8'h10 ;
			data[12393] <= 8'h10 ;
			data[12394] <= 8'h10 ;
			data[12395] <= 8'h10 ;
			data[12396] <= 8'h10 ;
			data[12397] <= 8'h10 ;
			data[12398] <= 8'h10 ;
			data[12399] <= 8'h10 ;
			data[12400] <= 8'h10 ;
			data[12401] <= 8'h10 ;
			data[12402] <= 8'h10 ;
			data[12403] <= 8'h10 ;
			data[12404] <= 8'h10 ;
			data[12405] <= 8'h10 ;
			data[12406] <= 8'h10 ;
			data[12407] <= 8'h10 ;
			data[12408] <= 8'h10 ;
			data[12409] <= 8'h10 ;
			data[12410] <= 8'h10 ;
			data[12411] <= 8'h10 ;
			data[12412] <= 8'h10 ;
			data[12413] <= 8'h10 ;
			data[12414] <= 8'h10 ;
			data[12415] <= 8'h10 ;
			data[12416] <= 8'h10 ;
			data[12417] <= 8'h10 ;
			data[12418] <= 8'h10 ;
			data[12419] <= 8'h10 ;
			data[12420] <= 8'h10 ;
			data[12421] <= 8'h10 ;
			data[12422] <= 8'h10 ;
			data[12423] <= 8'h10 ;
			data[12424] <= 8'h10 ;
			data[12425] <= 8'h10 ;
			data[12426] <= 8'h10 ;
			data[12427] <= 8'h10 ;
			data[12428] <= 8'h10 ;
			data[12429] <= 8'h10 ;
			data[12430] <= 8'h10 ;
			data[12431] <= 8'h10 ;
			data[12432] <= 8'h10 ;
			data[12433] <= 8'h10 ;
			data[12434] <= 8'h10 ;
			data[12435] <= 8'h10 ;
			data[12436] <= 8'h10 ;
			data[12437] <= 8'h10 ;
			data[12438] <= 8'h10 ;
			data[12439] <= 8'h10 ;
			data[12440] <= 8'h10 ;
			data[12441] <= 8'h10 ;
			data[12442] <= 8'h10 ;
			data[12443] <= 8'h10 ;
			data[12444] <= 8'h10 ;
			data[12445] <= 8'h10 ;
			data[12446] <= 8'h10 ;
			data[12447] <= 8'h10 ;
			data[12448] <= 8'h10 ;
			data[12449] <= 8'h10 ;
			data[12450] <= 8'h10 ;
			data[12451] <= 8'h10 ;
			data[12452] <= 8'h10 ;
			data[12453] <= 8'h10 ;
			data[12454] <= 8'h10 ;
			data[12455] <= 8'h10 ;
			data[12456] <= 8'h10 ;
			data[12457] <= 8'h10 ;
			data[12458] <= 8'h10 ;
			data[12459] <= 8'h10 ;
			data[12460] <= 8'h10 ;
			data[12461] <= 8'h10 ;
			data[12462] <= 8'h10 ;
			data[12463] <= 8'h10 ;
			data[12464] <= 8'h10 ;
			data[12465] <= 8'h10 ;
			data[12466] <= 8'h10 ;
			data[12467] <= 8'h10 ;
			data[12468] <= 8'h10 ;
			data[12469] <= 8'h10 ;
			data[12470] <= 8'h10 ;
			data[12471] <= 8'h10 ;
			data[12472] <= 8'h10 ;
			data[12473] <= 8'h10 ;
			data[12474] <= 8'h10 ;
			data[12475] <= 8'h10 ;
			data[12476] <= 8'h10 ;
			data[12477] <= 8'h10 ;
			data[12478] <= 8'h10 ;
			data[12479] <= 8'h10 ;
			data[12480] <= 8'h10 ;
			data[12481] <= 8'h10 ;
			data[12482] <= 8'h10 ;
			data[12483] <= 8'h10 ;
			data[12484] <= 8'h10 ;
			data[12485] <= 8'h10 ;
			data[12486] <= 8'h10 ;
			data[12487] <= 8'h10 ;
			data[12488] <= 8'h10 ;
			data[12489] <= 8'h10 ;
			data[12490] <= 8'h10 ;
			data[12491] <= 8'h10 ;
			data[12492] <= 8'h10 ;
			data[12493] <= 8'h10 ;
			data[12494] <= 8'h10 ;
			data[12495] <= 8'h10 ;
			data[12496] <= 8'h10 ;
			data[12497] <= 8'h10 ;
			data[12498] <= 8'h10 ;
			data[12499] <= 8'h10 ;
			data[12500] <= 8'h10 ;
			data[12501] <= 8'h10 ;
			data[12502] <= 8'h10 ;
			data[12503] <= 8'h10 ;
			data[12504] <= 8'h10 ;
			data[12505] <= 8'h10 ;
			data[12506] <= 8'h10 ;
			data[12507] <= 8'h10 ;
			data[12508] <= 8'h10 ;
			data[12509] <= 8'h10 ;
			data[12510] <= 8'h10 ;
			data[12511] <= 8'h10 ;
			data[12512] <= 8'h10 ;
			data[12513] <= 8'h10 ;
			data[12514] <= 8'h10 ;
			data[12515] <= 8'h10 ;
			data[12516] <= 8'h10 ;
			data[12517] <= 8'h10 ;
			data[12518] <= 8'h10 ;
			data[12519] <= 8'h10 ;
			data[12520] <= 8'h10 ;
			data[12521] <= 8'h10 ;
			data[12522] <= 8'h10 ;
			data[12523] <= 8'h10 ;
			data[12524] <= 8'h10 ;
			data[12525] <= 8'h10 ;
			data[12526] <= 8'h10 ;
			data[12527] <= 8'h10 ;
			data[12528] <= 8'h10 ;
			data[12529] <= 8'h10 ;
			data[12530] <= 8'h10 ;
			data[12531] <= 8'h10 ;
			data[12532] <= 8'h10 ;
			data[12533] <= 8'h10 ;
			data[12534] <= 8'h10 ;
			data[12535] <= 8'h10 ;
			data[12536] <= 8'h10 ;
			data[12537] <= 8'h10 ;
			data[12538] <= 8'h10 ;
			data[12539] <= 8'h10 ;
			data[12540] <= 8'h10 ;
			data[12541] <= 8'h10 ;
			data[12542] <= 8'h10 ;
			data[12543] <= 8'h10 ;
			data[12544] <= 8'h10 ;
			data[12545] <= 8'h10 ;
			data[12546] <= 8'h10 ;
			data[12547] <= 8'h10 ;
			data[12548] <= 8'h10 ;
			data[12549] <= 8'h10 ;
			data[12550] <= 8'h10 ;
			data[12551] <= 8'h10 ;
			data[12552] <= 8'h10 ;
			data[12553] <= 8'h10 ;
			data[12554] <= 8'h10 ;
			data[12555] <= 8'h10 ;
			data[12556] <= 8'h10 ;
			data[12557] <= 8'h10 ;
			data[12558] <= 8'h10 ;
			data[12559] <= 8'h10 ;
			data[12560] <= 8'h10 ;
			data[12561] <= 8'h10 ;
			data[12562] <= 8'h10 ;
			data[12563] <= 8'h10 ;
			data[12564] <= 8'h10 ;
			data[12565] <= 8'h10 ;
			data[12566] <= 8'h10 ;
			data[12567] <= 8'h10 ;
			data[12568] <= 8'h10 ;
			data[12569] <= 8'h10 ;
			data[12570] <= 8'h10 ;
			data[12571] <= 8'h10 ;
			data[12572] <= 8'h10 ;
			data[12573] <= 8'h10 ;
			data[12574] <= 8'h10 ;
			data[12575] <= 8'h10 ;
			data[12576] <= 8'h10 ;
			data[12577] <= 8'h10 ;
			data[12578] <= 8'h10 ;
			data[12579] <= 8'h10 ;
			data[12580] <= 8'h10 ;
			data[12581] <= 8'h10 ;
			data[12582] <= 8'h10 ;
			data[12583] <= 8'h10 ;
			data[12584] <= 8'h10 ;
			data[12585] <= 8'h10 ;
			data[12586] <= 8'h10 ;
			data[12587] <= 8'h10 ;
			data[12588] <= 8'h10 ;
			data[12589] <= 8'h10 ;
			data[12590] <= 8'h10 ;
			data[12591] <= 8'h10 ;
			data[12592] <= 8'h10 ;
			data[12593] <= 8'h10 ;
			data[12594] <= 8'h10 ;
			data[12595] <= 8'h10 ;
			data[12596] <= 8'h10 ;
			data[12597] <= 8'h10 ;
			data[12598] <= 8'h10 ;
			data[12599] <= 8'h10 ;
			data[12600] <= 8'h10 ;
			data[12601] <= 8'h10 ;
			data[12602] <= 8'h10 ;
			data[12603] <= 8'h10 ;
			data[12604] <= 8'h10 ;
			data[12605] <= 8'h10 ;
			data[12606] <= 8'h10 ;
			data[12607] <= 8'h10 ;
			data[12608] <= 8'h10 ;
			data[12609] <= 8'h10 ;
			data[12610] <= 8'h10 ;
			data[12611] <= 8'h10 ;
			data[12612] <= 8'h10 ;
			data[12613] <= 8'h10 ;
			data[12614] <= 8'h10 ;
			data[12615] <= 8'h10 ;
			data[12616] <= 8'h10 ;
			data[12617] <= 8'h10 ;
			data[12618] <= 8'h10 ;
			data[12619] <= 8'h10 ;
			data[12620] <= 8'h10 ;
			data[12621] <= 8'h10 ;
			data[12622] <= 8'h10 ;
			data[12623] <= 8'h10 ;
			data[12624] <= 8'h10 ;
			data[12625] <= 8'h10 ;
			data[12626] <= 8'h10 ;
			data[12627] <= 8'h10 ;
			data[12628] <= 8'h10 ;
			data[12629] <= 8'h10 ;
			data[12630] <= 8'h10 ;
			data[12631] <= 8'h10 ;
			data[12632] <= 8'h10 ;
			data[12633] <= 8'h10 ;
			data[12634] <= 8'h10 ;
			data[12635] <= 8'h10 ;
			data[12636] <= 8'h10 ;
			data[12637] <= 8'h10 ;
			data[12638] <= 8'h10 ;
			data[12639] <= 8'h10 ;
			data[12640] <= 8'h10 ;
			data[12641] <= 8'h10 ;
			data[12642] <= 8'h10 ;
			data[12643] <= 8'h10 ;
			data[12644] <= 8'h10 ;
			data[12645] <= 8'h10 ;
			data[12646] <= 8'h10 ;
			data[12647] <= 8'h10 ;
			data[12648] <= 8'h10 ;
			data[12649] <= 8'h10 ;
			data[12650] <= 8'h10 ;
			data[12651] <= 8'h10 ;
			data[12652] <= 8'h10 ;
			data[12653] <= 8'h10 ;
			data[12654] <= 8'h10 ;
			data[12655] <= 8'h10 ;
			data[12656] <= 8'h10 ;
			data[12657] <= 8'h10 ;
			data[12658] <= 8'h10 ;
			data[12659] <= 8'h10 ;
			data[12660] <= 8'h10 ;
			data[12661] <= 8'h10 ;
			data[12662] <= 8'h10 ;
			data[12663] <= 8'h10 ;
			data[12664] <= 8'h10 ;
			data[12665] <= 8'h10 ;
			data[12666] <= 8'h10 ;
			data[12667] <= 8'h10 ;
			data[12668] <= 8'h10 ;
			data[12669] <= 8'h10 ;
			data[12670] <= 8'h10 ;
			data[12671] <= 8'h10 ;
			data[12672] <= 8'h10 ;
			data[12673] <= 8'h10 ;
			data[12674] <= 8'h10 ;
			data[12675] <= 8'h10 ;
			data[12676] <= 8'h10 ;
			data[12677] <= 8'h10 ;
			data[12678] <= 8'h10 ;
			data[12679] <= 8'h10 ;
			data[12680] <= 8'h10 ;
			data[12681] <= 8'h10 ;
			data[12682] <= 8'h10 ;
			data[12683] <= 8'h10 ;
			data[12684] <= 8'h10 ;
			data[12685] <= 8'h10 ;
			data[12686] <= 8'h10 ;
			data[12687] <= 8'h10 ;
			data[12688] <= 8'h10 ;
			data[12689] <= 8'h10 ;
			data[12690] <= 8'h10 ;
			data[12691] <= 8'h10 ;
			data[12692] <= 8'h10 ;
			data[12693] <= 8'h10 ;
			data[12694] <= 8'h10 ;
			data[12695] <= 8'h10 ;
			data[12696] <= 8'h10 ;
			data[12697] <= 8'h10 ;
			data[12698] <= 8'h10 ;
			data[12699] <= 8'h10 ;
			data[12700] <= 8'h10 ;
			data[12701] <= 8'h10 ;
			data[12702] <= 8'h10 ;
			data[12703] <= 8'h10 ;
			data[12704] <= 8'h10 ;
			data[12705] <= 8'h10 ;
			data[12706] <= 8'h10 ;
			data[12707] <= 8'h10 ;
			data[12708] <= 8'h10 ;
			data[12709] <= 8'h10 ;
			data[12710] <= 8'h10 ;
			data[12711] <= 8'h10 ;
			data[12712] <= 8'h10 ;
			data[12713] <= 8'h10 ;
			data[12714] <= 8'h10 ;
			data[12715] <= 8'h10 ;
			data[12716] <= 8'h10 ;
			data[12717] <= 8'h10 ;
			data[12718] <= 8'h10 ;
			data[12719] <= 8'h10 ;
			data[12720] <= 8'h10 ;
			data[12721] <= 8'h10 ;
			data[12722] <= 8'h10 ;
			data[12723] <= 8'h10 ;
			data[12724] <= 8'h10 ;
			data[12725] <= 8'h10 ;
			data[12726] <= 8'h10 ;
			data[12727] <= 8'h10 ;
			data[12728] <= 8'h10 ;
			data[12729] <= 8'h10 ;
			data[12730] <= 8'h10 ;
			data[12731] <= 8'h10 ;
			data[12732] <= 8'h10 ;
			data[12733] <= 8'h10 ;
			data[12734] <= 8'h10 ;
			data[12735] <= 8'h10 ;
			data[12736] <= 8'h10 ;
			data[12737] <= 8'h10 ;
			data[12738] <= 8'h10 ;
			data[12739] <= 8'h10 ;
			data[12740] <= 8'h10 ;
			data[12741] <= 8'h10 ;
			data[12742] <= 8'h10 ;
			data[12743] <= 8'h10 ;
			data[12744] <= 8'h10 ;
			data[12745] <= 8'h10 ;
			data[12746] <= 8'h10 ;
			data[12747] <= 8'h10 ;
			data[12748] <= 8'h10 ;
			data[12749] <= 8'h10 ;
			data[12750] <= 8'h10 ;
			data[12751] <= 8'h10 ;
			data[12752] <= 8'h10 ;
			data[12753] <= 8'h10 ;
			data[12754] <= 8'h10 ;
			data[12755] <= 8'h10 ;
			data[12756] <= 8'h10 ;
			data[12757] <= 8'h10 ;
			data[12758] <= 8'h10 ;
			data[12759] <= 8'h10 ;
			data[12760] <= 8'h10 ;
			data[12761] <= 8'h10 ;
			data[12762] <= 8'h10 ;
			data[12763] <= 8'h10 ;
			data[12764] <= 8'h10 ;
			data[12765] <= 8'h10 ;
			data[12766] <= 8'h10 ;
			data[12767] <= 8'h10 ;
			data[12768] <= 8'h10 ;
			data[12769] <= 8'h10 ;
			data[12770] <= 8'h10 ;
			data[12771] <= 8'h10 ;
			data[12772] <= 8'h10 ;
			data[12773] <= 8'h10 ;
			data[12774] <= 8'h10 ;
			data[12775] <= 8'h10 ;
			data[12776] <= 8'h10 ;
			data[12777] <= 8'h10 ;
			data[12778] <= 8'h10 ;
			data[12779] <= 8'h10 ;
			data[12780] <= 8'h10 ;
			data[12781] <= 8'h10 ;
			data[12782] <= 8'h10 ;
			data[12783] <= 8'h10 ;
			data[12784] <= 8'h10 ;
			data[12785] <= 8'h10 ;
			data[12786] <= 8'h10 ;
			data[12787] <= 8'h10 ;
			data[12788] <= 8'h10 ;
			data[12789] <= 8'h10 ;
			data[12790] <= 8'h10 ;
			data[12791] <= 8'h10 ;
			data[12792] <= 8'h10 ;
			data[12793] <= 8'h10 ;
			data[12794] <= 8'h10 ;
			data[12795] <= 8'h10 ;
			data[12796] <= 8'h10 ;
			data[12797] <= 8'h10 ;
			data[12798] <= 8'h10 ;
			data[12799] <= 8'h10 ;
			data[12800] <= 8'h10 ;
			data[12801] <= 8'h10 ;
			data[12802] <= 8'h10 ;
			data[12803] <= 8'h10 ;
			data[12804] <= 8'h10 ;
			data[12805] <= 8'h10 ;
			data[12806] <= 8'h10 ;
			data[12807] <= 8'h10 ;
			data[12808] <= 8'h10 ;
			data[12809] <= 8'h10 ;
			data[12810] <= 8'h10 ;
			data[12811] <= 8'h10 ;
			data[12812] <= 8'h10 ;
			data[12813] <= 8'h10 ;
			data[12814] <= 8'h10 ;
			data[12815] <= 8'h10 ;
			data[12816] <= 8'h10 ;
			data[12817] <= 8'h10 ;
			data[12818] <= 8'h10 ;
			data[12819] <= 8'h10 ;
			data[12820] <= 8'h10 ;
			data[12821] <= 8'h10 ;
			data[12822] <= 8'h10 ;
			data[12823] <= 8'h10 ;
			data[12824] <= 8'h10 ;
			data[12825] <= 8'h10 ;
			data[12826] <= 8'h10 ;
			data[12827] <= 8'h10 ;
			data[12828] <= 8'h10 ;
			data[12829] <= 8'h10 ;
			data[12830] <= 8'h10 ;
			data[12831] <= 8'h10 ;
			data[12832] <= 8'h10 ;
			data[12833] <= 8'h10 ;
			data[12834] <= 8'h10 ;
			data[12835] <= 8'h10 ;
			data[12836] <= 8'h10 ;
			data[12837] <= 8'h10 ;
			data[12838] <= 8'h10 ;
			data[12839] <= 8'h10 ;
			data[12840] <= 8'h10 ;
			data[12841] <= 8'h10 ;
			data[12842] <= 8'h10 ;
			data[12843] <= 8'h10 ;
			data[12844] <= 8'h10 ;
			data[12845] <= 8'h10 ;
			data[12846] <= 8'h10 ;
			data[12847] <= 8'h10 ;
			data[12848] <= 8'h10 ;
			data[12849] <= 8'h10 ;
			data[12850] <= 8'h10 ;
			data[12851] <= 8'h10 ;
			data[12852] <= 8'h10 ;
			data[12853] <= 8'h10 ;
			data[12854] <= 8'h10 ;
			data[12855] <= 8'h10 ;
			data[12856] <= 8'h10 ;
			data[12857] <= 8'h10 ;
			data[12858] <= 8'h10 ;
			data[12859] <= 8'h10 ;
			data[12860] <= 8'h10 ;
			data[12861] <= 8'h10 ;
			data[12862] <= 8'h10 ;
			data[12863] <= 8'h10 ;
			data[12864] <= 8'h10 ;
			data[12865] <= 8'h10 ;
			data[12866] <= 8'h10 ;
			data[12867] <= 8'h10 ;
			data[12868] <= 8'h10 ;
			data[12869] <= 8'h10 ;
			data[12870] <= 8'h10 ;
			data[12871] <= 8'h10 ;
			data[12872] <= 8'h10 ;
			data[12873] <= 8'h10 ;
			data[12874] <= 8'h10 ;
			data[12875] <= 8'h10 ;
			data[12876] <= 8'h10 ;
			data[12877] <= 8'h10 ;
			data[12878] <= 8'h10 ;
			data[12879] <= 8'h10 ;
			data[12880] <= 8'h10 ;
			data[12881] <= 8'h10 ;
			data[12882] <= 8'h10 ;
			data[12883] <= 8'h10 ;
			data[12884] <= 8'h10 ;
			data[12885] <= 8'h10 ;
			data[12886] <= 8'h10 ;
			data[12887] <= 8'h10 ;
			data[12888] <= 8'h10 ;
			data[12889] <= 8'h10 ;
			data[12890] <= 8'h10 ;
			data[12891] <= 8'h10 ;
			data[12892] <= 8'h10 ;
			data[12893] <= 8'h10 ;
			data[12894] <= 8'h10 ;
			data[12895] <= 8'h10 ;
			data[12896] <= 8'h10 ;
			data[12897] <= 8'h10 ;
			data[12898] <= 8'h10 ;
			data[12899] <= 8'h10 ;
			data[12900] <= 8'h10 ;
			data[12901] <= 8'h10 ;
			data[12902] <= 8'h10 ;
			data[12903] <= 8'h10 ;
			data[12904] <= 8'h10 ;
			data[12905] <= 8'h10 ;
			data[12906] <= 8'h10 ;
			data[12907] <= 8'h10 ;
			data[12908] <= 8'h10 ;
			data[12909] <= 8'h10 ;
			data[12910] <= 8'h10 ;
			data[12911] <= 8'h10 ;
			data[12912] <= 8'h10 ;
			data[12913] <= 8'h10 ;
			data[12914] <= 8'h10 ;
			data[12915] <= 8'h10 ;
			data[12916] <= 8'h10 ;
			data[12917] <= 8'h10 ;
			data[12918] <= 8'h10 ;
			data[12919] <= 8'h10 ;
			data[12920] <= 8'h10 ;
			data[12921] <= 8'h10 ;
			data[12922] <= 8'h10 ;
			data[12923] <= 8'h10 ;
			data[12924] <= 8'h10 ;
			data[12925] <= 8'h10 ;
			data[12926] <= 8'h10 ;
			data[12927] <= 8'h10 ;
			data[12928] <= 8'h10 ;
			data[12929] <= 8'h10 ;
			data[12930] <= 8'h10 ;
			data[12931] <= 8'h10 ;
			data[12932] <= 8'h10 ;
			data[12933] <= 8'h10 ;
			data[12934] <= 8'h10 ;
			data[12935] <= 8'h10 ;
			data[12936] <= 8'h10 ;
			data[12937] <= 8'h10 ;
			data[12938] <= 8'h10 ;
			data[12939] <= 8'h10 ;
			data[12940] <= 8'h10 ;
			data[12941] <= 8'h10 ;
			data[12942] <= 8'h10 ;
			data[12943] <= 8'h10 ;
			data[12944] <= 8'h10 ;
			data[12945] <= 8'h10 ;
			data[12946] <= 8'h10 ;
			data[12947] <= 8'h10 ;
			data[12948] <= 8'h10 ;
			data[12949] <= 8'h10 ;
			data[12950] <= 8'h10 ;
			data[12951] <= 8'h10 ;
			data[12952] <= 8'h10 ;
			data[12953] <= 8'h10 ;
			data[12954] <= 8'h10 ;
			data[12955] <= 8'h10 ;
			data[12956] <= 8'h10 ;
			data[12957] <= 8'h10 ;
			data[12958] <= 8'h10 ;
			data[12959] <= 8'h10 ;
			data[12960] <= 8'h10 ;
			data[12961] <= 8'h10 ;
			data[12962] <= 8'h10 ;
			data[12963] <= 8'h10 ;
			data[12964] <= 8'h10 ;
			data[12965] <= 8'h10 ;
			data[12966] <= 8'h10 ;
			data[12967] <= 8'h10 ;
			data[12968] <= 8'h10 ;
			data[12969] <= 8'h10 ;
			data[12970] <= 8'h10 ;
			data[12971] <= 8'h10 ;
			data[12972] <= 8'h10 ;
			data[12973] <= 8'h10 ;
			data[12974] <= 8'h10 ;
			data[12975] <= 8'h10 ;
			data[12976] <= 8'h10 ;
			data[12977] <= 8'h10 ;
			data[12978] <= 8'h10 ;
			data[12979] <= 8'h10 ;
			data[12980] <= 8'h10 ;
			data[12981] <= 8'h10 ;
			data[12982] <= 8'h10 ;
			data[12983] <= 8'h10 ;
			data[12984] <= 8'h10 ;
			data[12985] <= 8'h10 ;
			data[12986] <= 8'h10 ;
			data[12987] <= 8'h10 ;
			data[12988] <= 8'h10 ;
			data[12989] <= 8'h10 ;
			data[12990] <= 8'h10 ;
			data[12991] <= 8'h10 ;
			data[12992] <= 8'h10 ;
			data[12993] <= 8'h10 ;
			data[12994] <= 8'h10 ;
			data[12995] <= 8'h10 ;
			data[12996] <= 8'h10 ;
			data[12997] <= 8'h10 ;
			data[12998] <= 8'h10 ;
			data[12999] <= 8'h10 ;
			data[13000] <= 8'h10 ;
			data[13001] <= 8'h10 ;
			data[13002] <= 8'h10 ;
			data[13003] <= 8'h10 ;
			data[13004] <= 8'h10 ;
			data[13005] <= 8'h10 ;
			data[13006] <= 8'h10 ;
			data[13007] <= 8'h10 ;
			data[13008] <= 8'h10 ;
			data[13009] <= 8'h10 ;
			data[13010] <= 8'h10 ;
			data[13011] <= 8'h10 ;
			data[13012] <= 8'h10 ;
			data[13013] <= 8'h10 ;
			data[13014] <= 8'h10 ;
			data[13015] <= 8'h10 ;
			data[13016] <= 8'h10 ;
			data[13017] <= 8'h10 ;
			data[13018] <= 8'h10 ;
			data[13019] <= 8'h10 ;
			data[13020] <= 8'h10 ;
			data[13021] <= 8'h10 ;
			data[13022] <= 8'h10 ;
			data[13023] <= 8'h10 ;
			data[13024] <= 8'h10 ;
			data[13025] <= 8'h10 ;
			data[13026] <= 8'h10 ;
			data[13027] <= 8'h10 ;
			data[13028] <= 8'h10 ;
			data[13029] <= 8'h10 ;
			data[13030] <= 8'h10 ;
			data[13031] <= 8'h10 ;
			data[13032] <= 8'h10 ;
			data[13033] <= 8'h10 ;
			data[13034] <= 8'h10 ;
			data[13035] <= 8'h10 ;
			data[13036] <= 8'h10 ;
			data[13037] <= 8'h10 ;
			data[13038] <= 8'h10 ;
			data[13039] <= 8'h10 ;
			data[13040] <= 8'h10 ;
			data[13041] <= 8'h10 ;
			data[13042] <= 8'h10 ;
			data[13043] <= 8'h10 ;
			data[13044] <= 8'h10 ;
			data[13045] <= 8'h10 ;
			data[13046] <= 8'h10 ;
			data[13047] <= 8'h10 ;
			data[13048] <= 8'h10 ;
			data[13049] <= 8'h10 ;
			data[13050] <= 8'h10 ;
			data[13051] <= 8'h10 ;
			data[13052] <= 8'h10 ;
			data[13053] <= 8'h10 ;
			data[13054] <= 8'h10 ;
			data[13055] <= 8'h10 ;
			data[13056] <= 8'h10 ;
			data[13057] <= 8'h10 ;
			data[13058] <= 8'h10 ;
			data[13059] <= 8'h10 ;
			data[13060] <= 8'h10 ;
			data[13061] <= 8'h10 ;
			data[13062] <= 8'h10 ;
			data[13063] <= 8'h10 ;
			data[13064] <= 8'h10 ;
			data[13065] <= 8'h10 ;
			data[13066] <= 8'h10 ;
			data[13067] <= 8'h10 ;
			data[13068] <= 8'h10 ;
			data[13069] <= 8'h10 ;
			data[13070] <= 8'h10 ;
			data[13071] <= 8'h10 ;
			data[13072] <= 8'h10 ;
			data[13073] <= 8'h10 ;
			data[13074] <= 8'h10 ;
			data[13075] <= 8'h10 ;
			data[13076] <= 8'h10 ;
			data[13077] <= 8'h10 ;
			data[13078] <= 8'h10 ;
			data[13079] <= 8'h10 ;
			data[13080] <= 8'h10 ;
			data[13081] <= 8'h10 ;
			data[13082] <= 8'h10 ;
			data[13083] <= 8'h10 ;
			data[13084] <= 8'h10 ;
			data[13085] <= 8'h10 ;
			data[13086] <= 8'h10 ;
			data[13087] <= 8'h10 ;
			data[13088] <= 8'h10 ;
			data[13089] <= 8'h10 ;
			data[13090] <= 8'h10 ;
			data[13091] <= 8'h10 ;
			data[13092] <= 8'h10 ;
			data[13093] <= 8'h10 ;
			data[13094] <= 8'h10 ;
			data[13095] <= 8'h10 ;
			data[13096] <= 8'h10 ;
			data[13097] <= 8'h10 ;
			data[13098] <= 8'h10 ;
			data[13099] <= 8'h10 ;
			data[13100] <= 8'h10 ;
			data[13101] <= 8'h10 ;
			data[13102] <= 8'h10 ;
			data[13103] <= 8'h10 ;
			data[13104] <= 8'h10 ;
			data[13105] <= 8'h10 ;
			data[13106] <= 8'h10 ;
			data[13107] <= 8'h10 ;
			data[13108] <= 8'h10 ;
			data[13109] <= 8'h10 ;
			data[13110] <= 8'h10 ;
			data[13111] <= 8'h10 ;
			data[13112] <= 8'h10 ;
			data[13113] <= 8'h10 ;
			data[13114] <= 8'h10 ;
			data[13115] <= 8'h10 ;
			data[13116] <= 8'h10 ;
			data[13117] <= 8'h10 ;
			data[13118] <= 8'h10 ;
			data[13119] <= 8'h10 ;
			data[13120] <= 8'h10 ;
			data[13121] <= 8'h10 ;
			data[13122] <= 8'h10 ;
			data[13123] <= 8'h10 ;
			data[13124] <= 8'h10 ;
			data[13125] <= 8'h10 ;
			data[13126] <= 8'h10 ;
			data[13127] <= 8'h10 ;
			data[13128] <= 8'h10 ;
			data[13129] <= 8'h10 ;
			data[13130] <= 8'h10 ;
			data[13131] <= 8'h10 ;
			data[13132] <= 8'h10 ;
			data[13133] <= 8'h10 ;
			data[13134] <= 8'h10 ;
			data[13135] <= 8'h10 ;
			data[13136] <= 8'h10 ;
			data[13137] <= 8'h10 ;
			data[13138] <= 8'h10 ;
			data[13139] <= 8'h10 ;
			data[13140] <= 8'h10 ;
			data[13141] <= 8'h10 ;
			data[13142] <= 8'h10 ;
			data[13143] <= 8'h10 ;
			data[13144] <= 8'h10 ;
			data[13145] <= 8'h10 ;
			data[13146] <= 8'h10 ;
			data[13147] <= 8'h10 ;
			data[13148] <= 8'h10 ;
			data[13149] <= 8'h10 ;
			data[13150] <= 8'h10 ;
			data[13151] <= 8'h10 ;
			data[13152] <= 8'h10 ;
			data[13153] <= 8'h10 ;
			data[13154] <= 8'h10 ;
			data[13155] <= 8'h10 ;
			data[13156] <= 8'h10 ;
			data[13157] <= 8'h10 ;
			data[13158] <= 8'h10 ;
			data[13159] <= 8'h10 ;
			data[13160] <= 8'h10 ;
			data[13161] <= 8'h10 ;
			data[13162] <= 8'h10 ;
			data[13163] <= 8'h10 ;
			data[13164] <= 8'h10 ;
			data[13165] <= 8'h10 ;
			data[13166] <= 8'h10 ;
			data[13167] <= 8'h10 ;
			data[13168] <= 8'h10 ;
			data[13169] <= 8'h10 ;
			data[13170] <= 8'h10 ;
			data[13171] <= 8'h10 ;
			data[13172] <= 8'h10 ;
			data[13173] <= 8'h10 ;
			data[13174] <= 8'h10 ;
			data[13175] <= 8'h10 ;
			data[13176] <= 8'h10 ;
			data[13177] <= 8'h10 ;
			data[13178] <= 8'h10 ;
			data[13179] <= 8'h10 ;
			data[13180] <= 8'h10 ;
			data[13181] <= 8'h10 ;
			data[13182] <= 8'h10 ;
			data[13183] <= 8'h10 ;
			data[13184] <= 8'h10 ;
			data[13185] <= 8'h10 ;
			data[13186] <= 8'h10 ;
			data[13187] <= 8'h10 ;
			data[13188] <= 8'h10 ;
			data[13189] <= 8'h10 ;
			data[13190] <= 8'h10 ;
			data[13191] <= 8'h10 ;
			data[13192] <= 8'h10 ;
			data[13193] <= 8'h10 ;
			data[13194] <= 8'h10 ;
			data[13195] <= 8'h10 ;
			data[13196] <= 8'h10 ;
			data[13197] <= 8'h10 ;
			data[13198] <= 8'h10 ;
			data[13199] <= 8'h10 ;
			data[13200] <= 8'h10 ;
			data[13201] <= 8'h10 ;
			data[13202] <= 8'h10 ;
			data[13203] <= 8'h10 ;
			data[13204] <= 8'h10 ;
			data[13205] <= 8'h10 ;
			data[13206] <= 8'h10 ;
			data[13207] <= 8'h10 ;
			data[13208] <= 8'h10 ;
			data[13209] <= 8'h10 ;
			data[13210] <= 8'h10 ;
			data[13211] <= 8'h10 ;
			data[13212] <= 8'h10 ;
			data[13213] <= 8'h10 ;
			data[13214] <= 8'h10 ;
			data[13215] <= 8'h10 ;
			data[13216] <= 8'h10 ;
			data[13217] <= 8'h10 ;
			data[13218] <= 8'h10 ;
			data[13219] <= 8'h10 ;
			data[13220] <= 8'h10 ;
			data[13221] <= 8'h10 ;
			data[13222] <= 8'h10 ;
			data[13223] <= 8'h10 ;
			data[13224] <= 8'h10 ;
			data[13225] <= 8'h10 ;
			data[13226] <= 8'h10 ;
			data[13227] <= 8'h10 ;
			data[13228] <= 8'h10 ;
			data[13229] <= 8'h10 ;
			data[13230] <= 8'h10 ;
			data[13231] <= 8'h10 ;
			data[13232] <= 8'h10 ;
			data[13233] <= 8'h10 ;
			data[13234] <= 8'h10 ;
			data[13235] <= 8'h10 ;
			data[13236] <= 8'h10 ;
			data[13237] <= 8'h10 ;
			data[13238] <= 8'h10 ;
			data[13239] <= 8'h10 ;
			data[13240] <= 8'h10 ;
			data[13241] <= 8'h10 ;
			data[13242] <= 8'h10 ;
			data[13243] <= 8'h10 ;
			data[13244] <= 8'h10 ;
			data[13245] <= 8'h10 ;
			data[13246] <= 8'h10 ;
			data[13247] <= 8'h10 ;
			data[13248] <= 8'h10 ;
			data[13249] <= 8'h10 ;
			data[13250] <= 8'h10 ;
			data[13251] <= 8'h10 ;
			data[13252] <= 8'h10 ;
			data[13253] <= 8'h10 ;
			data[13254] <= 8'h10 ;
			data[13255] <= 8'h10 ;
			data[13256] <= 8'h10 ;
			data[13257] <= 8'h10 ;
			data[13258] <= 8'h10 ;
			data[13259] <= 8'h10 ;
			data[13260] <= 8'h10 ;
			data[13261] <= 8'h10 ;
			data[13262] <= 8'h10 ;
			data[13263] <= 8'h10 ;
			data[13264] <= 8'h10 ;
			data[13265] <= 8'h10 ;
			data[13266] <= 8'h10 ;
			data[13267] <= 8'h10 ;
			data[13268] <= 8'h10 ;
			data[13269] <= 8'h10 ;
			data[13270] <= 8'h10 ;
			data[13271] <= 8'h10 ;
			data[13272] <= 8'h10 ;
			data[13273] <= 8'h10 ;
			data[13274] <= 8'h10 ;
			data[13275] <= 8'h10 ;
			data[13276] <= 8'h10 ;
			data[13277] <= 8'h10 ;
			data[13278] <= 8'h10 ;
			data[13279] <= 8'h10 ;
			data[13280] <= 8'h10 ;
			data[13281] <= 8'h10 ;
			data[13282] <= 8'h10 ;
			data[13283] <= 8'h10 ;
			data[13284] <= 8'h10 ;
			data[13285] <= 8'h10 ;
			data[13286] <= 8'h10 ;
			data[13287] <= 8'h10 ;
			data[13288] <= 8'h10 ;
			data[13289] <= 8'h10 ;
			data[13290] <= 8'h10 ;
			data[13291] <= 8'h10 ;
			data[13292] <= 8'h10 ;
			data[13293] <= 8'h10 ;
			data[13294] <= 8'h10 ;
			data[13295] <= 8'h10 ;
			data[13296] <= 8'h10 ;
			data[13297] <= 8'h10 ;
			data[13298] <= 8'h10 ;
			data[13299] <= 8'h10 ;
			data[13300] <= 8'h10 ;
			data[13301] <= 8'h10 ;
			data[13302] <= 8'h10 ;
			data[13303] <= 8'h10 ;
			data[13304] <= 8'h10 ;
			data[13305] <= 8'h10 ;
			data[13306] <= 8'h10 ;
			data[13307] <= 8'h10 ;
			data[13308] <= 8'h10 ;
			data[13309] <= 8'h10 ;
			data[13310] <= 8'h10 ;
			data[13311] <= 8'h10 ;
			data[13312] <= 8'h10 ;
			data[13313] <= 8'h10 ;
			data[13314] <= 8'h10 ;
			data[13315] <= 8'h10 ;
			data[13316] <= 8'h10 ;
			data[13317] <= 8'h10 ;
			data[13318] <= 8'h10 ;
			data[13319] <= 8'h10 ;
			data[13320] <= 8'h10 ;
			data[13321] <= 8'h10 ;
			data[13322] <= 8'h10 ;
			data[13323] <= 8'h10 ;
			data[13324] <= 8'h10 ;
			data[13325] <= 8'h10 ;
			data[13326] <= 8'h10 ;
			data[13327] <= 8'h10 ;
			data[13328] <= 8'h10 ;
			data[13329] <= 8'h10 ;
			data[13330] <= 8'h10 ;
			data[13331] <= 8'h10 ;
			data[13332] <= 8'h10 ;
			data[13333] <= 8'h10 ;
			data[13334] <= 8'h10 ;
			data[13335] <= 8'h10 ;
			data[13336] <= 8'h10 ;
			data[13337] <= 8'h10 ;
			data[13338] <= 8'h10 ;
			data[13339] <= 8'h10 ;
			data[13340] <= 8'h10 ;
			data[13341] <= 8'h10 ;
			data[13342] <= 8'h10 ;
			data[13343] <= 8'h10 ;
			data[13344] <= 8'h10 ;
			data[13345] <= 8'h10 ;
			data[13346] <= 8'h10 ;
			data[13347] <= 8'h10 ;
			data[13348] <= 8'h10 ;
			data[13349] <= 8'h10 ;
			data[13350] <= 8'h10 ;
			data[13351] <= 8'h10 ;
			data[13352] <= 8'h10 ;
			data[13353] <= 8'h10 ;
			data[13354] <= 8'h10 ;
			data[13355] <= 8'h10 ;
			data[13356] <= 8'h10 ;
			data[13357] <= 8'h10 ;
			data[13358] <= 8'h10 ;
			data[13359] <= 8'h10 ;
			data[13360] <= 8'h10 ;
			data[13361] <= 8'h10 ;
			data[13362] <= 8'h10 ;
			data[13363] <= 8'h10 ;
			data[13364] <= 8'h10 ;
			data[13365] <= 8'h10 ;
			data[13366] <= 8'h10 ;
			data[13367] <= 8'h10 ;
			data[13368] <= 8'h10 ;
			data[13369] <= 8'h10 ;
			data[13370] <= 8'h10 ;
			data[13371] <= 8'h10 ;
			data[13372] <= 8'h10 ;
			data[13373] <= 8'h10 ;
			data[13374] <= 8'h10 ;
			data[13375] <= 8'h10 ;
			data[13376] <= 8'h10 ;
			data[13377] <= 8'h10 ;
			data[13378] <= 8'h10 ;
			data[13379] <= 8'h10 ;
			data[13380] <= 8'h10 ;
			data[13381] <= 8'h10 ;
			data[13382] <= 8'h10 ;
			data[13383] <= 8'h10 ;
			data[13384] <= 8'h10 ;
			data[13385] <= 8'h10 ;
			data[13386] <= 8'h10 ;
			data[13387] <= 8'h10 ;
			data[13388] <= 8'h10 ;
			data[13389] <= 8'h10 ;
			data[13390] <= 8'h10 ;
			data[13391] <= 8'h10 ;
			data[13392] <= 8'h10 ;
			data[13393] <= 8'h10 ;
			data[13394] <= 8'h10 ;
			data[13395] <= 8'h10 ;
			data[13396] <= 8'h10 ;
			data[13397] <= 8'h10 ;
			data[13398] <= 8'h10 ;
			data[13399] <= 8'h10 ;
			data[13400] <= 8'h10 ;
			data[13401] <= 8'h10 ;
			data[13402] <= 8'h10 ;
			data[13403] <= 8'h10 ;
			data[13404] <= 8'h10 ;
			data[13405] <= 8'h10 ;
			data[13406] <= 8'h10 ;
			data[13407] <= 8'h10 ;
			data[13408] <= 8'h10 ;
			data[13409] <= 8'h10 ;
			data[13410] <= 8'h10 ;
			data[13411] <= 8'h10 ;
			data[13412] <= 8'h10 ;
			data[13413] <= 8'h10 ;
			data[13414] <= 8'h10 ;
			data[13415] <= 8'h10 ;
			data[13416] <= 8'h10 ;
			data[13417] <= 8'h10 ;
			data[13418] <= 8'h10 ;
			data[13419] <= 8'h10 ;
			data[13420] <= 8'h10 ;
			data[13421] <= 8'h10 ;
			data[13422] <= 8'h10 ;
			data[13423] <= 8'h10 ;
			data[13424] <= 8'h10 ;
			data[13425] <= 8'h10 ;
			data[13426] <= 8'h10 ;
			data[13427] <= 8'h10 ;
			data[13428] <= 8'h10 ;
			data[13429] <= 8'h10 ;
			data[13430] <= 8'h10 ;
			data[13431] <= 8'h10 ;
			data[13432] <= 8'h10 ;
			data[13433] <= 8'h10 ;
			data[13434] <= 8'h10 ;
			data[13435] <= 8'h10 ;
			data[13436] <= 8'h10 ;
			data[13437] <= 8'h10 ;
			data[13438] <= 8'h10 ;
			data[13439] <= 8'h10 ;
			data[13440] <= 8'h10 ;
			data[13441] <= 8'h10 ;
			data[13442] <= 8'h10 ;
			data[13443] <= 8'h10 ;
			data[13444] <= 8'h10 ;
			data[13445] <= 8'h10 ;
			data[13446] <= 8'h10 ;
			data[13447] <= 8'h10 ;
			data[13448] <= 8'h10 ;
			data[13449] <= 8'h10 ;
			data[13450] <= 8'h10 ;
			data[13451] <= 8'h10 ;
			data[13452] <= 8'h10 ;
			data[13453] <= 8'h10 ;
			data[13454] <= 8'h10 ;
			data[13455] <= 8'h10 ;
			data[13456] <= 8'h10 ;
			data[13457] <= 8'h10 ;
			data[13458] <= 8'h10 ;
			data[13459] <= 8'h10 ;
			data[13460] <= 8'h10 ;
			data[13461] <= 8'h10 ;
			data[13462] <= 8'h10 ;
			data[13463] <= 8'h10 ;
			data[13464] <= 8'h10 ;
			data[13465] <= 8'h10 ;
			data[13466] <= 8'h10 ;
			data[13467] <= 8'h10 ;
			data[13468] <= 8'h10 ;
			data[13469] <= 8'h10 ;
			data[13470] <= 8'h10 ;
			data[13471] <= 8'h10 ;
			data[13472] <= 8'h10 ;
			data[13473] <= 8'h10 ;
			data[13474] <= 8'h10 ;
			data[13475] <= 8'h10 ;
			data[13476] <= 8'h10 ;
			data[13477] <= 8'h10 ;
			data[13478] <= 8'h10 ;
			data[13479] <= 8'h10 ;
			data[13480] <= 8'h10 ;
			data[13481] <= 8'h10 ;
			data[13482] <= 8'h10 ;
			data[13483] <= 8'h10 ;
			data[13484] <= 8'h10 ;
			data[13485] <= 8'h10 ;
			data[13486] <= 8'h10 ;
			data[13487] <= 8'h10 ;
			data[13488] <= 8'h10 ;
			data[13489] <= 8'h10 ;
			data[13490] <= 8'h10 ;
			data[13491] <= 8'h10 ;
			data[13492] <= 8'h10 ;
			data[13493] <= 8'h10 ;
			data[13494] <= 8'h10 ;
			data[13495] <= 8'h10 ;
			data[13496] <= 8'h10 ;
			data[13497] <= 8'h10 ;
			data[13498] <= 8'h10 ;
			data[13499] <= 8'h10 ;
			data[13500] <= 8'h10 ;
			data[13501] <= 8'h10 ;
			data[13502] <= 8'h10 ;
			data[13503] <= 8'h10 ;
			data[13504] <= 8'h10 ;
			data[13505] <= 8'h10 ;
			data[13506] <= 8'h10 ;
			data[13507] <= 8'h10 ;
			data[13508] <= 8'h10 ;
			data[13509] <= 8'h10 ;
			data[13510] <= 8'h10 ;
			data[13511] <= 8'h10 ;
			data[13512] <= 8'h10 ;
			data[13513] <= 8'h10 ;
			data[13514] <= 8'h10 ;
			data[13515] <= 8'h10 ;
			data[13516] <= 8'h10 ;
			data[13517] <= 8'h10 ;
			data[13518] <= 8'h10 ;
			data[13519] <= 8'h10 ;
			data[13520] <= 8'h10 ;
			data[13521] <= 8'h10 ;
			data[13522] <= 8'h10 ;
			data[13523] <= 8'h10 ;
			data[13524] <= 8'h10 ;
			data[13525] <= 8'h10 ;
			data[13526] <= 8'h10 ;
			data[13527] <= 8'h10 ;
			data[13528] <= 8'h10 ;
			data[13529] <= 8'h10 ;
			data[13530] <= 8'h10 ;
			data[13531] <= 8'h10 ;
			data[13532] <= 8'h10 ;
			data[13533] <= 8'h10 ;
			data[13534] <= 8'h10 ;
			data[13535] <= 8'h10 ;
			data[13536] <= 8'h10 ;
			data[13537] <= 8'h10 ;
			data[13538] <= 8'h10 ;
			data[13539] <= 8'h10 ;
			data[13540] <= 8'h10 ;
			data[13541] <= 8'h10 ;
			data[13542] <= 8'h10 ;
			data[13543] <= 8'h10 ;
			data[13544] <= 8'h10 ;
			data[13545] <= 8'h10 ;
			data[13546] <= 8'h10 ;
			data[13547] <= 8'h10 ;
			data[13548] <= 8'h10 ;
			data[13549] <= 8'h10 ;
			data[13550] <= 8'h10 ;
			data[13551] <= 8'h10 ;
			data[13552] <= 8'h10 ;
			data[13553] <= 8'h10 ;
			data[13554] <= 8'h10 ;
			data[13555] <= 8'h10 ;
			data[13556] <= 8'h10 ;
			data[13557] <= 8'h10 ;
			data[13558] <= 8'h10 ;
			data[13559] <= 8'h10 ;
			data[13560] <= 8'h10 ;
			data[13561] <= 8'h10 ;
			data[13562] <= 8'h10 ;
			data[13563] <= 8'h10 ;
			data[13564] <= 8'h10 ;
			data[13565] <= 8'h10 ;
			data[13566] <= 8'h10 ;
			data[13567] <= 8'h10 ;
			data[13568] <= 8'h10 ;
			data[13569] <= 8'h10 ;
			data[13570] <= 8'h10 ;
			data[13571] <= 8'h10 ;
			data[13572] <= 8'h10 ;
			data[13573] <= 8'h10 ;
			data[13574] <= 8'h10 ;
			data[13575] <= 8'h10 ;
			data[13576] <= 8'h10 ;
			data[13577] <= 8'h10 ;
			data[13578] <= 8'h10 ;
			data[13579] <= 8'h10 ;
			data[13580] <= 8'h10 ;
			data[13581] <= 8'h10 ;
			data[13582] <= 8'h10 ;
			data[13583] <= 8'h10 ;
			data[13584] <= 8'h10 ;
			data[13585] <= 8'h10 ;
			data[13586] <= 8'h10 ;
			data[13587] <= 8'h10 ;
			data[13588] <= 8'h10 ;
			data[13589] <= 8'h10 ;
			data[13590] <= 8'h10 ;
			data[13591] <= 8'h10 ;
			data[13592] <= 8'h10 ;
			data[13593] <= 8'h10 ;
			data[13594] <= 8'h10 ;
			data[13595] <= 8'h10 ;
			data[13596] <= 8'h10 ;
			data[13597] <= 8'h10 ;
			data[13598] <= 8'h10 ;
			data[13599] <= 8'h10 ;
			data[13600] <= 8'h10 ;
			data[13601] <= 8'h10 ;
			data[13602] <= 8'h10 ;
			data[13603] <= 8'h10 ;
			data[13604] <= 8'h10 ;
			data[13605] <= 8'h10 ;
			data[13606] <= 8'h10 ;
			data[13607] <= 8'h10 ;
			data[13608] <= 8'h10 ;
			data[13609] <= 8'h10 ;
			data[13610] <= 8'h10 ;
			data[13611] <= 8'h10 ;
			data[13612] <= 8'h10 ;
			data[13613] <= 8'h10 ;
			data[13614] <= 8'h10 ;
			data[13615] <= 8'h10 ;
			data[13616] <= 8'h10 ;
			data[13617] <= 8'h10 ;
			data[13618] <= 8'h10 ;
			data[13619] <= 8'h10 ;
			data[13620] <= 8'h10 ;
			data[13621] <= 8'h10 ;
			data[13622] <= 8'h10 ;
			data[13623] <= 8'h10 ;
			data[13624] <= 8'h10 ;
			data[13625] <= 8'h10 ;
			data[13626] <= 8'h10 ;
			data[13627] <= 8'h10 ;
			data[13628] <= 8'h10 ;
			data[13629] <= 8'h10 ;
			data[13630] <= 8'h10 ;
			data[13631] <= 8'h10 ;
			data[13632] <= 8'h10 ;
			data[13633] <= 8'h10 ;
			data[13634] <= 8'h10 ;
			data[13635] <= 8'h10 ;
			data[13636] <= 8'h10 ;
			data[13637] <= 8'h10 ;
			data[13638] <= 8'h10 ;
			data[13639] <= 8'h10 ;
			data[13640] <= 8'h10 ;
			data[13641] <= 8'h10 ;
			data[13642] <= 8'h10 ;
			data[13643] <= 8'h10 ;
			data[13644] <= 8'h10 ;
			data[13645] <= 8'h10 ;
			data[13646] <= 8'h10 ;
			data[13647] <= 8'h10 ;
			data[13648] <= 8'h10 ;
			data[13649] <= 8'h10 ;
			data[13650] <= 8'h10 ;
			data[13651] <= 8'h10 ;
			data[13652] <= 8'h10 ;
			data[13653] <= 8'h10 ;
			data[13654] <= 8'h10 ;
			data[13655] <= 8'h10 ;
			data[13656] <= 8'h10 ;
			data[13657] <= 8'h10 ;
			data[13658] <= 8'h10 ;
			data[13659] <= 8'h10 ;
			data[13660] <= 8'h10 ;
			data[13661] <= 8'h10 ;
			data[13662] <= 8'h10 ;
			data[13663] <= 8'h10 ;
			data[13664] <= 8'h10 ;
			data[13665] <= 8'h10 ;
			data[13666] <= 8'h10 ;
			data[13667] <= 8'h10 ;
			data[13668] <= 8'h10 ;
			data[13669] <= 8'h10 ;
			data[13670] <= 8'h10 ;
			data[13671] <= 8'h10 ;
			data[13672] <= 8'h10 ;
			data[13673] <= 8'h10 ;
			data[13674] <= 8'h10 ;
			data[13675] <= 8'h10 ;
			data[13676] <= 8'h10 ;
			data[13677] <= 8'h10 ;
			data[13678] <= 8'h10 ;
			data[13679] <= 8'h10 ;
			data[13680] <= 8'h10 ;
			data[13681] <= 8'h10 ;
			data[13682] <= 8'h10 ;
			data[13683] <= 8'h10 ;
			data[13684] <= 8'h10 ;
			data[13685] <= 8'h10 ;
			data[13686] <= 8'h10 ;
			data[13687] <= 8'h10 ;
			data[13688] <= 8'h10 ;
			data[13689] <= 8'h10 ;
			data[13690] <= 8'h10 ;
			data[13691] <= 8'h10 ;
			data[13692] <= 8'h10 ;
			data[13693] <= 8'h10 ;
			data[13694] <= 8'h10 ;
			data[13695] <= 8'h10 ;
			data[13696] <= 8'h10 ;
			data[13697] <= 8'h10 ;
			data[13698] <= 8'h10 ;
			data[13699] <= 8'h10 ;
			data[13700] <= 8'h10 ;
			data[13701] <= 8'h10 ;
			data[13702] <= 8'h10 ;
			data[13703] <= 8'h10 ;
			data[13704] <= 8'h10 ;
			data[13705] <= 8'h10 ;
			data[13706] <= 8'h10 ;
			data[13707] <= 8'h10 ;
			data[13708] <= 8'h10 ;
			data[13709] <= 8'h10 ;
			data[13710] <= 8'h10 ;
			data[13711] <= 8'h10 ;
			data[13712] <= 8'h10 ;
			data[13713] <= 8'h10 ;
			data[13714] <= 8'h10 ;
			data[13715] <= 8'h10 ;
			data[13716] <= 8'h10 ;
			data[13717] <= 8'h10 ;
			data[13718] <= 8'h10 ;
			data[13719] <= 8'h10 ;
			data[13720] <= 8'h10 ;
			data[13721] <= 8'h10 ;
			data[13722] <= 8'h10 ;
			data[13723] <= 8'h10 ;
			data[13724] <= 8'h10 ;
			data[13725] <= 8'h10 ;
			data[13726] <= 8'h10 ;
			data[13727] <= 8'h10 ;
			data[13728] <= 8'h10 ;
			data[13729] <= 8'h10 ;
			data[13730] <= 8'h10 ;
			data[13731] <= 8'h10 ;
			data[13732] <= 8'h10 ;
			data[13733] <= 8'h10 ;
			data[13734] <= 8'h10 ;
			data[13735] <= 8'h10 ;
			data[13736] <= 8'h10 ;
			data[13737] <= 8'h10 ;
			data[13738] <= 8'h10 ;
			data[13739] <= 8'h10 ;
			data[13740] <= 8'h10 ;
			data[13741] <= 8'h10 ;
			data[13742] <= 8'h10 ;
			data[13743] <= 8'h10 ;
			data[13744] <= 8'h10 ;
			data[13745] <= 8'h10 ;
			data[13746] <= 8'h10 ;
			data[13747] <= 8'h10 ;
			data[13748] <= 8'h10 ;
			data[13749] <= 8'h10 ;
			data[13750] <= 8'h10 ;
			data[13751] <= 8'h10 ;
			data[13752] <= 8'h10 ;
			data[13753] <= 8'h10 ;
			data[13754] <= 8'h10 ;
			data[13755] <= 8'h10 ;
			data[13756] <= 8'h10 ;
			data[13757] <= 8'h10 ;
			data[13758] <= 8'h10 ;
			data[13759] <= 8'h10 ;
			data[13760] <= 8'h10 ;
			data[13761] <= 8'h10 ;
			data[13762] <= 8'h10 ;
			data[13763] <= 8'h10 ;
			data[13764] <= 8'h10 ;
			data[13765] <= 8'h10 ;
			data[13766] <= 8'h10 ;
			data[13767] <= 8'h10 ;
			data[13768] <= 8'h10 ;
			data[13769] <= 8'h10 ;
			data[13770] <= 8'h10 ;
			data[13771] <= 8'h10 ;
			data[13772] <= 8'h10 ;
			data[13773] <= 8'h10 ;
			data[13774] <= 8'h10 ;
			data[13775] <= 8'h10 ;
			data[13776] <= 8'h10 ;
			data[13777] <= 8'h10 ;
			data[13778] <= 8'h10 ;
			data[13779] <= 8'h10 ;
			data[13780] <= 8'h10 ;
			data[13781] <= 8'h10 ;
			data[13782] <= 8'h10 ;
			data[13783] <= 8'h10 ;
			data[13784] <= 8'h10 ;
			data[13785] <= 8'h10 ;
			data[13786] <= 8'h10 ;
			data[13787] <= 8'h10 ;
			data[13788] <= 8'h10 ;
			data[13789] <= 8'h10 ;
			data[13790] <= 8'h10 ;
			data[13791] <= 8'h10 ;
			data[13792] <= 8'h10 ;
			data[13793] <= 8'h10 ;
			data[13794] <= 8'h10 ;
			data[13795] <= 8'h10 ;
			data[13796] <= 8'h10 ;
			data[13797] <= 8'h10 ;
			data[13798] <= 8'h10 ;
			data[13799] <= 8'h10 ;
			data[13800] <= 8'h10 ;
			data[13801] <= 8'h10 ;
			data[13802] <= 8'h10 ;
			data[13803] <= 8'h10 ;
			data[13804] <= 8'h10 ;
			data[13805] <= 8'h10 ;
			data[13806] <= 8'h10 ;
			data[13807] <= 8'h10 ;
			data[13808] <= 8'h10 ;
			data[13809] <= 8'h10 ;
			data[13810] <= 8'h10 ;
			data[13811] <= 8'h10 ;
			data[13812] <= 8'h10 ;
			data[13813] <= 8'h10 ;
			data[13814] <= 8'h10 ;
			data[13815] <= 8'h10 ;
			data[13816] <= 8'h10 ;
			data[13817] <= 8'h10 ;
			data[13818] <= 8'h10 ;
			data[13819] <= 8'h10 ;
			data[13820] <= 8'h10 ;
			data[13821] <= 8'h10 ;
			data[13822] <= 8'h10 ;
			data[13823] <= 8'h10 ;
			data[13824] <= 8'h10 ;
			data[13825] <= 8'h10 ;
			data[13826] <= 8'h10 ;
			data[13827] <= 8'h10 ;
			data[13828] <= 8'h10 ;
			data[13829] <= 8'h10 ;
			data[13830] <= 8'h10 ;
			data[13831] <= 8'h10 ;
			data[13832] <= 8'h10 ;
			data[13833] <= 8'h10 ;
			data[13834] <= 8'h10 ;
			data[13835] <= 8'h10 ;
			data[13836] <= 8'h10 ;
			data[13837] <= 8'h10 ;
			data[13838] <= 8'h10 ;
			data[13839] <= 8'h10 ;
			data[13840] <= 8'h10 ;
			data[13841] <= 8'h10 ;
			data[13842] <= 8'h10 ;
			data[13843] <= 8'h10 ;
			data[13844] <= 8'h10 ;
			data[13845] <= 8'h10 ;
			data[13846] <= 8'h10 ;
			data[13847] <= 8'h10 ;
			data[13848] <= 8'h10 ;
			data[13849] <= 8'h10 ;
			data[13850] <= 8'h10 ;
			data[13851] <= 8'h10 ;
			data[13852] <= 8'h10 ;
			data[13853] <= 8'h10 ;
			data[13854] <= 8'h10 ;
			data[13855] <= 8'h10 ;
			data[13856] <= 8'h10 ;
			data[13857] <= 8'h10 ;
			data[13858] <= 8'h10 ;
			data[13859] <= 8'h10 ;
			data[13860] <= 8'h10 ;
			data[13861] <= 8'h10 ;
			data[13862] <= 8'h10 ;
			data[13863] <= 8'h10 ;
			data[13864] <= 8'h10 ;
			data[13865] <= 8'h10 ;
			data[13866] <= 8'h10 ;
			data[13867] <= 8'h10 ;
			data[13868] <= 8'h10 ;
			data[13869] <= 8'h10 ;
			data[13870] <= 8'h10 ;
			data[13871] <= 8'h10 ;
			data[13872] <= 8'h10 ;
			data[13873] <= 8'h10 ;
			data[13874] <= 8'h10 ;
			data[13875] <= 8'h10 ;
			data[13876] <= 8'h10 ;
			data[13877] <= 8'h10 ;
			data[13878] <= 8'h10 ;
			data[13879] <= 8'h10 ;
			data[13880] <= 8'h10 ;
			data[13881] <= 8'h10 ;
			data[13882] <= 8'h10 ;
			data[13883] <= 8'h10 ;
			data[13884] <= 8'h10 ;
			data[13885] <= 8'h10 ;
			data[13886] <= 8'h10 ;
			data[13887] <= 8'h10 ;
			data[13888] <= 8'h10 ;
			data[13889] <= 8'h10 ;
			data[13890] <= 8'h10 ;
			data[13891] <= 8'h10 ;
			data[13892] <= 8'h10 ;
			data[13893] <= 8'h10 ;
			data[13894] <= 8'h10 ;
			data[13895] <= 8'h10 ;
			data[13896] <= 8'h10 ;
			data[13897] <= 8'h10 ;
			data[13898] <= 8'h10 ;
			data[13899] <= 8'h10 ;
			data[13900] <= 8'h10 ;
			data[13901] <= 8'h10 ;
			data[13902] <= 8'h10 ;
			data[13903] <= 8'h10 ;
			data[13904] <= 8'h10 ;
			data[13905] <= 8'h10 ;
			data[13906] <= 8'h10 ;
			data[13907] <= 8'h10 ;
			data[13908] <= 8'h10 ;
			data[13909] <= 8'h10 ;
			data[13910] <= 8'h10 ;
			data[13911] <= 8'h10 ;
			data[13912] <= 8'h10 ;
			data[13913] <= 8'h10 ;
			data[13914] <= 8'h10 ;
			data[13915] <= 8'h10 ;
			data[13916] <= 8'h10 ;
			data[13917] <= 8'h10 ;
			data[13918] <= 8'h10 ;
			data[13919] <= 8'h10 ;
			data[13920] <= 8'h10 ;
			data[13921] <= 8'h10 ;
			data[13922] <= 8'h10 ;
			data[13923] <= 8'h10 ;
			data[13924] <= 8'h10 ;
			data[13925] <= 8'h10 ;
			data[13926] <= 8'h10 ;
			data[13927] <= 8'h10 ;
			data[13928] <= 8'h10 ;
			data[13929] <= 8'h10 ;
			data[13930] <= 8'h10 ;
			data[13931] <= 8'h10 ;
			data[13932] <= 8'h10 ;
			data[13933] <= 8'h10 ;
			data[13934] <= 8'h10 ;
			data[13935] <= 8'h10 ;
			data[13936] <= 8'h10 ;
			data[13937] <= 8'h10 ;
			data[13938] <= 8'h10 ;
			data[13939] <= 8'h10 ;
			data[13940] <= 8'h10 ;
			data[13941] <= 8'h10 ;
			data[13942] <= 8'h10 ;
			data[13943] <= 8'h10 ;
			data[13944] <= 8'h10 ;
			data[13945] <= 8'h10 ;
			data[13946] <= 8'h10 ;
			data[13947] <= 8'h10 ;
			data[13948] <= 8'h10 ;
			data[13949] <= 8'h10 ;
			data[13950] <= 8'h10 ;
			data[13951] <= 8'h10 ;
			data[13952] <= 8'h10 ;
			data[13953] <= 8'h10 ;
			data[13954] <= 8'h10 ;
			data[13955] <= 8'h10 ;
			data[13956] <= 8'h10 ;
			data[13957] <= 8'h10 ;
			data[13958] <= 8'h10 ;
			data[13959] <= 8'h10 ;
			data[13960] <= 8'h10 ;
			data[13961] <= 8'h10 ;
			data[13962] <= 8'h10 ;
			data[13963] <= 8'h10 ;
			data[13964] <= 8'h10 ;
			data[13965] <= 8'h10 ;
			data[13966] <= 8'h10 ;
			data[13967] <= 8'h10 ;
			data[13968] <= 8'h10 ;
			data[13969] <= 8'h10 ;
			data[13970] <= 8'h10 ;
			data[13971] <= 8'h10 ;
			data[13972] <= 8'h10 ;
			data[13973] <= 8'h10 ;
			data[13974] <= 8'h10 ;
			data[13975] <= 8'h10 ;
			data[13976] <= 8'h10 ;
			data[13977] <= 8'h10 ;
			data[13978] <= 8'h10 ;
			data[13979] <= 8'h10 ;
			data[13980] <= 8'h10 ;
			data[13981] <= 8'h10 ;
			data[13982] <= 8'h10 ;
			data[13983] <= 8'h10 ;
			data[13984] <= 8'h10 ;
			data[13985] <= 8'h10 ;
			data[13986] <= 8'h10 ;
			data[13987] <= 8'h10 ;
			data[13988] <= 8'h10 ;
			data[13989] <= 8'h10 ;
			data[13990] <= 8'h10 ;
			data[13991] <= 8'h10 ;
			data[13992] <= 8'h10 ;
			data[13993] <= 8'h10 ;
			data[13994] <= 8'h10 ;
			data[13995] <= 8'h10 ;
			data[13996] <= 8'h10 ;
			data[13997] <= 8'h10 ;
			data[13998] <= 8'h10 ;
			data[13999] <= 8'h10 ;
			data[14000] <= 8'h10 ;
			data[14001] <= 8'h10 ;
			data[14002] <= 8'h10 ;
			data[14003] <= 8'h10 ;
			data[14004] <= 8'h10 ;
			data[14005] <= 8'h10 ;
			data[14006] <= 8'h10 ;
			data[14007] <= 8'h10 ;
			data[14008] <= 8'h10 ;
			data[14009] <= 8'h10 ;
			data[14010] <= 8'h10 ;
			data[14011] <= 8'h10 ;
			data[14012] <= 8'h10 ;
			data[14013] <= 8'h10 ;
			data[14014] <= 8'h10 ;
			data[14015] <= 8'h10 ;
			data[14016] <= 8'h10 ;
			data[14017] <= 8'h10 ;
			data[14018] <= 8'h10 ;
			data[14019] <= 8'h10 ;
			data[14020] <= 8'h10 ;
			data[14021] <= 8'h10 ;
			data[14022] <= 8'h10 ;
			data[14023] <= 8'h10 ;
			data[14024] <= 8'h10 ;
			data[14025] <= 8'h10 ;
			data[14026] <= 8'h10 ;
			data[14027] <= 8'h10 ;
			data[14028] <= 8'h10 ;
			data[14029] <= 8'h10 ;
			data[14030] <= 8'h10 ;
			data[14031] <= 8'h10 ;
			data[14032] <= 8'h10 ;
			data[14033] <= 8'h10 ;
			data[14034] <= 8'h10 ;
			data[14035] <= 8'h10 ;
			data[14036] <= 8'h10 ;
			data[14037] <= 8'h10 ;
			data[14038] <= 8'h10 ;
			data[14039] <= 8'h10 ;
			data[14040] <= 8'h10 ;
			data[14041] <= 8'h10 ;
			data[14042] <= 8'h10 ;
			data[14043] <= 8'h10 ;
			data[14044] <= 8'h10 ;
			data[14045] <= 8'h10 ;
			data[14046] <= 8'h10 ;
			data[14047] <= 8'h10 ;
			data[14048] <= 8'h10 ;
			data[14049] <= 8'h10 ;
			data[14050] <= 8'h10 ;
			data[14051] <= 8'h10 ;
			data[14052] <= 8'h10 ;
			data[14053] <= 8'h10 ;
			data[14054] <= 8'h10 ;
			data[14055] <= 8'h10 ;
			data[14056] <= 8'h10 ;
			data[14057] <= 8'h10 ;
			data[14058] <= 8'h10 ;
			data[14059] <= 8'h10 ;
			data[14060] <= 8'h10 ;
			data[14061] <= 8'h10 ;
			data[14062] <= 8'h10 ;
			data[14063] <= 8'h10 ;
			data[14064] <= 8'h10 ;
			data[14065] <= 8'h10 ;
			data[14066] <= 8'h10 ;
			data[14067] <= 8'h10 ;
			data[14068] <= 8'h10 ;
			data[14069] <= 8'h10 ;
			data[14070] <= 8'h10 ;
			data[14071] <= 8'h10 ;
			data[14072] <= 8'h10 ;
			data[14073] <= 8'h10 ;
			data[14074] <= 8'h10 ;
			data[14075] <= 8'h10 ;
			data[14076] <= 8'h10 ;
			data[14077] <= 8'h10 ;
			data[14078] <= 8'h10 ;
			data[14079] <= 8'h10 ;
			data[14080] <= 8'h10 ;
			data[14081] <= 8'h10 ;
			data[14082] <= 8'h10 ;
			data[14083] <= 8'h10 ;
			data[14084] <= 8'h10 ;
			data[14085] <= 8'h10 ;
			data[14086] <= 8'h10 ;
			data[14087] <= 8'h10 ;
			data[14088] <= 8'h10 ;
			data[14089] <= 8'h10 ;
			data[14090] <= 8'h10 ;
			data[14091] <= 8'h10 ;
			data[14092] <= 8'h10 ;
			data[14093] <= 8'h10 ;
			data[14094] <= 8'h10 ;
			data[14095] <= 8'h10 ;
			data[14096] <= 8'h10 ;
			data[14097] <= 8'h10 ;
			data[14098] <= 8'h10 ;
			data[14099] <= 8'h10 ;
			data[14100] <= 8'h10 ;
			data[14101] <= 8'h10 ;
			data[14102] <= 8'h10 ;
			data[14103] <= 8'h10 ;
			data[14104] <= 8'h10 ;
			data[14105] <= 8'h10 ;
			data[14106] <= 8'h10 ;
			data[14107] <= 8'h10 ;
			data[14108] <= 8'h10 ;
			data[14109] <= 8'h10 ;
			data[14110] <= 8'h10 ;
			data[14111] <= 8'h10 ;
			data[14112] <= 8'h10 ;
			data[14113] <= 8'h10 ;
			data[14114] <= 8'h10 ;
			data[14115] <= 8'h10 ;
			data[14116] <= 8'h10 ;
			data[14117] <= 8'h10 ;
			data[14118] <= 8'h10 ;
			data[14119] <= 8'h10 ;
			data[14120] <= 8'h10 ;
			data[14121] <= 8'h10 ;
			data[14122] <= 8'h10 ;
			data[14123] <= 8'h10 ;
			data[14124] <= 8'h10 ;
			data[14125] <= 8'h10 ;
			data[14126] <= 8'h10 ;
			data[14127] <= 8'h10 ;
			data[14128] <= 8'h10 ;
			data[14129] <= 8'h10 ;
			data[14130] <= 8'h10 ;
			data[14131] <= 8'h10 ;
			data[14132] <= 8'h10 ;
			data[14133] <= 8'h10 ;
			data[14134] <= 8'h10 ;
			data[14135] <= 8'h10 ;
			data[14136] <= 8'h10 ;
			data[14137] <= 8'h10 ;
			data[14138] <= 8'h10 ;
			data[14139] <= 8'h10 ;
			data[14140] <= 8'h10 ;
			data[14141] <= 8'h10 ;
			data[14142] <= 8'h10 ;
			data[14143] <= 8'h10 ;
			data[14144] <= 8'h10 ;
			data[14145] <= 8'h10 ;
			data[14146] <= 8'h10 ;
			data[14147] <= 8'h10 ;
			data[14148] <= 8'h10 ;
			data[14149] <= 8'h10 ;
			data[14150] <= 8'h10 ;
			data[14151] <= 8'h10 ;
			data[14152] <= 8'h10 ;
			data[14153] <= 8'h10 ;
			data[14154] <= 8'h10 ;
			data[14155] <= 8'h10 ;
			data[14156] <= 8'h10 ;
			data[14157] <= 8'h10 ;
			data[14158] <= 8'h10 ;
			data[14159] <= 8'h10 ;
			data[14160] <= 8'h10 ;
			data[14161] <= 8'h10 ;
			data[14162] <= 8'h10 ;
			data[14163] <= 8'h10 ;
			data[14164] <= 8'h10 ;
			data[14165] <= 8'h10 ;
			data[14166] <= 8'h10 ;
			data[14167] <= 8'h10 ;
			data[14168] <= 8'h10 ;
			data[14169] <= 8'h10 ;
			data[14170] <= 8'h10 ;
			data[14171] <= 8'h10 ;
			data[14172] <= 8'h10 ;
			data[14173] <= 8'h10 ;
			data[14174] <= 8'h10 ;
			data[14175] <= 8'h10 ;
			data[14176] <= 8'h10 ;
			data[14177] <= 8'h10 ;
			data[14178] <= 8'h10 ;
			data[14179] <= 8'h10 ;
			data[14180] <= 8'h10 ;
			data[14181] <= 8'h10 ;
			data[14182] <= 8'h10 ;
			data[14183] <= 8'h10 ;
			data[14184] <= 8'h10 ;
			data[14185] <= 8'h10 ;
			data[14186] <= 8'h10 ;
			data[14187] <= 8'h10 ;
			data[14188] <= 8'h10 ;
			data[14189] <= 8'h10 ;
			data[14190] <= 8'h10 ;
			data[14191] <= 8'h10 ;
			data[14192] <= 8'h10 ;
			data[14193] <= 8'h10 ;
			data[14194] <= 8'h10 ;
			data[14195] <= 8'h10 ;
			data[14196] <= 8'h10 ;
			data[14197] <= 8'h10 ;
			data[14198] <= 8'h10 ;
			data[14199] <= 8'h10 ;
			data[14200] <= 8'h10 ;
			data[14201] <= 8'h10 ;
			data[14202] <= 8'h10 ;
			data[14203] <= 8'h10 ;
			data[14204] <= 8'h10 ;
			data[14205] <= 8'h10 ;
			data[14206] <= 8'h10 ;
			data[14207] <= 8'h10 ;
			data[14208] <= 8'h10 ;
			data[14209] <= 8'h10 ;
			data[14210] <= 8'h10 ;
			data[14211] <= 8'h10 ;
			data[14212] <= 8'h10 ;
			data[14213] <= 8'h10 ;
			data[14214] <= 8'h10 ;
			data[14215] <= 8'h10 ;
			data[14216] <= 8'h10 ;
			data[14217] <= 8'h10 ;
			data[14218] <= 8'h10 ;
			data[14219] <= 8'h10 ;
			data[14220] <= 8'h10 ;
			data[14221] <= 8'h10 ;
			data[14222] <= 8'h10 ;
			data[14223] <= 8'h10 ;
			data[14224] <= 8'h10 ;
			data[14225] <= 8'h10 ;
			data[14226] <= 8'h10 ;
			data[14227] <= 8'h10 ;
			data[14228] <= 8'h10 ;
			data[14229] <= 8'h10 ;
			data[14230] <= 8'h10 ;
			data[14231] <= 8'h10 ;
			data[14232] <= 8'h10 ;
			data[14233] <= 8'h10 ;
			data[14234] <= 8'h10 ;
			data[14235] <= 8'h10 ;
			data[14236] <= 8'h10 ;
			data[14237] <= 8'h10 ;
			data[14238] <= 8'h10 ;
			data[14239] <= 8'h10 ;
			data[14240] <= 8'h10 ;
			data[14241] <= 8'h10 ;
			data[14242] <= 8'h10 ;
			data[14243] <= 8'h10 ;
			data[14244] <= 8'h10 ;
			data[14245] <= 8'h10 ;
			data[14246] <= 8'h10 ;
			data[14247] <= 8'h10 ;
			data[14248] <= 8'h10 ;
			data[14249] <= 8'h10 ;
			data[14250] <= 8'h10 ;
			data[14251] <= 8'h10 ;
			data[14252] <= 8'h10 ;
			data[14253] <= 8'h10 ;
			data[14254] <= 8'h10 ;
			data[14255] <= 8'h10 ;
			data[14256] <= 8'h10 ;
			data[14257] <= 8'h10 ;
			data[14258] <= 8'h10 ;
			data[14259] <= 8'h10 ;
			data[14260] <= 8'h10 ;
			data[14261] <= 8'h10 ;
			data[14262] <= 8'h10 ;
			data[14263] <= 8'h10 ;
			data[14264] <= 8'h10 ;
			data[14265] <= 8'h10 ;
			data[14266] <= 8'h10 ;
			data[14267] <= 8'h10 ;
			data[14268] <= 8'h10 ;
			data[14269] <= 8'h10 ;
			data[14270] <= 8'h10 ;
			data[14271] <= 8'h10 ;
			data[14272] <= 8'h10 ;
			data[14273] <= 8'h10 ;
			data[14274] <= 8'h10 ;
			data[14275] <= 8'h10 ;
			data[14276] <= 8'h10 ;
			data[14277] <= 8'h10 ;
			data[14278] <= 8'h10 ;
			data[14279] <= 8'h10 ;
			data[14280] <= 8'h10 ;
			data[14281] <= 8'h10 ;
			data[14282] <= 8'h10 ;
			data[14283] <= 8'h10 ;
			data[14284] <= 8'h10 ;
			data[14285] <= 8'h10 ;
			data[14286] <= 8'h10 ;
			data[14287] <= 8'h10 ;
			data[14288] <= 8'h10 ;
			data[14289] <= 8'h10 ;
			data[14290] <= 8'h10 ;
			data[14291] <= 8'h10 ;
			data[14292] <= 8'h10 ;
			data[14293] <= 8'h10 ;
			data[14294] <= 8'h10 ;
			data[14295] <= 8'h10 ;
			data[14296] <= 8'h10 ;
			data[14297] <= 8'h10 ;
			data[14298] <= 8'h10 ;
			data[14299] <= 8'h10 ;
			data[14300] <= 8'h10 ;
			data[14301] <= 8'h10 ;
			data[14302] <= 8'h10 ;
			data[14303] <= 8'h10 ;
			data[14304] <= 8'h10 ;
			data[14305] <= 8'h10 ;
			data[14306] <= 8'h10 ;
			data[14307] <= 8'h10 ;
			data[14308] <= 8'h10 ;
			data[14309] <= 8'h10 ;
			data[14310] <= 8'h10 ;
			data[14311] <= 8'h10 ;
			data[14312] <= 8'h10 ;
			data[14313] <= 8'h10 ;
			data[14314] <= 8'h10 ;
			data[14315] <= 8'h10 ;
			data[14316] <= 8'h10 ;
			data[14317] <= 8'h10 ;
			data[14318] <= 8'h10 ;
			data[14319] <= 8'h10 ;
			data[14320] <= 8'h10 ;
			data[14321] <= 8'h10 ;
			data[14322] <= 8'h10 ;
			data[14323] <= 8'h10 ;
			data[14324] <= 8'h10 ;
			data[14325] <= 8'h10 ;
			data[14326] <= 8'h10 ;
			data[14327] <= 8'h10 ;
			data[14328] <= 8'h10 ;
			data[14329] <= 8'h10 ;
			data[14330] <= 8'h10 ;
			data[14331] <= 8'h10 ;
			data[14332] <= 8'h10 ;
			data[14333] <= 8'h10 ;
			data[14334] <= 8'h10 ;
			data[14335] <= 8'h10 ;
			data[14336] <= 8'h10 ;
			data[14337] <= 8'h10 ;
			data[14338] <= 8'h10 ;
			data[14339] <= 8'h10 ;
			data[14340] <= 8'h10 ;
			data[14341] <= 8'h10 ;
			data[14342] <= 8'h10 ;
			data[14343] <= 8'h10 ;
			data[14344] <= 8'h10 ;
			data[14345] <= 8'h10 ;
			data[14346] <= 8'h10 ;
			data[14347] <= 8'h10 ;
			data[14348] <= 8'h10 ;
			data[14349] <= 8'h10 ;
			data[14350] <= 8'h10 ;
			data[14351] <= 8'h10 ;
			data[14352] <= 8'h10 ;
			data[14353] <= 8'h10 ;
			data[14354] <= 8'h10 ;
			data[14355] <= 8'h10 ;
			data[14356] <= 8'h10 ;
			data[14357] <= 8'h10 ;
			data[14358] <= 8'h10 ;
			data[14359] <= 8'h10 ;
			data[14360] <= 8'h10 ;
			data[14361] <= 8'h10 ;
			data[14362] <= 8'h10 ;
			data[14363] <= 8'h10 ;
			data[14364] <= 8'h10 ;
			data[14365] <= 8'h10 ;
			data[14366] <= 8'h10 ;
			data[14367] <= 8'h10 ;
			data[14368] <= 8'h10 ;
			data[14369] <= 8'h10 ;
			data[14370] <= 8'h10 ;
			data[14371] <= 8'h10 ;
			data[14372] <= 8'h10 ;
			data[14373] <= 8'h10 ;
			data[14374] <= 8'h10 ;
			data[14375] <= 8'h10 ;
			data[14376] <= 8'h10 ;
			data[14377] <= 8'h10 ;
			data[14378] <= 8'h10 ;
			data[14379] <= 8'h10 ;
			data[14380] <= 8'h10 ;
			data[14381] <= 8'h10 ;
			data[14382] <= 8'h10 ;
			data[14383] <= 8'h10 ;
			data[14384] <= 8'h10 ;
			data[14385] <= 8'h10 ;
			data[14386] <= 8'h10 ;
			data[14387] <= 8'h10 ;
			data[14388] <= 8'h10 ;
			data[14389] <= 8'h10 ;
			data[14390] <= 8'h10 ;
			data[14391] <= 8'h10 ;
			data[14392] <= 8'h10 ;
			data[14393] <= 8'h10 ;
			data[14394] <= 8'h10 ;
			data[14395] <= 8'h10 ;
			data[14396] <= 8'h10 ;
			data[14397] <= 8'h10 ;
			data[14398] <= 8'h10 ;
			data[14399] <= 8'h10 ;
			data[14400] <= 8'h10 ;
			data[14401] <= 8'h10 ;
			data[14402] <= 8'h10 ;
			data[14403] <= 8'h10 ;
			data[14404] <= 8'h10 ;
			data[14405] <= 8'h10 ;
			data[14406] <= 8'h10 ;
			data[14407] <= 8'h10 ;
			data[14408] <= 8'h10 ;
			data[14409] <= 8'h10 ;
			data[14410] <= 8'h10 ;
			data[14411] <= 8'h10 ;
			data[14412] <= 8'h10 ;
			data[14413] <= 8'h10 ;
			data[14414] <= 8'h10 ;
			data[14415] <= 8'h10 ;
			data[14416] <= 8'h10 ;
			data[14417] <= 8'h10 ;
			data[14418] <= 8'h10 ;
			data[14419] <= 8'h10 ;
			data[14420] <= 8'h10 ;
			data[14421] <= 8'h10 ;
			data[14422] <= 8'h10 ;
			data[14423] <= 8'h10 ;
			data[14424] <= 8'h10 ;
			data[14425] <= 8'h10 ;
			data[14426] <= 8'h10 ;
			data[14427] <= 8'h10 ;
			data[14428] <= 8'h10 ;
			data[14429] <= 8'h10 ;
			data[14430] <= 8'h10 ;
			data[14431] <= 8'h10 ;
			data[14432] <= 8'h10 ;
			data[14433] <= 8'h10 ;
			data[14434] <= 8'h10 ;
			data[14435] <= 8'h10 ;
			data[14436] <= 8'h10 ;
			data[14437] <= 8'h10 ;
			data[14438] <= 8'h10 ;
			data[14439] <= 8'h10 ;
			data[14440] <= 8'h10 ;
			data[14441] <= 8'h10 ;
			data[14442] <= 8'h10 ;
			data[14443] <= 8'h10 ;
			data[14444] <= 8'h10 ;
			data[14445] <= 8'h10 ;
			data[14446] <= 8'h10 ;
			data[14447] <= 8'h10 ;
			data[14448] <= 8'h10 ;
			data[14449] <= 8'h10 ;
			data[14450] <= 8'h10 ;
			data[14451] <= 8'h10 ;
			data[14452] <= 8'h10 ;
			data[14453] <= 8'h10 ;
			data[14454] <= 8'h10 ;
			data[14455] <= 8'h10 ;
			data[14456] <= 8'h10 ;
			data[14457] <= 8'h10 ;
			data[14458] <= 8'h10 ;
			data[14459] <= 8'h10 ;
			data[14460] <= 8'h10 ;
			data[14461] <= 8'h10 ;
			data[14462] <= 8'h10 ;
			data[14463] <= 8'h10 ;
			data[14464] <= 8'h10 ;
			data[14465] <= 8'h10 ;
			data[14466] <= 8'h10 ;
			data[14467] <= 8'h10 ;
			data[14468] <= 8'h10 ;
			data[14469] <= 8'h10 ;
			data[14470] <= 8'h10 ;
			data[14471] <= 8'h10 ;
			data[14472] <= 8'h10 ;
			data[14473] <= 8'h10 ;
			data[14474] <= 8'h10 ;
			data[14475] <= 8'h10 ;
			data[14476] <= 8'h10 ;
			data[14477] <= 8'h10 ;
			data[14478] <= 8'h10 ;
			data[14479] <= 8'h10 ;
			data[14480] <= 8'h10 ;
			data[14481] <= 8'h10 ;
			data[14482] <= 8'h10 ;
			data[14483] <= 8'h10 ;
			data[14484] <= 8'h10 ;
			data[14485] <= 8'h10 ;
			data[14486] <= 8'h10 ;
			data[14487] <= 8'h10 ;
			data[14488] <= 8'h10 ;
			data[14489] <= 8'h10 ;
			data[14490] <= 8'h10 ;
			data[14491] <= 8'h10 ;
			data[14492] <= 8'h10 ;
			data[14493] <= 8'h10 ;
			data[14494] <= 8'h10 ;
			data[14495] <= 8'h10 ;
			data[14496] <= 8'h10 ;
			data[14497] <= 8'h10 ;
			data[14498] <= 8'h10 ;
			data[14499] <= 8'h10 ;
			data[14500] <= 8'h10 ;
			data[14501] <= 8'h10 ;
			data[14502] <= 8'h10 ;
			data[14503] <= 8'h10 ;
			data[14504] <= 8'h10 ;
			data[14505] <= 8'h10 ;
			data[14506] <= 8'h10 ;
			data[14507] <= 8'h10 ;
			data[14508] <= 8'h10 ;
			data[14509] <= 8'h10 ;
			data[14510] <= 8'h10 ;
			data[14511] <= 8'h10 ;
			data[14512] <= 8'h10 ;
			data[14513] <= 8'h10 ;
			data[14514] <= 8'h10 ;
			data[14515] <= 8'h10 ;
			data[14516] <= 8'h10 ;
			data[14517] <= 8'h10 ;
			data[14518] <= 8'h10 ;
			data[14519] <= 8'h10 ;
			data[14520] <= 8'h10 ;
			data[14521] <= 8'h10 ;
			data[14522] <= 8'h10 ;
			data[14523] <= 8'h10 ;
			data[14524] <= 8'h10 ;
			data[14525] <= 8'h10 ;
			data[14526] <= 8'h10 ;
			data[14527] <= 8'h10 ;
			data[14528] <= 8'h10 ;
			data[14529] <= 8'h10 ;
			data[14530] <= 8'h10 ;
			data[14531] <= 8'h10 ;
			data[14532] <= 8'h10 ;
			data[14533] <= 8'h10 ;
			data[14534] <= 8'h10 ;
			data[14535] <= 8'h10 ;
			data[14536] <= 8'h10 ;
			data[14537] <= 8'h10 ;
			data[14538] <= 8'h10 ;
			data[14539] <= 8'h10 ;
			data[14540] <= 8'h10 ;
			data[14541] <= 8'h10 ;
			data[14542] <= 8'h10 ;
			data[14543] <= 8'h10 ;
			data[14544] <= 8'h10 ;
			data[14545] <= 8'h10 ;
			data[14546] <= 8'h10 ;
			data[14547] <= 8'h10 ;
			data[14548] <= 8'h10 ;
			data[14549] <= 8'h10 ;
			data[14550] <= 8'h10 ;
			data[14551] <= 8'h10 ;
			data[14552] <= 8'h10 ;
			data[14553] <= 8'h10 ;
			data[14554] <= 8'h10 ;
			data[14555] <= 8'h10 ;
			data[14556] <= 8'h10 ;
			data[14557] <= 8'h10 ;
			data[14558] <= 8'h10 ;
			data[14559] <= 8'h10 ;
			data[14560] <= 8'h10 ;
			data[14561] <= 8'h10 ;
			data[14562] <= 8'h10 ;
			data[14563] <= 8'h10 ;
			data[14564] <= 8'h10 ;
			data[14565] <= 8'h10 ;
			data[14566] <= 8'h10 ;
			data[14567] <= 8'h10 ;
			data[14568] <= 8'h10 ;
			data[14569] <= 8'h10 ;
			data[14570] <= 8'h10 ;
			data[14571] <= 8'h10 ;
			data[14572] <= 8'h10 ;
			data[14573] <= 8'h10 ;
			data[14574] <= 8'h10 ;
			data[14575] <= 8'h10 ;
			data[14576] <= 8'h10 ;
			data[14577] <= 8'h10 ;
			data[14578] <= 8'h10 ;
			data[14579] <= 8'h10 ;
			data[14580] <= 8'h10 ;
			data[14581] <= 8'h10 ;
			data[14582] <= 8'h10 ;
			data[14583] <= 8'h10 ;
			data[14584] <= 8'h10 ;
			data[14585] <= 8'h10 ;
			data[14586] <= 8'h10 ;
			data[14587] <= 8'h10 ;
			data[14588] <= 8'h10 ;
			data[14589] <= 8'h10 ;
			data[14590] <= 8'h10 ;
			data[14591] <= 8'h10 ;
			data[14592] <= 8'h10 ;
			data[14593] <= 8'h10 ;
			data[14594] <= 8'h10 ;
			data[14595] <= 8'h10 ;
			data[14596] <= 8'h10 ;
			data[14597] <= 8'h10 ;
			data[14598] <= 8'h10 ;
			data[14599] <= 8'h10 ;
			data[14600] <= 8'h10 ;
			data[14601] <= 8'h10 ;
			data[14602] <= 8'h10 ;
			data[14603] <= 8'h10 ;
			data[14604] <= 8'h10 ;
			data[14605] <= 8'h10 ;
			data[14606] <= 8'h10 ;
			data[14607] <= 8'h10 ;
			data[14608] <= 8'h10 ;
			data[14609] <= 8'h10 ;
			data[14610] <= 8'h10 ;
			data[14611] <= 8'h10 ;
			data[14612] <= 8'h10 ;
			data[14613] <= 8'h10 ;
			data[14614] <= 8'h10 ;
			data[14615] <= 8'h10 ;
			data[14616] <= 8'h10 ;
			data[14617] <= 8'h10 ;
			data[14618] <= 8'h10 ;
			data[14619] <= 8'h10 ;
			data[14620] <= 8'h10 ;
			data[14621] <= 8'h10 ;
			data[14622] <= 8'h10 ;
			data[14623] <= 8'h10 ;
			data[14624] <= 8'h10 ;
			data[14625] <= 8'h10 ;
			data[14626] <= 8'h10 ;
			data[14627] <= 8'h10 ;
			data[14628] <= 8'h10 ;
			data[14629] <= 8'h10 ;
			data[14630] <= 8'h10 ;
			data[14631] <= 8'h10 ;
			data[14632] <= 8'h10 ;
			data[14633] <= 8'h10 ;
			data[14634] <= 8'h10 ;
			data[14635] <= 8'h10 ;
			data[14636] <= 8'h10 ;
			data[14637] <= 8'h10 ;
			data[14638] <= 8'h10 ;
			data[14639] <= 8'h10 ;
			data[14640] <= 8'h10 ;
			data[14641] <= 8'h10 ;
			data[14642] <= 8'h10 ;
			data[14643] <= 8'h10 ;
			data[14644] <= 8'h10 ;
			data[14645] <= 8'h10 ;
			data[14646] <= 8'h10 ;
			data[14647] <= 8'h10 ;
			data[14648] <= 8'h10 ;
			data[14649] <= 8'h10 ;
			data[14650] <= 8'h10 ;
			data[14651] <= 8'h10 ;
			data[14652] <= 8'h10 ;
			data[14653] <= 8'h10 ;
			data[14654] <= 8'h10 ;
			data[14655] <= 8'h10 ;
			data[14656] <= 8'h10 ;
			data[14657] <= 8'h10 ;
			data[14658] <= 8'h10 ;
			data[14659] <= 8'h10 ;
			data[14660] <= 8'h10 ;
			data[14661] <= 8'h10 ;
			data[14662] <= 8'h10 ;
			data[14663] <= 8'h10 ;
			data[14664] <= 8'h10 ;
			data[14665] <= 8'h10 ;
			data[14666] <= 8'h10 ;
			data[14667] <= 8'h10 ;
			data[14668] <= 8'h10 ;
			data[14669] <= 8'h10 ;
			data[14670] <= 8'h10 ;
			data[14671] <= 8'h10 ;
			data[14672] <= 8'h10 ;
			data[14673] <= 8'h10 ;
			data[14674] <= 8'h10 ;
			data[14675] <= 8'h10 ;
			data[14676] <= 8'h10 ;
			data[14677] <= 8'h10 ;
			data[14678] <= 8'h10 ;
			data[14679] <= 8'h10 ;
			data[14680] <= 8'h10 ;
			data[14681] <= 8'h10 ;
			data[14682] <= 8'h10 ;
			data[14683] <= 8'h10 ;
			data[14684] <= 8'h10 ;
			data[14685] <= 8'h10 ;
			data[14686] <= 8'h10 ;
			data[14687] <= 8'h10 ;
			data[14688] <= 8'h10 ;
			data[14689] <= 8'h10 ;
			data[14690] <= 8'h10 ;
			data[14691] <= 8'h10 ;
			data[14692] <= 8'h10 ;
			data[14693] <= 8'h10 ;
			data[14694] <= 8'h10 ;
			data[14695] <= 8'h10 ;
			data[14696] <= 8'h10 ;
			data[14697] <= 8'h10 ;
			data[14698] <= 8'h10 ;
			data[14699] <= 8'h10 ;
			data[14700] <= 8'h10 ;
			data[14701] <= 8'h10 ;
			data[14702] <= 8'h10 ;
			data[14703] <= 8'h10 ;
			data[14704] <= 8'h10 ;
			data[14705] <= 8'h10 ;
			data[14706] <= 8'h10 ;
			data[14707] <= 8'h10 ;
			data[14708] <= 8'h10 ;
			data[14709] <= 8'h10 ;
			data[14710] <= 8'h10 ;
			data[14711] <= 8'h10 ;
			data[14712] <= 8'h10 ;
			data[14713] <= 8'h10 ;
			data[14714] <= 8'h10 ;
			data[14715] <= 8'h10 ;
			data[14716] <= 8'h10 ;
			data[14717] <= 8'h10 ;
			data[14718] <= 8'h10 ;
			data[14719] <= 8'h10 ;
			data[14720] <= 8'h10 ;
			data[14721] <= 8'h10 ;
			data[14722] <= 8'h10 ;
			data[14723] <= 8'h10 ;
			data[14724] <= 8'h10 ;
			data[14725] <= 8'h10 ;
			data[14726] <= 8'h10 ;
			data[14727] <= 8'h10 ;
			data[14728] <= 8'h10 ;
			data[14729] <= 8'h10 ;
			data[14730] <= 8'h10 ;
			data[14731] <= 8'h10 ;
			data[14732] <= 8'h10 ;
			data[14733] <= 8'h10 ;
			data[14734] <= 8'h10 ;
			data[14735] <= 8'h10 ;
			data[14736] <= 8'h10 ;
			data[14737] <= 8'h10 ;
			data[14738] <= 8'h10 ;
			data[14739] <= 8'h10 ;
			data[14740] <= 8'h10 ;
			data[14741] <= 8'h10 ;
			data[14742] <= 8'h10 ;
			data[14743] <= 8'h10 ;
			data[14744] <= 8'h10 ;
			data[14745] <= 8'h10 ;
			data[14746] <= 8'h10 ;
			data[14747] <= 8'h10 ;
			data[14748] <= 8'h10 ;
			data[14749] <= 8'h10 ;
			data[14750] <= 8'h10 ;
			data[14751] <= 8'h10 ;
			data[14752] <= 8'h10 ;
			data[14753] <= 8'h10 ;
			data[14754] <= 8'h10 ;
			data[14755] <= 8'h10 ;
			data[14756] <= 8'h10 ;
			data[14757] <= 8'h10 ;
			data[14758] <= 8'h10 ;
			data[14759] <= 8'h10 ;
			data[14760] <= 8'h10 ;
			data[14761] <= 8'h10 ;
			data[14762] <= 8'h10 ;
			data[14763] <= 8'h10 ;
			data[14764] <= 8'h10 ;
			data[14765] <= 8'h10 ;
			data[14766] <= 8'h10 ;
			data[14767] <= 8'h10 ;
			data[14768] <= 8'h10 ;
			data[14769] <= 8'h10 ;
			data[14770] <= 8'h10 ;
			data[14771] <= 8'h10 ;
			data[14772] <= 8'h10 ;
			data[14773] <= 8'h10 ;
			data[14774] <= 8'h10 ;
			data[14775] <= 8'h10 ;
			data[14776] <= 8'h10 ;
			data[14777] <= 8'h10 ;
			data[14778] <= 8'h10 ;
			data[14779] <= 8'h10 ;
			data[14780] <= 8'h10 ;
			data[14781] <= 8'h10 ;
			data[14782] <= 8'h10 ;
			data[14783] <= 8'h10 ;
			data[14784] <= 8'h10 ;
			data[14785] <= 8'h10 ;
			data[14786] <= 8'h10 ;
			data[14787] <= 8'h10 ;
			data[14788] <= 8'h10 ;
			data[14789] <= 8'h10 ;
			data[14790] <= 8'h10 ;
			data[14791] <= 8'h10 ;
			data[14792] <= 8'h10 ;
			data[14793] <= 8'h10 ;
			data[14794] <= 8'h10 ;
			data[14795] <= 8'h10 ;
			data[14796] <= 8'h10 ;
			data[14797] <= 8'h10 ;
			data[14798] <= 8'h10 ;
			data[14799] <= 8'h10 ;
			data[14800] <= 8'h10 ;
			data[14801] <= 8'h10 ;
			data[14802] <= 8'h10 ;
			data[14803] <= 8'h10 ;
			data[14804] <= 8'h10 ;
			data[14805] <= 8'h10 ;
			data[14806] <= 8'h10 ;
			data[14807] <= 8'h10 ;
			data[14808] <= 8'h10 ;
			data[14809] <= 8'h10 ;
			data[14810] <= 8'h10 ;
			data[14811] <= 8'h10 ;
			data[14812] <= 8'h10 ;
			data[14813] <= 8'h10 ;
			data[14814] <= 8'h10 ;
			data[14815] <= 8'h10 ;
			data[14816] <= 8'h10 ;
			data[14817] <= 8'h10 ;
			data[14818] <= 8'h10 ;
			data[14819] <= 8'h10 ;
			data[14820] <= 8'h10 ;
			data[14821] <= 8'h10 ;
			data[14822] <= 8'h10 ;
			data[14823] <= 8'h10 ;
			data[14824] <= 8'h10 ;
			data[14825] <= 8'h10 ;
			data[14826] <= 8'h10 ;
			data[14827] <= 8'h10 ;
			data[14828] <= 8'h10 ;
			data[14829] <= 8'h10 ;
			data[14830] <= 8'h10 ;
			data[14831] <= 8'h10 ;
			data[14832] <= 8'h10 ;
			data[14833] <= 8'h10 ;
			data[14834] <= 8'h10 ;
			data[14835] <= 8'h10 ;
			data[14836] <= 8'h10 ;
			data[14837] <= 8'h10 ;
			data[14838] <= 8'h10 ;
			data[14839] <= 8'h10 ;
			data[14840] <= 8'h10 ;
			data[14841] <= 8'h10 ;
			data[14842] <= 8'h10 ;
			data[14843] <= 8'h10 ;
			data[14844] <= 8'h10 ;
			data[14845] <= 8'h10 ;
			data[14846] <= 8'h10 ;
			data[14847] <= 8'h10 ;
			data[14848] <= 8'h10 ;
			data[14849] <= 8'h10 ;
			data[14850] <= 8'h10 ;
			data[14851] <= 8'h10 ;
			data[14852] <= 8'h10 ;
			data[14853] <= 8'h10 ;
			data[14854] <= 8'h10 ;
			data[14855] <= 8'h10 ;
			data[14856] <= 8'h10 ;
			data[14857] <= 8'h10 ;
			data[14858] <= 8'h10 ;
			data[14859] <= 8'h10 ;
			data[14860] <= 8'h10 ;
			data[14861] <= 8'h10 ;
			data[14862] <= 8'h10 ;
			data[14863] <= 8'h10 ;
			data[14864] <= 8'h10 ;
			data[14865] <= 8'h10 ;
			data[14866] <= 8'h10 ;
			data[14867] <= 8'h10 ;
			data[14868] <= 8'h10 ;
			data[14869] <= 8'h10 ;
			data[14870] <= 8'h10 ;
			data[14871] <= 8'h10 ;
			data[14872] <= 8'h10 ;
			data[14873] <= 8'h10 ;
			data[14874] <= 8'h10 ;
			data[14875] <= 8'h10 ;
			data[14876] <= 8'h10 ;
			data[14877] <= 8'h10 ;
			data[14878] <= 8'h10 ;
			data[14879] <= 8'h10 ;
			data[14880] <= 8'h10 ;
			data[14881] <= 8'h10 ;
			data[14882] <= 8'h10 ;
			data[14883] <= 8'h10 ;
			data[14884] <= 8'h10 ;
			data[14885] <= 8'h10 ;
			data[14886] <= 8'h10 ;
			data[14887] <= 8'h10 ;
			data[14888] <= 8'h10 ;
			data[14889] <= 8'h10 ;
			data[14890] <= 8'h10 ;
			data[14891] <= 8'h10 ;
			data[14892] <= 8'h10 ;
			data[14893] <= 8'h10 ;
			data[14894] <= 8'h10 ;
			data[14895] <= 8'h10 ;
			data[14896] <= 8'h10 ;
			data[14897] <= 8'h10 ;
			data[14898] <= 8'h10 ;
			data[14899] <= 8'h10 ;
			data[14900] <= 8'h10 ;
			data[14901] <= 8'h10 ;
			data[14902] <= 8'h10 ;
			data[14903] <= 8'h10 ;
			data[14904] <= 8'h10 ;
			data[14905] <= 8'h10 ;
			data[14906] <= 8'h10 ;
			data[14907] <= 8'h10 ;
			data[14908] <= 8'h10 ;
			data[14909] <= 8'h10 ;
			data[14910] <= 8'h10 ;
			data[14911] <= 8'h10 ;
			data[14912] <= 8'h10 ;
			data[14913] <= 8'h10 ;
			data[14914] <= 8'h10 ;
			data[14915] <= 8'h10 ;
			data[14916] <= 8'h10 ;
			data[14917] <= 8'h10 ;
			data[14918] <= 8'h10 ;
			data[14919] <= 8'h10 ;
			data[14920] <= 8'h10 ;
			data[14921] <= 8'h10 ;
			data[14922] <= 8'h10 ;
			data[14923] <= 8'h10 ;
			data[14924] <= 8'h10 ;
			data[14925] <= 8'h10 ;
			data[14926] <= 8'h10 ;
			data[14927] <= 8'h10 ;
			data[14928] <= 8'h10 ;
			data[14929] <= 8'h10 ;
			data[14930] <= 8'h10 ;
			data[14931] <= 8'h10 ;
			data[14932] <= 8'h10 ;
			data[14933] <= 8'h10 ;
			data[14934] <= 8'h10 ;
			data[14935] <= 8'h10 ;
			data[14936] <= 8'h10 ;
			data[14937] <= 8'h10 ;
			data[14938] <= 8'h10 ;
			data[14939] <= 8'h10 ;
			data[14940] <= 8'h10 ;
			data[14941] <= 8'h10 ;
			data[14942] <= 8'h10 ;
			data[14943] <= 8'h10 ;
			data[14944] <= 8'h10 ;
			data[14945] <= 8'h10 ;
			data[14946] <= 8'h10 ;
			data[14947] <= 8'h10 ;
			data[14948] <= 8'h10 ;
			data[14949] <= 8'h10 ;
			data[14950] <= 8'h10 ;
			data[14951] <= 8'h10 ;
			data[14952] <= 8'h10 ;
			data[14953] <= 8'h10 ;
			data[14954] <= 8'h10 ;
			data[14955] <= 8'h10 ;
			data[14956] <= 8'h10 ;
			data[14957] <= 8'h10 ;
			data[14958] <= 8'h10 ;
			data[14959] <= 8'h10 ;
			data[14960] <= 8'h10 ;
			data[14961] <= 8'h10 ;
			data[14962] <= 8'h10 ;
			data[14963] <= 8'h10 ;
			data[14964] <= 8'h10 ;
			data[14965] <= 8'h10 ;
			data[14966] <= 8'h10 ;
			data[14967] <= 8'h10 ;
			data[14968] <= 8'h10 ;
			data[14969] <= 8'h10 ;
			data[14970] <= 8'h10 ;
			data[14971] <= 8'h10 ;
			data[14972] <= 8'h10 ;
			data[14973] <= 8'h10 ;
			data[14974] <= 8'h10 ;
			data[14975] <= 8'h10 ;
			data[14976] <= 8'h10 ;
			data[14977] <= 8'h10 ;
			data[14978] <= 8'h10 ;
			data[14979] <= 8'h10 ;
			data[14980] <= 8'h10 ;
			data[14981] <= 8'h10 ;
			data[14982] <= 8'h10 ;
			data[14983] <= 8'h10 ;
			data[14984] <= 8'h10 ;
			data[14985] <= 8'h10 ;
			data[14986] <= 8'h10 ;
			data[14987] <= 8'h10 ;
			data[14988] <= 8'h10 ;
			data[14989] <= 8'h10 ;
			data[14990] <= 8'h10 ;
			data[14991] <= 8'h10 ;
			data[14992] <= 8'h10 ;
			data[14993] <= 8'h10 ;
			data[14994] <= 8'h10 ;
			data[14995] <= 8'h10 ;
			data[14996] <= 8'h10 ;
			data[14997] <= 8'h10 ;
			data[14998] <= 8'h10 ;
			data[14999] <= 8'h10 ;
			data[15000] <= 8'h10 ;
			data[15001] <= 8'h10 ;
			data[15002] <= 8'h10 ;
			data[15003] <= 8'h10 ;
			data[15004] <= 8'h10 ;
			data[15005] <= 8'h10 ;
			data[15006] <= 8'h10 ;
			data[15007] <= 8'h10 ;
			data[15008] <= 8'h10 ;
			data[15009] <= 8'h10 ;
			data[15010] <= 8'h10 ;
			data[15011] <= 8'h10 ;
			data[15012] <= 8'h10 ;
			data[15013] <= 8'h10 ;
			data[15014] <= 8'h10 ;
			data[15015] <= 8'h10 ;
			data[15016] <= 8'h10 ;
			data[15017] <= 8'h10 ;
			data[15018] <= 8'h10 ;
			data[15019] <= 8'h10 ;
			data[15020] <= 8'h10 ;
			data[15021] <= 8'h10 ;
			data[15022] <= 8'h10 ;
			data[15023] <= 8'h10 ;
			data[15024] <= 8'h10 ;
			data[15025] <= 8'h10 ;
			data[15026] <= 8'h10 ;
			data[15027] <= 8'h10 ;
			data[15028] <= 8'h10 ;
			data[15029] <= 8'h10 ;
			data[15030] <= 8'h10 ;
			data[15031] <= 8'h10 ;
			data[15032] <= 8'h10 ;
			data[15033] <= 8'h10 ;
			data[15034] <= 8'h10 ;
			data[15035] <= 8'h10 ;
			data[15036] <= 8'h10 ;
			data[15037] <= 8'h10 ;
			data[15038] <= 8'h10 ;
			data[15039] <= 8'h10 ;
			data[15040] <= 8'h10 ;
			data[15041] <= 8'h10 ;
			data[15042] <= 8'h10 ;
			data[15043] <= 8'h10 ;
			data[15044] <= 8'h10 ;
			data[15045] <= 8'h10 ;
			data[15046] <= 8'h10 ;
			data[15047] <= 8'h10 ;
			data[15048] <= 8'h10 ;
			data[15049] <= 8'h10 ;
			data[15050] <= 8'h10 ;
			data[15051] <= 8'h10 ;
			data[15052] <= 8'h10 ;
			data[15053] <= 8'h10 ;
			data[15054] <= 8'h10 ;
			data[15055] <= 8'h10 ;
			data[15056] <= 8'h10 ;
			data[15057] <= 8'h10 ;
			data[15058] <= 8'h10 ;
			data[15059] <= 8'h10 ;
			data[15060] <= 8'h10 ;
			data[15061] <= 8'h10 ;
			data[15062] <= 8'h10 ;
			data[15063] <= 8'h10 ;
			data[15064] <= 8'h10 ;
			data[15065] <= 8'h10 ;
			data[15066] <= 8'h10 ;
			data[15067] <= 8'h10 ;
			data[15068] <= 8'h10 ;
			data[15069] <= 8'h10 ;
			data[15070] <= 8'h10 ;
			data[15071] <= 8'h10 ;
			data[15072] <= 8'h10 ;
			data[15073] <= 8'h10 ;
			data[15074] <= 8'h10 ;
			data[15075] <= 8'h10 ;
			data[15076] <= 8'h10 ;
			data[15077] <= 8'h10 ;
			data[15078] <= 8'h10 ;
			data[15079] <= 8'h10 ;
			data[15080] <= 8'h10 ;
			data[15081] <= 8'h10 ;
			data[15082] <= 8'h10 ;
			data[15083] <= 8'h10 ;
			data[15084] <= 8'h10 ;
			data[15085] <= 8'h10 ;
			data[15086] <= 8'h10 ;
			data[15087] <= 8'h10 ;
			data[15088] <= 8'h10 ;
			data[15089] <= 8'h10 ;
			data[15090] <= 8'h10 ;
			data[15091] <= 8'h10 ;
			data[15092] <= 8'h10 ;
			data[15093] <= 8'h10 ;
			data[15094] <= 8'h10 ;
			data[15095] <= 8'h10 ;
			data[15096] <= 8'h10 ;
			data[15097] <= 8'h10 ;
			data[15098] <= 8'h10 ;
			data[15099] <= 8'h10 ;
			data[15100] <= 8'h10 ;
			data[15101] <= 8'h10 ;
			data[15102] <= 8'h10 ;
			data[15103] <= 8'h10 ;
			data[15104] <= 8'h10 ;
			data[15105] <= 8'h10 ;
			data[15106] <= 8'h10 ;
			data[15107] <= 8'h10 ;
			data[15108] <= 8'h10 ;
			data[15109] <= 8'h10 ;
			data[15110] <= 8'h10 ;
			data[15111] <= 8'h10 ;
			data[15112] <= 8'h10 ;
			data[15113] <= 8'h10 ;
			data[15114] <= 8'h10 ;
			data[15115] <= 8'h10 ;
			data[15116] <= 8'h10 ;
			data[15117] <= 8'h10 ;
			data[15118] <= 8'h10 ;
			data[15119] <= 8'h10 ;
			data[15120] <= 8'h10 ;
			data[15121] <= 8'h10 ;
			data[15122] <= 8'h10 ;
			data[15123] <= 8'h10 ;
			data[15124] <= 8'h10 ;
			data[15125] <= 8'h10 ;
			data[15126] <= 8'h10 ;
			data[15127] <= 8'h10 ;
			data[15128] <= 8'h10 ;
			data[15129] <= 8'h10 ;
			data[15130] <= 8'h10 ;
			data[15131] <= 8'h10 ;
			data[15132] <= 8'h10 ;
			data[15133] <= 8'h10 ;
			data[15134] <= 8'h10 ;
			data[15135] <= 8'h10 ;
			data[15136] <= 8'h10 ;
			data[15137] <= 8'h10 ;
			data[15138] <= 8'h10 ;
			data[15139] <= 8'h10 ;
			data[15140] <= 8'h10 ;
			data[15141] <= 8'h10 ;
			data[15142] <= 8'h10 ;
			data[15143] <= 8'h10 ;
			data[15144] <= 8'h10 ;
			data[15145] <= 8'h10 ;
			data[15146] <= 8'h10 ;
			data[15147] <= 8'h10 ;
			data[15148] <= 8'h10 ;
			data[15149] <= 8'h10 ;
			data[15150] <= 8'h10 ;
			data[15151] <= 8'h10 ;
			data[15152] <= 8'h10 ;
			data[15153] <= 8'h10 ;
			data[15154] <= 8'h10 ;
			data[15155] <= 8'h10 ;
			data[15156] <= 8'h10 ;
			data[15157] <= 8'h10 ;
			data[15158] <= 8'h10 ;
			data[15159] <= 8'h10 ;
			data[15160] <= 8'h10 ;
			data[15161] <= 8'h10 ;
			data[15162] <= 8'h10 ;
			data[15163] <= 8'h10 ;
			data[15164] <= 8'h10 ;
			data[15165] <= 8'h10 ;
			data[15166] <= 8'h10 ;
			data[15167] <= 8'h10 ;
			data[15168] <= 8'h10 ;
			data[15169] <= 8'h10 ;
			data[15170] <= 8'h10 ;
			data[15171] <= 8'h10 ;
			data[15172] <= 8'h10 ;
			data[15173] <= 8'h10 ;
			data[15174] <= 8'h10 ;
			data[15175] <= 8'h10 ;
			data[15176] <= 8'h10 ;
			data[15177] <= 8'h10 ;
			data[15178] <= 8'h10 ;
			data[15179] <= 8'h10 ;
			data[15180] <= 8'h10 ;
			data[15181] <= 8'h10 ;
			data[15182] <= 8'h10 ;
			data[15183] <= 8'h10 ;
			data[15184] <= 8'h10 ;
			data[15185] <= 8'h10 ;
			data[15186] <= 8'h10 ;
			data[15187] <= 8'h10 ;
			data[15188] <= 8'h10 ;
			data[15189] <= 8'h10 ;
			data[15190] <= 8'h10 ;
			data[15191] <= 8'h10 ;
			data[15192] <= 8'h10 ;
			data[15193] <= 8'h10 ;
			data[15194] <= 8'h10 ;
			data[15195] <= 8'h10 ;
			data[15196] <= 8'h10 ;
			data[15197] <= 8'h10 ;
			data[15198] <= 8'h10 ;
			data[15199] <= 8'h10 ;
			data[15200] <= 8'h10 ;
			data[15201] <= 8'h10 ;
			data[15202] <= 8'h10 ;
			data[15203] <= 8'h10 ;
			data[15204] <= 8'h10 ;
			data[15205] <= 8'h10 ;
			data[15206] <= 8'h10 ;
			data[15207] <= 8'h10 ;
			data[15208] <= 8'h10 ;
			data[15209] <= 8'h10 ;
			data[15210] <= 8'h10 ;
			data[15211] <= 8'h10 ;
			data[15212] <= 8'h10 ;
			data[15213] <= 8'h10 ;
			data[15214] <= 8'h10 ;
			data[15215] <= 8'h10 ;
			data[15216] <= 8'h10 ;
			data[15217] <= 8'h10 ;
			data[15218] <= 8'h10 ;
			data[15219] <= 8'h10 ;
			data[15220] <= 8'h10 ;
			data[15221] <= 8'h10 ;
			data[15222] <= 8'h10 ;
			data[15223] <= 8'h10 ;
			data[15224] <= 8'h10 ;
			data[15225] <= 8'h10 ;
			data[15226] <= 8'h10 ;
			data[15227] <= 8'h10 ;
			data[15228] <= 8'h10 ;
			data[15229] <= 8'h10 ;
			data[15230] <= 8'h10 ;
			data[15231] <= 8'h10 ;
			data[15232] <= 8'h10 ;
			data[15233] <= 8'h10 ;
			data[15234] <= 8'h10 ;
			data[15235] <= 8'h10 ;
			data[15236] <= 8'h10 ;
			data[15237] <= 8'h10 ;
			data[15238] <= 8'h10 ;
			data[15239] <= 8'h10 ;
			data[15240] <= 8'h10 ;
			data[15241] <= 8'h10 ;
			data[15242] <= 8'h10 ;
			data[15243] <= 8'h10 ;
			data[15244] <= 8'h10 ;
			data[15245] <= 8'h10 ;
			data[15246] <= 8'h10 ;
			data[15247] <= 8'h10 ;
			data[15248] <= 8'h10 ;
			data[15249] <= 8'h10 ;
			data[15250] <= 8'h10 ;
			data[15251] <= 8'h10 ;
			data[15252] <= 8'h10 ;
			data[15253] <= 8'h10 ;
			data[15254] <= 8'h10 ;
			data[15255] <= 8'h10 ;
			data[15256] <= 8'h10 ;
			data[15257] <= 8'h10 ;
			data[15258] <= 8'h10 ;
			data[15259] <= 8'h10 ;
			data[15260] <= 8'h10 ;
			data[15261] <= 8'h10 ;
			data[15262] <= 8'h10 ;
			data[15263] <= 8'h10 ;
			data[15264] <= 8'h10 ;
			data[15265] <= 8'h10 ;
			data[15266] <= 8'h10 ;
			data[15267] <= 8'h10 ;
			data[15268] <= 8'h10 ;
			data[15269] <= 8'h10 ;
			data[15270] <= 8'h10 ;
			data[15271] <= 8'h10 ;
			data[15272] <= 8'h10 ;
			data[15273] <= 8'h10 ;
			data[15274] <= 8'h10 ;
			data[15275] <= 8'h10 ;
			data[15276] <= 8'h10 ;
			data[15277] <= 8'h10 ;
			data[15278] <= 8'h10 ;
			data[15279] <= 8'h10 ;
			data[15280] <= 8'h10 ;
			data[15281] <= 8'h10 ;
			data[15282] <= 8'h10 ;
			data[15283] <= 8'h10 ;
			data[15284] <= 8'h10 ;
			data[15285] <= 8'h10 ;
			data[15286] <= 8'h10 ;
			data[15287] <= 8'h10 ;
			data[15288] <= 8'h10 ;
			data[15289] <= 8'h10 ;
			data[15290] <= 8'h10 ;
			data[15291] <= 8'h10 ;
			data[15292] <= 8'h10 ;
			data[15293] <= 8'h10 ;
			data[15294] <= 8'h10 ;
			data[15295] <= 8'h10 ;
			data[15296] <= 8'h10 ;
			data[15297] <= 8'h10 ;
			data[15298] <= 8'h10 ;
			data[15299] <= 8'h10 ;
			data[15300] <= 8'h10 ;
			data[15301] <= 8'h10 ;
			data[15302] <= 8'h10 ;
			data[15303] <= 8'h10 ;
			data[15304] <= 8'h10 ;
			data[15305] <= 8'h10 ;
			data[15306] <= 8'h10 ;
			data[15307] <= 8'h10 ;
			data[15308] <= 8'h10 ;
			data[15309] <= 8'h10 ;
			data[15310] <= 8'h10 ;
			data[15311] <= 8'h10 ;
			data[15312] <= 8'h10 ;
			data[15313] <= 8'h10 ;
			data[15314] <= 8'h10 ;
			data[15315] <= 8'h10 ;
			data[15316] <= 8'h10 ;
			data[15317] <= 8'h10 ;
			data[15318] <= 8'h10 ;
			data[15319] <= 8'h10 ;
			data[15320] <= 8'h10 ;
			data[15321] <= 8'h10 ;
			data[15322] <= 8'h10 ;
			data[15323] <= 8'h10 ;
			data[15324] <= 8'h10 ;
			data[15325] <= 8'h10 ;
			data[15326] <= 8'h10 ;
			data[15327] <= 8'h10 ;
			data[15328] <= 8'h10 ;
			data[15329] <= 8'h10 ;
			data[15330] <= 8'h10 ;
			data[15331] <= 8'h10 ;
			data[15332] <= 8'h10 ;
			data[15333] <= 8'h10 ;
			data[15334] <= 8'h10 ;
			data[15335] <= 8'h10 ;
			data[15336] <= 8'h10 ;
			data[15337] <= 8'h10 ;
			data[15338] <= 8'h10 ;
			data[15339] <= 8'h10 ;
			data[15340] <= 8'h10 ;
			data[15341] <= 8'h10 ;
			data[15342] <= 8'h10 ;
			data[15343] <= 8'h10 ;
			data[15344] <= 8'h10 ;
			data[15345] <= 8'h10 ;
			data[15346] <= 8'h10 ;
			data[15347] <= 8'h10 ;
			data[15348] <= 8'h10 ;
			data[15349] <= 8'h10 ;
			data[15350] <= 8'h10 ;
			data[15351] <= 8'h10 ;
			data[15352] <= 8'h10 ;
			data[15353] <= 8'h10 ;
			data[15354] <= 8'h10 ;
			data[15355] <= 8'h10 ;
			data[15356] <= 8'h10 ;
			data[15357] <= 8'h10 ;
			data[15358] <= 8'h10 ;
			data[15359] <= 8'h10 ;
			data[15360] <= 8'h10 ;
			data[15361] <= 8'h10 ;
			data[15362] <= 8'h10 ;
			data[15363] <= 8'h10 ;
			data[15364] <= 8'h10 ;
			data[15365] <= 8'h10 ;
			data[15366] <= 8'h10 ;
			data[15367] <= 8'h10 ;
			data[15368] <= 8'h10 ;
			data[15369] <= 8'h10 ;
			data[15370] <= 8'h10 ;
			data[15371] <= 8'h10 ;
			data[15372] <= 8'h10 ;
			data[15373] <= 8'h10 ;
			data[15374] <= 8'h10 ;
			data[15375] <= 8'h10 ;
			data[15376] <= 8'h10 ;
			data[15377] <= 8'h10 ;
			data[15378] <= 8'h10 ;
			data[15379] <= 8'h10 ;
			data[15380] <= 8'h10 ;
			data[15381] <= 8'h10 ;
			data[15382] <= 8'h10 ;
			data[15383] <= 8'h10 ;
			data[15384] <= 8'h10 ;
			data[15385] <= 8'h10 ;
			data[15386] <= 8'h10 ;
			data[15387] <= 8'h10 ;
			data[15388] <= 8'h10 ;
			data[15389] <= 8'h10 ;
			data[15390] <= 8'h10 ;
			data[15391] <= 8'h10 ;
			data[15392] <= 8'h10 ;
			data[15393] <= 8'h10 ;
			data[15394] <= 8'h10 ;
			data[15395] <= 8'h10 ;
			data[15396] <= 8'h10 ;
			data[15397] <= 8'h10 ;
			data[15398] <= 8'h10 ;
			data[15399] <= 8'h10 ;
			data[15400] <= 8'h10 ;
			data[15401] <= 8'h10 ;
			data[15402] <= 8'h10 ;
			data[15403] <= 8'h10 ;
			data[15404] <= 8'h10 ;
			data[15405] <= 8'h10 ;
			data[15406] <= 8'h10 ;
			data[15407] <= 8'h10 ;
			data[15408] <= 8'h10 ;
			data[15409] <= 8'h10 ;
			data[15410] <= 8'h10 ;
			data[15411] <= 8'h10 ;
			data[15412] <= 8'h10 ;
			data[15413] <= 8'h10 ;
			data[15414] <= 8'h10 ;
			data[15415] <= 8'h10 ;
			data[15416] <= 8'h10 ;
			data[15417] <= 8'h10 ;
			data[15418] <= 8'h10 ;
			data[15419] <= 8'h10 ;
			data[15420] <= 8'h10 ;
			data[15421] <= 8'h10 ;
			data[15422] <= 8'h10 ;
			data[15423] <= 8'h10 ;
			data[15424] <= 8'h10 ;
			data[15425] <= 8'h10 ;
			data[15426] <= 8'h10 ;
			data[15427] <= 8'h10 ;
			data[15428] <= 8'h10 ;
			data[15429] <= 8'h10 ;
			data[15430] <= 8'h10 ;
			data[15431] <= 8'h10 ;
			data[15432] <= 8'h10 ;
			data[15433] <= 8'h10 ;
			data[15434] <= 8'h10 ;
			data[15435] <= 8'h10 ;
			data[15436] <= 8'h10 ;
			data[15437] <= 8'h10 ;
			data[15438] <= 8'h10 ;
			data[15439] <= 8'h10 ;
			data[15440] <= 8'h10 ;
			data[15441] <= 8'h10 ;
			data[15442] <= 8'h10 ;
			data[15443] <= 8'h10 ;
			data[15444] <= 8'h10 ;
			data[15445] <= 8'h10 ;
			data[15446] <= 8'h10 ;
			data[15447] <= 8'h10 ;
			data[15448] <= 8'h10 ;
			data[15449] <= 8'h10 ;
			data[15450] <= 8'h10 ;
			data[15451] <= 8'h10 ;
			data[15452] <= 8'h10 ;
			data[15453] <= 8'h10 ;
			data[15454] <= 8'h10 ;
			data[15455] <= 8'h10 ;
			data[15456] <= 8'h10 ;
			data[15457] <= 8'h10 ;
			data[15458] <= 8'h10 ;
			data[15459] <= 8'h10 ;
			data[15460] <= 8'h10 ;
			data[15461] <= 8'h10 ;
			data[15462] <= 8'h10 ;
			data[15463] <= 8'h10 ;
			data[15464] <= 8'h10 ;
			data[15465] <= 8'h10 ;
			data[15466] <= 8'h10 ;
			data[15467] <= 8'h10 ;
			data[15468] <= 8'h10 ;
			data[15469] <= 8'h10 ;
			data[15470] <= 8'h10 ;
			data[15471] <= 8'h10 ;
			data[15472] <= 8'h10 ;
			data[15473] <= 8'h10 ;
			data[15474] <= 8'h10 ;
			data[15475] <= 8'h10 ;
			data[15476] <= 8'h10 ;
			data[15477] <= 8'h10 ;
			data[15478] <= 8'h10 ;
			data[15479] <= 8'h10 ;
			data[15480] <= 8'h10 ;
			data[15481] <= 8'h10 ;
			data[15482] <= 8'h10 ;
			data[15483] <= 8'h10 ;
			data[15484] <= 8'h10 ;
			data[15485] <= 8'h10 ;
			data[15486] <= 8'h10 ;
			data[15487] <= 8'h10 ;
			data[15488] <= 8'h10 ;
			data[15489] <= 8'h10 ;
			data[15490] <= 8'h10 ;
			data[15491] <= 8'h10 ;
			data[15492] <= 8'h10 ;
			data[15493] <= 8'h10 ;
			data[15494] <= 8'h10 ;
			data[15495] <= 8'h10 ;
			data[15496] <= 8'h10 ;
			data[15497] <= 8'h10 ;
			data[15498] <= 8'h10 ;
			data[15499] <= 8'h10 ;
			data[15500] <= 8'h10 ;
			data[15501] <= 8'h10 ;
			data[15502] <= 8'h10 ;
			data[15503] <= 8'h10 ;
			data[15504] <= 8'h10 ;
			data[15505] <= 8'h10 ;
			data[15506] <= 8'h10 ;
			data[15507] <= 8'h10 ;
			data[15508] <= 8'h10 ;
			data[15509] <= 8'h10 ;
			data[15510] <= 8'h10 ;
			data[15511] <= 8'h10 ;
			data[15512] <= 8'h10 ;
			data[15513] <= 8'h10 ;
			data[15514] <= 8'h10 ;
			data[15515] <= 8'h10 ;
			data[15516] <= 8'h10 ;
			data[15517] <= 8'h10 ;
			data[15518] <= 8'h10 ;
			data[15519] <= 8'h10 ;
			data[15520] <= 8'h10 ;
			data[15521] <= 8'h10 ;
			data[15522] <= 8'h10 ;
			data[15523] <= 8'h10 ;
			data[15524] <= 8'h10 ;
			data[15525] <= 8'h10 ;
			data[15526] <= 8'h10 ;
			data[15527] <= 8'h10 ;
			data[15528] <= 8'h10 ;
			data[15529] <= 8'h10 ;
			data[15530] <= 8'h10 ;
			data[15531] <= 8'h10 ;
			data[15532] <= 8'h10 ;
			data[15533] <= 8'h10 ;
			data[15534] <= 8'h10 ;
			data[15535] <= 8'h10 ;
			data[15536] <= 8'h10 ;
			data[15537] <= 8'h10 ;
			data[15538] <= 8'h10 ;
			data[15539] <= 8'h10 ;
			data[15540] <= 8'h10 ;
			data[15541] <= 8'h10 ;
			data[15542] <= 8'h10 ;
			data[15543] <= 8'h10 ;
			data[15544] <= 8'h10 ;
			data[15545] <= 8'h10 ;
			data[15546] <= 8'h10 ;
			data[15547] <= 8'h10 ;
			data[15548] <= 8'h10 ;
			data[15549] <= 8'h10 ;
			data[15550] <= 8'h10 ;
			data[15551] <= 8'h10 ;
			data[15552] <= 8'h10 ;
			data[15553] <= 8'h10 ;
			data[15554] <= 8'h10 ;
			data[15555] <= 8'h10 ;
			data[15556] <= 8'h10 ;
			data[15557] <= 8'h10 ;
			data[15558] <= 8'h10 ;
			data[15559] <= 8'h10 ;
			data[15560] <= 8'h10 ;
			data[15561] <= 8'h10 ;
			data[15562] <= 8'h10 ;
			data[15563] <= 8'h10 ;
			data[15564] <= 8'h10 ;
			data[15565] <= 8'h10 ;
			data[15566] <= 8'h10 ;
			data[15567] <= 8'h10 ;
			data[15568] <= 8'h10 ;
			data[15569] <= 8'h10 ;
			data[15570] <= 8'h10 ;
			data[15571] <= 8'h10 ;
			data[15572] <= 8'h10 ;
			data[15573] <= 8'h10 ;
			data[15574] <= 8'h10 ;
			data[15575] <= 8'h10 ;
			data[15576] <= 8'h10 ;
			data[15577] <= 8'h10 ;
			data[15578] <= 8'h10 ;
			data[15579] <= 8'h10 ;
			data[15580] <= 8'h10 ;
			data[15581] <= 8'h10 ;
			data[15582] <= 8'h10 ;
			data[15583] <= 8'h10 ;
			data[15584] <= 8'h10 ;
			data[15585] <= 8'h10 ;
			data[15586] <= 8'h10 ;
			data[15587] <= 8'h10 ;
			data[15588] <= 8'h10 ;
			data[15589] <= 8'h10 ;
			data[15590] <= 8'h10 ;
			data[15591] <= 8'h10 ;
			data[15592] <= 8'h10 ;
			data[15593] <= 8'h10 ;
			data[15594] <= 8'h10 ;
			data[15595] <= 8'h10 ;
			data[15596] <= 8'h10 ;
			data[15597] <= 8'h10 ;
			data[15598] <= 8'h10 ;
			data[15599] <= 8'h10 ;
			data[15600] <= 8'h10 ;
			data[15601] <= 8'h10 ;
			data[15602] <= 8'h10 ;
			data[15603] <= 8'h10 ;
			data[15604] <= 8'h10 ;
			data[15605] <= 8'h10 ;
			data[15606] <= 8'h10 ;
			data[15607] <= 8'h10 ;
			data[15608] <= 8'h10 ;
			data[15609] <= 8'h10 ;
			data[15610] <= 8'h10 ;
			data[15611] <= 8'h10 ;
			data[15612] <= 8'h10 ;
			data[15613] <= 8'h10 ;
			data[15614] <= 8'h10 ;
			data[15615] <= 8'h10 ;
			data[15616] <= 8'h10 ;
			data[15617] <= 8'h10 ;
			data[15618] <= 8'h10 ;
			data[15619] <= 8'h10 ;
			data[15620] <= 8'h10 ;
			data[15621] <= 8'h10 ;
			data[15622] <= 8'h10 ;
			data[15623] <= 8'h10 ;
			data[15624] <= 8'h10 ;
			data[15625] <= 8'h10 ;
			data[15626] <= 8'h10 ;
			data[15627] <= 8'h10 ;
			data[15628] <= 8'h10 ;
			data[15629] <= 8'h10 ;
			data[15630] <= 8'h10 ;
			data[15631] <= 8'h10 ;
			data[15632] <= 8'h10 ;
			data[15633] <= 8'h10 ;
			data[15634] <= 8'h10 ;
			data[15635] <= 8'h10 ;
			data[15636] <= 8'h10 ;
			data[15637] <= 8'h10 ;
			data[15638] <= 8'h10 ;
			data[15639] <= 8'h10 ;
			data[15640] <= 8'h10 ;
			data[15641] <= 8'h10 ;
			data[15642] <= 8'h10 ;
			data[15643] <= 8'h10 ;
			data[15644] <= 8'h10 ;
			data[15645] <= 8'h10 ;
			data[15646] <= 8'h10 ;
			data[15647] <= 8'h10 ;
			data[15648] <= 8'h10 ;
			data[15649] <= 8'h10 ;
			data[15650] <= 8'h10 ;
			data[15651] <= 8'h10 ;
			data[15652] <= 8'h10 ;
			data[15653] <= 8'h10 ;
			data[15654] <= 8'h10 ;
			data[15655] <= 8'h10 ;
			data[15656] <= 8'h10 ;
			data[15657] <= 8'h10 ;
			data[15658] <= 8'h10 ;
			data[15659] <= 8'h10 ;
			data[15660] <= 8'h10 ;
			data[15661] <= 8'h10 ;
			data[15662] <= 8'h10 ;
			data[15663] <= 8'h10 ;
			data[15664] <= 8'h10 ;
			data[15665] <= 8'h10 ;
			data[15666] <= 8'h10 ;
			data[15667] <= 8'h10 ;
			data[15668] <= 8'h10 ;
			data[15669] <= 8'h10 ;
			data[15670] <= 8'h10 ;
			data[15671] <= 8'h10 ;
			data[15672] <= 8'h10 ;
			data[15673] <= 8'h10 ;
			data[15674] <= 8'h10 ;
			data[15675] <= 8'h10 ;
			data[15676] <= 8'h10 ;
			data[15677] <= 8'h10 ;
			data[15678] <= 8'h10 ;
			data[15679] <= 8'h10 ;
			data[15680] <= 8'h10 ;
			data[15681] <= 8'h10 ;
			data[15682] <= 8'h10 ;
			data[15683] <= 8'h10 ;
			data[15684] <= 8'h10 ;
			data[15685] <= 8'h10 ;
			data[15686] <= 8'h10 ;
			data[15687] <= 8'h10 ;
			data[15688] <= 8'h10 ;
			data[15689] <= 8'h10 ;
			data[15690] <= 8'h10 ;
			data[15691] <= 8'h10 ;
			data[15692] <= 8'h10 ;
			data[15693] <= 8'h10 ;
			data[15694] <= 8'h10 ;
			data[15695] <= 8'h10 ;
			data[15696] <= 8'h10 ;
			data[15697] <= 8'h10 ;
			data[15698] <= 8'h10 ;
			data[15699] <= 8'h10 ;
			data[15700] <= 8'h10 ;
			data[15701] <= 8'h10 ;
			data[15702] <= 8'h10 ;
			data[15703] <= 8'h10 ;
			data[15704] <= 8'h10 ;
			data[15705] <= 8'h10 ;
			data[15706] <= 8'h10 ;
			data[15707] <= 8'h10 ;
			data[15708] <= 8'h10 ;
			data[15709] <= 8'h10 ;
			data[15710] <= 8'h10 ;
			data[15711] <= 8'h10 ;
			data[15712] <= 8'h10 ;
			data[15713] <= 8'h10 ;
			data[15714] <= 8'h10 ;
			data[15715] <= 8'h10 ;
			data[15716] <= 8'h10 ;
			data[15717] <= 8'h10 ;
			data[15718] <= 8'h10 ;
			data[15719] <= 8'h10 ;
			data[15720] <= 8'h10 ;
			data[15721] <= 8'h10 ;
			data[15722] <= 8'h10 ;
			data[15723] <= 8'h10 ;
			data[15724] <= 8'h10 ;
			data[15725] <= 8'h10 ;
			data[15726] <= 8'h10 ;
			data[15727] <= 8'h10 ;
			data[15728] <= 8'h10 ;
			data[15729] <= 8'h10 ;
			data[15730] <= 8'h10 ;
			data[15731] <= 8'h10 ;
			data[15732] <= 8'h10 ;
			data[15733] <= 8'h10 ;
			data[15734] <= 8'h10 ;
			data[15735] <= 8'h10 ;
			data[15736] <= 8'h10 ;
			data[15737] <= 8'h10 ;
			data[15738] <= 8'h10 ;
			data[15739] <= 8'h10 ;
			data[15740] <= 8'h10 ;
			data[15741] <= 8'h10 ;
			data[15742] <= 8'h10 ;
			data[15743] <= 8'h10 ;
			data[15744] <= 8'h10 ;
			data[15745] <= 8'h10 ;
			data[15746] <= 8'h10 ;
			data[15747] <= 8'h10 ;
			data[15748] <= 8'h10 ;
			data[15749] <= 8'h10 ;
			data[15750] <= 8'h10 ;
			data[15751] <= 8'h10 ;
			data[15752] <= 8'h10 ;
			data[15753] <= 8'h10 ;
			data[15754] <= 8'h10 ;
			data[15755] <= 8'h10 ;
			data[15756] <= 8'h10 ;
			data[15757] <= 8'h10 ;
			data[15758] <= 8'h10 ;
			data[15759] <= 8'h10 ;
			data[15760] <= 8'h10 ;
			data[15761] <= 8'h10 ;
			data[15762] <= 8'h10 ;
			data[15763] <= 8'h10 ;
			data[15764] <= 8'h10 ;
			data[15765] <= 8'h10 ;
			data[15766] <= 8'h10 ;
			data[15767] <= 8'h10 ;
			data[15768] <= 8'h10 ;
			data[15769] <= 8'h10 ;
			data[15770] <= 8'h10 ;
			data[15771] <= 8'h10 ;
			data[15772] <= 8'h10 ;
			data[15773] <= 8'h10 ;
			data[15774] <= 8'h10 ;
			data[15775] <= 8'h10 ;
			data[15776] <= 8'h10 ;
			data[15777] <= 8'h10 ;
			data[15778] <= 8'h10 ;
			data[15779] <= 8'h10 ;
			data[15780] <= 8'h10 ;
			data[15781] <= 8'h10 ;
			data[15782] <= 8'h10 ;
			data[15783] <= 8'h10 ;
			data[15784] <= 8'h10 ;
			data[15785] <= 8'h10 ;
			data[15786] <= 8'h10 ;
			data[15787] <= 8'h10 ;
			data[15788] <= 8'h10 ;
			data[15789] <= 8'h10 ;
			data[15790] <= 8'h10 ;
			data[15791] <= 8'h10 ;
			data[15792] <= 8'h10 ;
			data[15793] <= 8'h10 ;
			data[15794] <= 8'h10 ;
			data[15795] <= 8'h10 ;
			data[15796] <= 8'h10 ;
			data[15797] <= 8'h10 ;
			data[15798] <= 8'h10 ;
			data[15799] <= 8'h10 ;
			data[15800] <= 8'h10 ;
			data[15801] <= 8'h10 ;
			data[15802] <= 8'h10 ;
			data[15803] <= 8'h10 ;
			data[15804] <= 8'h10 ;
			data[15805] <= 8'h10 ;
			data[15806] <= 8'h10 ;
			data[15807] <= 8'h10 ;
			data[15808] <= 8'h10 ;
			data[15809] <= 8'h10 ;
			data[15810] <= 8'h10 ;
			data[15811] <= 8'h10 ;
			data[15812] <= 8'h10 ;
			data[15813] <= 8'h10 ;
			data[15814] <= 8'h10 ;
			data[15815] <= 8'h10 ;
			data[15816] <= 8'h10 ;
			data[15817] <= 8'h10 ;
			data[15818] <= 8'h10 ;
			data[15819] <= 8'h10 ;
			data[15820] <= 8'h10 ;
			data[15821] <= 8'h10 ;
			data[15822] <= 8'h10 ;
			data[15823] <= 8'h10 ;
			data[15824] <= 8'h10 ;
			data[15825] <= 8'h10 ;
			data[15826] <= 8'h10 ;
			data[15827] <= 8'h10 ;
			data[15828] <= 8'h10 ;
			data[15829] <= 8'h10 ;
			data[15830] <= 8'h10 ;
			data[15831] <= 8'h10 ;
			data[15832] <= 8'h10 ;
			data[15833] <= 8'h10 ;
			data[15834] <= 8'h10 ;
			data[15835] <= 8'h10 ;
			data[15836] <= 8'h10 ;
			data[15837] <= 8'h10 ;
			data[15838] <= 8'h10 ;
			data[15839] <= 8'h10 ;
			data[15840] <= 8'h10 ;
			data[15841] <= 8'h10 ;
			data[15842] <= 8'h10 ;
			data[15843] <= 8'h10 ;
			data[15844] <= 8'h10 ;
			data[15845] <= 8'h10 ;
			data[15846] <= 8'h10 ;
			data[15847] <= 8'h10 ;
			data[15848] <= 8'h10 ;
			data[15849] <= 8'h10 ;
			data[15850] <= 8'h10 ;
			data[15851] <= 8'h10 ;
			data[15852] <= 8'h10 ;
			data[15853] <= 8'h10 ;
			data[15854] <= 8'h10 ;
			data[15855] <= 8'h10 ;
			data[15856] <= 8'h10 ;
			data[15857] <= 8'h10 ;
			data[15858] <= 8'h10 ;
			data[15859] <= 8'h10 ;
			data[15860] <= 8'h10 ;
			data[15861] <= 8'h10 ;
			data[15862] <= 8'h10 ;
			data[15863] <= 8'h10 ;
			data[15864] <= 8'h10 ;
			data[15865] <= 8'h10 ;
			data[15866] <= 8'h10 ;
			data[15867] <= 8'h10 ;
			data[15868] <= 8'h10 ;
			data[15869] <= 8'h10 ;
			data[15870] <= 8'h10 ;
			data[15871] <= 8'h10 ;
			data[15872] <= 8'h10 ;
			data[15873] <= 8'h10 ;
			data[15874] <= 8'h10 ;
			data[15875] <= 8'h10 ;
			data[15876] <= 8'h10 ;
			data[15877] <= 8'h10 ;
			data[15878] <= 8'h10 ;
			data[15879] <= 8'h10 ;
			data[15880] <= 8'h10 ;
			data[15881] <= 8'h10 ;
			data[15882] <= 8'h10 ;
			data[15883] <= 8'h10 ;
			data[15884] <= 8'h10 ;
			data[15885] <= 8'h10 ;
			data[15886] <= 8'h10 ;
			data[15887] <= 8'h10 ;
			data[15888] <= 8'h10 ;
			data[15889] <= 8'h10 ;
			data[15890] <= 8'h10 ;
			data[15891] <= 8'h10 ;
			data[15892] <= 8'h10 ;
			data[15893] <= 8'h10 ;
			data[15894] <= 8'h10 ;
			data[15895] <= 8'h10 ;
			data[15896] <= 8'h10 ;
			data[15897] <= 8'h10 ;
			data[15898] <= 8'h10 ;
			data[15899] <= 8'h10 ;
			data[15900] <= 8'h10 ;
			data[15901] <= 8'h10 ;
			data[15902] <= 8'h10 ;
			data[15903] <= 8'h10 ;
			data[15904] <= 8'h10 ;
			data[15905] <= 8'h10 ;
			data[15906] <= 8'h10 ;
			data[15907] <= 8'h10 ;
			data[15908] <= 8'h10 ;
			data[15909] <= 8'h10 ;
			data[15910] <= 8'h10 ;
			data[15911] <= 8'h10 ;
			data[15912] <= 8'h10 ;
			data[15913] <= 8'h10 ;
			data[15914] <= 8'h10 ;
			data[15915] <= 8'h10 ;
			data[15916] <= 8'h10 ;
			data[15917] <= 8'h10 ;
			data[15918] <= 8'h10 ;
			data[15919] <= 8'h10 ;
			data[15920] <= 8'h10 ;
			data[15921] <= 8'h10 ;
			data[15922] <= 8'h10 ;
			data[15923] <= 8'h10 ;
			data[15924] <= 8'h10 ;
			data[15925] <= 8'h10 ;
			data[15926] <= 8'h10 ;
			data[15927] <= 8'h10 ;
			data[15928] <= 8'h10 ;
			data[15929] <= 8'h10 ;
			data[15930] <= 8'h10 ;
			data[15931] <= 8'h10 ;
			data[15932] <= 8'h10 ;
			data[15933] <= 8'h10 ;
			data[15934] <= 8'h10 ;
			data[15935] <= 8'h10 ;
			data[15936] <= 8'h10 ;
			data[15937] <= 8'h10 ;
			data[15938] <= 8'h10 ;
			data[15939] <= 8'h10 ;
			data[15940] <= 8'h10 ;
			data[15941] <= 8'h10 ;
			data[15942] <= 8'h10 ;
			data[15943] <= 8'h10 ;
			data[15944] <= 8'h10 ;
			data[15945] <= 8'h10 ;
			data[15946] <= 8'h10 ;
			data[15947] <= 8'h10 ;
			data[15948] <= 8'h10 ;
			data[15949] <= 8'h10 ;
			data[15950] <= 8'h10 ;
			data[15951] <= 8'h10 ;
			data[15952] <= 8'h10 ;
			data[15953] <= 8'h10 ;
			data[15954] <= 8'h10 ;
			data[15955] <= 8'h10 ;
			data[15956] <= 8'h10 ;
			data[15957] <= 8'h10 ;
			data[15958] <= 8'h10 ;
			data[15959] <= 8'h10 ;
			data[15960] <= 8'h10 ;
			data[15961] <= 8'h10 ;
			data[15962] <= 8'h10 ;
			data[15963] <= 8'h10 ;
			data[15964] <= 8'h10 ;
			data[15965] <= 8'h10 ;
			data[15966] <= 8'h10 ;
			data[15967] <= 8'h10 ;
			data[15968] <= 8'h10 ;
			data[15969] <= 8'h10 ;
			data[15970] <= 8'h10 ;
			data[15971] <= 8'h10 ;
			data[15972] <= 8'h10 ;
			data[15973] <= 8'h10 ;
			data[15974] <= 8'h10 ;
			data[15975] <= 8'h10 ;
			data[15976] <= 8'h10 ;
			data[15977] <= 8'h10 ;
			data[15978] <= 8'h10 ;
			data[15979] <= 8'h10 ;
			data[15980] <= 8'h10 ;
			data[15981] <= 8'h10 ;
			data[15982] <= 8'h10 ;
			data[15983] <= 8'h10 ;
			data[15984] <= 8'h10 ;
			data[15985] <= 8'h10 ;
			data[15986] <= 8'h10 ;
			data[15987] <= 8'h10 ;
			data[15988] <= 8'h10 ;
			data[15989] <= 8'h10 ;
			data[15990] <= 8'h10 ;
			data[15991] <= 8'h10 ;
			data[15992] <= 8'h10 ;
			data[15993] <= 8'h10 ;
			data[15994] <= 8'h10 ;
			data[15995] <= 8'h10 ;
			data[15996] <= 8'h10 ;
			data[15997] <= 8'h10 ;
			data[15998] <= 8'h10 ;
			data[15999] <= 8'h10 ;
			data[16000] <= 8'h10 ;
			data[16001] <= 8'h10 ;
			data[16002] <= 8'h10 ;
			data[16003] <= 8'h10 ;
			data[16004] <= 8'h10 ;
			data[16005] <= 8'h10 ;
			data[16006] <= 8'h10 ;
			data[16007] <= 8'h10 ;
			data[16008] <= 8'h10 ;
			data[16009] <= 8'h10 ;
			data[16010] <= 8'h10 ;
			data[16011] <= 8'h10 ;
			data[16012] <= 8'h10 ;
			data[16013] <= 8'h10 ;
			data[16014] <= 8'h10 ;
			data[16015] <= 8'h10 ;
			data[16016] <= 8'h10 ;
			data[16017] <= 8'h10 ;
			data[16018] <= 8'h10 ;
			data[16019] <= 8'h10 ;
			data[16020] <= 8'h10 ;
			data[16021] <= 8'h10 ;
			data[16022] <= 8'h10 ;
			data[16023] <= 8'h10 ;
			data[16024] <= 8'h10 ;
			data[16025] <= 8'h10 ;
			data[16026] <= 8'h10 ;
			data[16027] <= 8'h10 ;
			data[16028] <= 8'h10 ;
			data[16029] <= 8'h10 ;
			data[16030] <= 8'h10 ;
			data[16031] <= 8'h10 ;
			data[16032] <= 8'h10 ;
			data[16033] <= 8'h10 ;
			data[16034] <= 8'h10 ;
			data[16035] <= 8'h10 ;
			data[16036] <= 8'h10 ;
			data[16037] <= 8'h10 ;
			data[16038] <= 8'h10 ;
			data[16039] <= 8'h10 ;
			data[16040] <= 8'h10 ;
			data[16041] <= 8'h10 ;
			data[16042] <= 8'h10 ;
			data[16043] <= 8'h10 ;
			data[16044] <= 8'h10 ;
			data[16045] <= 8'h10 ;
			data[16046] <= 8'h10 ;
			data[16047] <= 8'h10 ;
			data[16048] <= 8'h10 ;
			data[16049] <= 8'h10 ;
			data[16050] <= 8'h10 ;
			data[16051] <= 8'h10 ;
			data[16052] <= 8'h10 ;
			data[16053] <= 8'h10 ;
			data[16054] <= 8'h10 ;
			data[16055] <= 8'h10 ;
			data[16056] <= 8'h10 ;
			data[16057] <= 8'h10 ;
			data[16058] <= 8'h10 ;
			data[16059] <= 8'h10 ;
			data[16060] <= 8'h10 ;
			data[16061] <= 8'h10 ;
			data[16062] <= 8'h10 ;
			data[16063] <= 8'h10 ;
			data[16064] <= 8'h10 ;
			data[16065] <= 8'h10 ;
			data[16066] <= 8'h10 ;
			data[16067] <= 8'h10 ;
			data[16068] <= 8'h10 ;
			data[16069] <= 8'h10 ;
			data[16070] <= 8'h10 ;
			data[16071] <= 8'h10 ;
			data[16072] <= 8'h10 ;
			data[16073] <= 8'h10 ;
			data[16074] <= 8'h10 ;
			data[16075] <= 8'h10 ;
			data[16076] <= 8'h10 ;
			data[16077] <= 8'h10 ;
			data[16078] <= 8'h10 ;
			data[16079] <= 8'h10 ;
			data[16080] <= 8'h10 ;
			data[16081] <= 8'h10 ;
			data[16082] <= 8'h10 ;
			data[16083] <= 8'h10 ;
			data[16084] <= 8'h10 ;
			data[16085] <= 8'h10 ;
			data[16086] <= 8'h10 ;
			data[16087] <= 8'h10 ;
			data[16088] <= 8'h10 ;
			data[16089] <= 8'h10 ;
			data[16090] <= 8'h10 ;
			data[16091] <= 8'h10 ;
			data[16092] <= 8'h10 ;
			data[16093] <= 8'h10 ;
			data[16094] <= 8'h10 ;
			data[16095] <= 8'h10 ;
			data[16096] <= 8'h10 ;
			data[16097] <= 8'h10 ;
			data[16098] <= 8'h10 ;
			data[16099] <= 8'h10 ;
			data[16100] <= 8'h10 ;
			data[16101] <= 8'h10 ;
			data[16102] <= 8'h10 ;
			data[16103] <= 8'h10 ;
			data[16104] <= 8'h10 ;
			data[16105] <= 8'h10 ;
			data[16106] <= 8'h10 ;
			data[16107] <= 8'h10 ;
			data[16108] <= 8'h10 ;
			data[16109] <= 8'h10 ;
			data[16110] <= 8'h10 ;
			data[16111] <= 8'h10 ;
			data[16112] <= 8'h10 ;
			data[16113] <= 8'h10 ;
			data[16114] <= 8'h10 ;
			data[16115] <= 8'h10 ;
			data[16116] <= 8'h10 ;
			data[16117] <= 8'h10 ;
			data[16118] <= 8'h10 ;
			data[16119] <= 8'h10 ;
			data[16120] <= 8'h10 ;
			data[16121] <= 8'h10 ;
			data[16122] <= 8'h10 ;
			data[16123] <= 8'h10 ;
			data[16124] <= 8'h10 ;
			data[16125] <= 8'h10 ;
			data[16126] <= 8'h10 ;
			data[16127] <= 8'h10 ;
			data[16128] <= 8'h10 ;
			data[16129] <= 8'h10 ;
			data[16130] <= 8'h10 ;
			data[16131] <= 8'h10 ;
			data[16132] <= 8'h10 ;
			data[16133] <= 8'h10 ;
			data[16134] <= 8'h10 ;
			data[16135] <= 8'h10 ;
			data[16136] <= 8'h10 ;
			data[16137] <= 8'h10 ;
			data[16138] <= 8'h10 ;
			data[16139] <= 8'h10 ;
			data[16140] <= 8'h10 ;
			data[16141] <= 8'h10 ;
			data[16142] <= 8'h10 ;
			data[16143] <= 8'h10 ;
			data[16144] <= 8'h10 ;
			data[16145] <= 8'h10 ;
			data[16146] <= 8'h10 ;
			data[16147] <= 8'h10 ;
			data[16148] <= 8'h10 ;
			data[16149] <= 8'h10 ;
			data[16150] <= 8'h10 ;
			data[16151] <= 8'h10 ;
			data[16152] <= 8'h10 ;
			data[16153] <= 8'h10 ;
			data[16154] <= 8'h10 ;
			data[16155] <= 8'h10 ;
			data[16156] <= 8'h10 ;
			data[16157] <= 8'h10 ;
			data[16158] <= 8'h10 ;
			data[16159] <= 8'h10 ;
			data[16160] <= 8'h10 ;
			data[16161] <= 8'h10 ;
			data[16162] <= 8'h10 ;
			data[16163] <= 8'h10 ;
			data[16164] <= 8'h10 ;
			data[16165] <= 8'h10 ;
			data[16166] <= 8'h10 ;
			data[16167] <= 8'h10 ;
			data[16168] <= 8'h10 ;
			data[16169] <= 8'h10 ;
			data[16170] <= 8'h10 ;
			data[16171] <= 8'h10 ;
			data[16172] <= 8'h10 ;
			data[16173] <= 8'h10 ;
			data[16174] <= 8'h10 ;
			data[16175] <= 8'h10 ;
			data[16176] <= 8'h10 ;
			data[16177] <= 8'h10 ;
			data[16178] <= 8'h10 ;
			data[16179] <= 8'h10 ;
			data[16180] <= 8'h10 ;
			data[16181] <= 8'h10 ;
			data[16182] <= 8'h10 ;
			data[16183] <= 8'h10 ;
			data[16184] <= 8'h10 ;
			data[16185] <= 8'h10 ;
			data[16186] <= 8'h10 ;
			data[16187] <= 8'h10 ;
			data[16188] <= 8'h10 ;
			data[16189] <= 8'h10 ;
			data[16190] <= 8'h10 ;
			data[16191] <= 8'h10 ;
			data[16192] <= 8'h10 ;
			data[16193] <= 8'h10 ;
			data[16194] <= 8'h10 ;
			data[16195] <= 8'h10 ;
			data[16196] <= 8'h10 ;
			data[16197] <= 8'h10 ;
			data[16198] <= 8'h10 ;
			data[16199] <= 8'h10 ;
			data[16200] <= 8'h10 ;
			data[16201] <= 8'h10 ;
			data[16202] <= 8'h10 ;
			data[16203] <= 8'h10 ;
			data[16204] <= 8'h10 ;
			data[16205] <= 8'h10 ;
			data[16206] <= 8'h10 ;
			data[16207] <= 8'h10 ;
			data[16208] <= 8'h10 ;
			data[16209] <= 8'h10 ;
			data[16210] <= 8'h10 ;
			data[16211] <= 8'h10 ;
			data[16212] <= 8'h10 ;
			data[16213] <= 8'h10 ;
			data[16214] <= 8'h10 ;
			data[16215] <= 8'h10 ;
			data[16216] <= 8'h10 ;
			data[16217] <= 8'h10 ;
			data[16218] <= 8'h10 ;
			data[16219] <= 8'h10 ;
			data[16220] <= 8'h10 ;
			data[16221] <= 8'h10 ;
			data[16222] <= 8'h10 ;
			data[16223] <= 8'h10 ;
			data[16224] <= 8'h10 ;
			data[16225] <= 8'h10 ;
			data[16226] <= 8'h10 ;
			data[16227] <= 8'h10 ;
			data[16228] <= 8'h10 ;
			data[16229] <= 8'h10 ;
			data[16230] <= 8'h10 ;
			data[16231] <= 8'h10 ;
			data[16232] <= 8'h10 ;
			data[16233] <= 8'h10 ;
			data[16234] <= 8'h10 ;
			data[16235] <= 8'h10 ;
			data[16236] <= 8'h10 ;
			data[16237] <= 8'h10 ;
			data[16238] <= 8'h10 ;
			data[16239] <= 8'h10 ;
			data[16240] <= 8'h10 ;
			data[16241] <= 8'h10 ;
			data[16242] <= 8'h10 ;
			data[16243] <= 8'h10 ;
			data[16244] <= 8'h10 ;
			data[16245] <= 8'h10 ;
			data[16246] <= 8'h10 ;
			data[16247] <= 8'h10 ;
			data[16248] <= 8'h10 ;
			data[16249] <= 8'h10 ;
			data[16250] <= 8'h10 ;
			data[16251] <= 8'h10 ;
			data[16252] <= 8'h10 ;
			data[16253] <= 8'h10 ;
			data[16254] <= 8'h10 ;
			data[16255] <= 8'h10 ;
			data[16256] <= 8'h10 ;
			data[16257] <= 8'h10 ;
			data[16258] <= 8'h10 ;
			data[16259] <= 8'h10 ;
			data[16260] <= 8'h10 ;
			data[16261] <= 8'h10 ;
			data[16262] <= 8'h10 ;
			data[16263] <= 8'h10 ;
			data[16264] <= 8'h10 ;
			data[16265] <= 8'h10 ;
			data[16266] <= 8'h10 ;
			data[16267] <= 8'h10 ;
			data[16268] <= 8'h10 ;
			data[16269] <= 8'h10 ;
			data[16270] <= 8'h10 ;
			data[16271] <= 8'h10 ;
			data[16272] <= 8'h10 ;
			data[16273] <= 8'h10 ;
			data[16274] <= 8'h10 ;
			data[16275] <= 8'h10 ;
			data[16276] <= 8'h10 ;
			data[16277] <= 8'h10 ;
			data[16278] <= 8'h10 ;
			data[16279] <= 8'h10 ;
			data[16280] <= 8'h10 ;
			data[16281] <= 8'h10 ;
			data[16282] <= 8'h10 ;
			data[16283] <= 8'h10 ;
			data[16284] <= 8'h10 ;
			data[16285] <= 8'h10 ;
			data[16286] <= 8'h10 ;
			data[16287] <= 8'h10 ;
			data[16288] <= 8'h10 ;
			data[16289] <= 8'h10 ;
			data[16290] <= 8'h10 ;
			data[16291] <= 8'h10 ;
			data[16292] <= 8'h10 ;
			data[16293] <= 8'h10 ;
			data[16294] <= 8'h10 ;
			data[16295] <= 8'h10 ;
			data[16296] <= 8'h10 ;
			data[16297] <= 8'h10 ;
			data[16298] <= 8'h10 ;
			data[16299] <= 8'h10 ;
			data[16300] <= 8'h10 ;
			data[16301] <= 8'h10 ;
			data[16302] <= 8'h10 ;
			data[16303] <= 8'h10 ;
			data[16304] <= 8'h10 ;
			data[16305] <= 8'h10 ;
			data[16306] <= 8'h10 ;
			data[16307] <= 8'h10 ;
			data[16308] <= 8'h10 ;
			data[16309] <= 8'h10 ;
			data[16310] <= 8'h10 ;
			data[16311] <= 8'h10 ;
			data[16312] <= 8'h10 ;
			data[16313] <= 8'h10 ;
			data[16314] <= 8'h10 ;
			data[16315] <= 8'h10 ;
			data[16316] <= 8'h10 ;
			data[16317] <= 8'h10 ;
			data[16318] <= 8'h10 ;
			data[16319] <= 8'h10 ;
			data[16320] <= 8'h10 ;
			data[16321] <= 8'h10 ;
			data[16322] <= 8'h10 ;
			data[16323] <= 8'h10 ;
			data[16324] <= 8'h10 ;
			data[16325] <= 8'h10 ;
			data[16326] <= 8'h10 ;
			data[16327] <= 8'h10 ;
			data[16328] <= 8'h10 ;
			data[16329] <= 8'h10 ;
			data[16330] <= 8'h10 ;
			data[16331] <= 8'h10 ;
			data[16332] <= 8'h10 ;
			data[16333] <= 8'h10 ;
			data[16334] <= 8'h10 ;
			data[16335] <= 8'h10 ;
			data[16336] <= 8'h10 ;
			data[16337] <= 8'h10 ;
			data[16338] <= 8'h10 ;
			data[16339] <= 8'h10 ;
			data[16340] <= 8'h10 ;
			data[16341] <= 8'h10 ;
			data[16342] <= 8'h10 ;
			data[16343] <= 8'h10 ;
			data[16344] <= 8'h10 ;
			data[16345] <= 8'h10 ;
			data[16346] <= 8'h10 ;
			data[16347] <= 8'h10 ;
			data[16348] <= 8'h10 ;
			data[16349] <= 8'h10 ;
			data[16350] <= 8'h10 ;
			data[16351] <= 8'h10 ;
			data[16352] <= 8'h10 ;
			data[16353] <= 8'h10 ;
			data[16354] <= 8'h10 ;
			data[16355] <= 8'h10 ;
			data[16356] <= 8'h10 ;
			data[16357] <= 8'h10 ;
			data[16358] <= 8'h10 ;
			data[16359] <= 8'h10 ;
			data[16360] <= 8'h10 ;
			data[16361] <= 8'h10 ;
			data[16362] <= 8'h10 ;
			data[16363] <= 8'h10 ;
			data[16364] <= 8'h10 ;
			data[16365] <= 8'h10 ;
			data[16366] <= 8'h10 ;
			data[16367] <= 8'h10 ;
			data[16368] <= 8'h10 ;
			data[16369] <= 8'h10 ;
			data[16370] <= 8'h10 ;
			data[16371] <= 8'h10 ;
			data[16372] <= 8'h10 ;
			data[16373] <= 8'h10 ;
			data[16374] <= 8'h10 ;
			data[16375] <= 8'h10 ;
			data[16376] <= 8'h10 ;
			data[16377] <= 8'h10 ;
			data[16378] <= 8'h10 ;
			data[16379] <= 8'h10 ;
			data[16380] <= 8'h10 ;
			data[16381] <= 8'h10 ;
			data[16382] <= 8'h10 ;
			data[16383] <= 8'h10 ;
			data[16384] <= 8'h10 ;
			data[16385] <= 8'h10 ;
			data[16386] <= 8'h10 ;
			data[16387] <= 8'h10 ;
			data[16388] <= 8'h10 ;
			data[16389] <= 8'h10 ;
			data[16390] <= 8'h10 ;
			data[16391] <= 8'h10 ;
			data[16392] <= 8'h10 ;
			data[16393] <= 8'h10 ;
			data[16394] <= 8'h10 ;
			data[16395] <= 8'h10 ;
			data[16396] <= 8'h10 ;
			data[16397] <= 8'h10 ;
			data[16398] <= 8'h10 ;
			data[16399] <= 8'h10 ;
			data[16400] <= 8'h10 ;
			data[16401] <= 8'h10 ;
			data[16402] <= 8'h10 ;
			data[16403] <= 8'h10 ;
			data[16404] <= 8'h10 ;
			data[16405] <= 8'h10 ;
			data[16406] <= 8'h10 ;
			data[16407] <= 8'h10 ;
			data[16408] <= 8'h10 ;
			data[16409] <= 8'h10 ;
			data[16410] <= 8'h10 ;
			data[16411] <= 8'h10 ;
			data[16412] <= 8'h10 ;
			data[16413] <= 8'h10 ;
			data[16414] <= 8'h10 ;
			data[16415] <= 8'h10 ;
			data[16416] <= 8'h10 ;
			data[16417] <= 8'h10 ;
			data[16418] <= 8'h10 ;
			data[16419] <= 8'h10 ;
			data[16420] <= 8'h10 ;
			data[16421] <= 8'h10 ;
			data[16422] <= 8'h10 ;
			data[16423] <= 8'h10 ;
			data[16424] <= 8'h10 ;
			data[16425] <= 8'h10 ;
			data[16426] <= 8'h10 ;
			data[16427] <= 8'h10 ;
			data[16428] <= 8'h10 ;
			data[16429] <= 8'h10 ;
			data[16430] <= 8'h10 ;
			data[16431] <= 8'h10 ;
			data[16432] <= 8'h10 ;
			data[16433] <= 8'h10 ;
			data[16434] <= 8'h10 ;
			data[16435] <= 8'h10 ;
			data[16436] <= 8'h10 ;
			data[16437] <= 8'h10 ;
			data[16438] <= 8'h10 ;
			data[16439] <= 8'h10 ;
			data[16440] <= 8'h10 ;
			data[16441] <= 8'h10 ;
			data[16442] <= 8'h10 ;
			data[16443] <= 8'h10 ;
			data[16444] <= 8'h10 ;
			data[16445] <= 8'h10 ;
			data[16446] <= 8'h10 ;
			data[16447] <= 8'h10 ;
			data[16448] <= 8'h10 ;
			data[16449] <= 8'h10 ;
			data[16450] <= 8'h10 ;
			data[16451] <= 8'h10 ;
			data[16452] <= 8'h10 ;
			data[16453] <= 8'h10 ;
			data[16454] <= 8'h10 ;
			data[16455] <= 8'h10 ;
			data[16456] <= 8'h10 ;
			data[16457] <= 8'h10 ;
			data[16458] <= 8'h10 ;
			data[16459] <= 8'h10 ;
			data[16460] <= 8'h10 ;
			data[16461] <= 8'h10 ;
			data[16462] <= 8'h10 ;
			data[16463] <= 8'h10 ;
			data[16464] <= 8'h10 ;
			data[16465] <= 8'h10 ;
			data[16466] <= 8'h10 ;
			data[16467] <= 8'h10 ;
			data[16468] <= 8'h10 ;
			data[16469] <= 8'h10 ;
			data[16470] <= 8'h10 ;
			data[16471] <= 8'h10 ;
			data[16472] <= 8'h10 ;
			data[16473] <= 8'h10 ;
			data[16474] <= 8'h10 ;
			data[16475] <= 8'h10 ;
			data[16476] <= 8'h10 ;
			data[16477] <= 8'h10 ;
			data[16478] <= 8'h10 ;
			data[16479] <= 8'h10 ;
			data[16480] <= 8'h10 ;
			data[16481] <= 8'h10 ;
			data[16482] <= 8'h10 ;
			data[16483] <= 8'h10 ;
			data[16484] <= 8'h10 ;
			data[16485] <= 8'h10 ;
			data[16486] <= 8'h10 ;
			data[16487] <= 8'h10 ;
			data[16488] <= 8'h10 ;
			data[16489] <= 8'h10 ;
			data[16490] <= 8'h10 ;
			data[16491] <= 8'h10 ;
			data[16492] <= 8'h10 ;
			data[16493] <= 8'h10 ;
			data[16494] <= 8'h10 ;
			data[16495] <= 8'h10 ;
			data[16496] <= 8'h10 ;
			data[16497] <= 8'h10 ;
			data[16498] <= 8'h10 ;
			data[16499] <= 8'h10 ;
			data[16500] <= 8'h10 ;
			data[16501] <= 8'h10 ;
			data[16502] <= 8'h10 ;
			data[16503] <= 8'h10 ;
			data[16504] <= 8'h10 ;
			data[16505] <= 8'h10 ;
			data[16506] <= 8'h10 ;
			data[16507] <= 8'h10 ;
			data[16508] <= 8'h10 ;
			data[16509] <= 8'h10 ;
			data[16510] <= 8'h10 ;
			data[16511] <= 8'h10 ;
			data[16512] <= 8'h10 ;
			data[16513] <= 8'h10 ;
			data[16514] <= 8'h10 ;
			data[16515] <= 8'h10 ;
			data[16516] <= 8'h10 ;
			data[16517] <= 8'h10 ;
			data[16518] <= 8'h10 ;
			data[16519] <= 8'h10 ;
			data[16520] <= 8'h10 ;
			data[16521] <= 8'h10 ;
			data[16522] <= 8'h10 ;
			data[16523] <= 8'h10 ;
			data[16524] <= 8'h10 ;
			data[16525] <= 8'h10 ;
			data[16526] <= 8'h10 ;
			data[16527] <= 8'h10 ;
			data[16528] <= 8'h10 ;
			data[16529] <= 8'h10 ;
			data[16530] <= 8'h10 ;
			data[16531] <= 8'h10 ;
			data[16532] <= 8'h10 ;
			data[16533] <= 8'h10 ;
			data[16534] <= 8'h10 ;
			data[16535] <= 8'h10 ;
			data[16536] <= 8'h10 ;
			data[16537] <= 8'h10 ;
			data[16538] <= 8'h10 ;
			data[16539] <= 8'h10 ;
			data[16540] <= 8'h10 ;
			data[16541] <= 8'h10 ;
			data[16542] <= 8'h10 ;
			data[16543] <= 8'h10 ;
			data[16544] <= 8'h10 ;
			data[16545] <= 8'h10 ;
			data[16546] <= 8'h10 ;
			data[16547] <= 8'h10 ;
			data[16548] <= 8'h10 ;
			data[16549] <= 8'h10 ;
			data[16550] <= 8'h10 ;
			data[16551] <= 8'h10 ;
			data[16552] <= 8'h10 ;
			data[16553] <= 8'h10 ;
			data[16554] <= 8'h10 ;
			data[16555] <= 8'h10 ;
			data[16556] <= 8'h10 ;
			data[16557] <= 8'h10 ;
			data[16558] <= 8'h10 ;
			data[16559] <= 8'h10 ;
			data[16560] <= 8'h10 ;
			data[16561] <= 8'h10 ;
			data[16562] <= 8'h10 ;
			data[16563] <= 8'h10 ;
			data[16564] <= 8'h10 ;
			data[16565] <= 8'h10 ;
			data[16566] <= 8'h10 ;
			data[16567] <= 8'h10 ;
			data[16568] <= 8'h10 ;
			data[16569] <= 8'h10 ;
			data[16570] <= 8'h10 ;
			data[16571] <= 8'h10 ;
			data[16572] <= 8'h10 ;
			data[16573] <= 8'h10 ;
			data[16574] <= 8'h10 ;
			data[16575] <= 8'h10 ;
			data[16576] <= 8'h10 ;
			data[16577] <= 8'h10 ;
			data[16578] <= 8'h10 ;
			data[16579] <= 8'h10 ;
			data[16580] <= 8'h10 ;
			data[16581] <= 8'h10 ;
			data[16582] <= 8'h10 ;
			data[16583] <= 8'h10 ;
			data[16584] <= 8'h10 ;
			data[16585] <= 8'h10 ;
			data[16586] <= 8'h10 ;
			data[16587] <= 8'h10 ;
			data[16588] <= 8'h10 ;
			data[16589] <= 8'h10 ;
			data[16590] <= 8'h10 ;
			data[16591] <= 8'h10 ;
			data[16592] <= 8'h10 ;
			data[16593] <= 8'h10 ;
			data[16594] <= 8'h10 ;
			data[16595] <= 8'h10 ;
			data[16596] <= 8'h10 ;
			data[16597] <= 8'h10 ;
			data[16598] <= 8'h10 ;
			data[16599] <= 8'h10 ;
			data[16600] <= 8'h10 ;
			data[16601] <= 8'h10 ;
			data[16602] <= 8'h10 ;
			data[16603] <= 8'h10 ;
			data[16604] <= 8'h10 ;
			data[16605] <= 8'h10 ;
			data[16606] <= 8'h10 ;
			data[16607] <= 8'h10 ;
			data[16608] <= 8'h10 ;
			data[16609] <= 8'h10 ;
			data[16610] <= 8'h10 ;
			data[16611] <= 8'h10 ;
			data[16612] <= 8'h10 ;
			data[16613] <= 8'h10 ;
			data[16614] <= 8'h10 ;
			data[16615] <= 8'h10 ;
			data[16616] <= 8'h10 ;
			data[16617] <= 8'h10 ;
			data[16618] <= 8'h10 ;
			data[16619] <= 8'h10 ;
			data[16620] <= 8'h10 ;
			data[16621] <= 8'h10 ;
			data[16622] <= 8'h10 ;
			data[16623] <= 8'h10 ;
			data[16624] <= 8'h10 ;
			data[16625] <= 8'h10 ;
			data[16626] <= 8'h10 ;
			data[16627] <= 8'h10 ;
			data[16628] <= 8'h10 ;
			data[16629] <= 8'h10 ;
			data[16630] <= 8'h10 ;
			data[16631] <= 8'h10 ;
			data[16632] <= 8'h10 ;
			data[16633] <= 8'h10 ;
			data[16634] <= 8'h10 ;
			data[16635] <= 8'h10 ;
			data[16636] <= 8'h10 ;
			data[16637] <= 8'h10 ;
			data[16638] <= 8'h10 ;
			data[16639] <= 8'h10 ;
			data[16640] <= 8'h10 ;
			data[16641] <= 8'h10 ;
			data[16642] <= 8'h10 ;
			data[16643] <= 8'h10 ;
			data[16644] <= 8'h10 ;
			data[16645] <= 8'h10 ;
			data[16646] <= 8'h10 ;
			data[16647] <= 8'h10 ;
			data[16648] <= 8'h10 ;
			data[16649] <= 8'h10 ;
			data[16650] <= 8'h10 ;
			data[16651] <= 8'h10 ;
			data[16652] <= 8'h10 ;
			data[16653] <= 8'h10 ;
			data[16654] <= 8'h10 ;
			data[16655] <= 8'h10 ;
			data[16656] <= 8'h10 ;
			data[16657] <= 8'h10 ;
			data[16658] <= 8'h10 ;
			data[16659] <= 8'h10 ;
			data[16660] <= 8'h10 ;
			data[16661] <= 8'h10 ;
			data[16662] <= 8'h10 ;
			data[16663] <= 8'h10 ;
			data[16664] <= 8'h10 ;
			data[16665] <= 8'h10 ;
			data[16666] <= 8'h10 ;
			data[16667] <= 8'h10 ;
			data[16668] <= 8'h10 ;
			data[16669] <= 8'h10 ;
			data[16670] <= 8'h10 ;
			data[16671] <= 8'h10 ;
			data[16672] <= 8'h10 ;
			data[16673] <= 8'h10 ;
			data[16674] <= 8'h10 ;
			data[16675] <= 8'h10 ;
			data[16676] <= 8'h10 ;
			data[16677] <= 8'h10 ;
			data[16678] <= 8'h10 ;
			data[16679] <= 8'h10 ;
			data[16680] <= 8'h10 ;
			data[16681] <= 8'h10 ;
			data[16682] <= 8'h10 ;
			data[16683] <= 8'h10 ;
			data[16684] <= 8'h10 ;
			data[16685] <= 8'h10 ;
			data[16686] <= 8'h10 ;
			data[16687] <= 8'h10 ;
			data[16688] <= 8'h10 ;
			data[16689] <= 8'h10 ;
			data[16690] <= 8'h10 ;
			data[16691] <= 8'h10 ;
			data[16692] <= 8'h10 ;
			data[16693] <= 8'h10 ;
			data[16694] <= 8'h10 ;
			data[16695] <= 8'h10 ;
			data[16696] <= 8'h10 ;
			data[16697] <= 8'h10 ;
			data[16698] <= 8'h10 ;
			data[16699] <= 8'h10 ;
			data[16700] <= 8'h10 ;
			data[16701] <= 8'h10 ;
			data[16702] <= 8'h10 ;
			data[16703] <= 8'h10 ;
			data[16704] <= 8'h10 ;
			data[16705] <= 8'h10 ;
			data[16706] <= 8'h10 ;
			data[16707] <= 8'h10 ;
			data[16708] <= 8'h10 ;
			data[16709] <= 8'h10 ;
			data[16710] <= 8'h10 ;
			data[16711] <= 8'h10 ;
			data[16712] <= 8'h10 ;
			data[16713] <= 8'h10 ;
			data[16714] <= 8'h10 ;
			data[16715] <= 8'h10 ;
			data[16716] <= 8'h10 ;
			data[16717] <= 8'h10 ;
			data[16718] <= 8'h10 ;
			data[16719] <= 8'h10 ;
			data[16720] <= 8'h10 ;
			data[16721] <= 8'h10 ;
			data[16722] <= 8'h10 ;
			data[16723] <= 8'h10 ;
			data[16724] <= 8'h10 ;
			data[16725] <= 8'h10 ;
			data[16726] <= 8'h10 ;
			data[16727] <= 8'h10 ;
			data[16728] <= 8'h10 ;
			data[16729] <= 8'h10 ;
			data[16730] <= 8'h10 ;
			data[16731] <= 8'h10 ;
			data[16732] <= 8'h10 ;
			data[16733] <= 8'h10 ;
			data[16734] <= 8'h10 ;
			data[16735] <= 8'h10 ;
			data[16736] <= 8'h10 ;
			data[16737] <= 8'h10 ;
			data[16738] <= 8'h10 ;
			data[16739] <= 8'h10 ;
			data[16740] <= 8'h10 ;
			data[16741] <= 8'h10 ;
			data[16742] <= 8'h10 ;
			data[16743] <= 8'h10 ;
			data[16744] <= 8'h10 ;
			data[16745] <= 8'h10 ;
			data[16746] <= 8'h10 ;
			data[16747] <= 8'h10 ;
			data[16748] <= 8'h10 ;
			data[16749] <= 8'h10 ;
			data[16750] <= 8'h10 ;
			data[16751] <= 8'h10 ;
			data[16752] <= 8'h10 ;
			data[16753] <= 8'h10 ;
			data[16754] <= 8'h10 ;
			data[16755] <= 8'h10 ;
			data[16756] <= 8'h10 ;
			data[16757] <= 8'h10 ;
			data[16758] <= 8'h10 ;
			data[16759] <= 8'h10 ;
			data[16760] <= 8'h10 ;
			data[16761] <= 8'h10 ;
			data[16762] <= 8'h10 ;
			data[16763] <= 8'h10 ;
			data[16764] <= 8'h10 ;
			data[16765] <= 8'h10 ;
			data[16766] <= 8'h10 ;
			data[16767] <= 8'h10 ;
			data[16768] <= 8'h10 ;
			data[16769] <= 8'h10 ;
			data[16770] <= 8'h10 ;
			data[16771] <= 8'h10 ;
			data[16772] <= 8'h10 ;
			data[16773] <= 8'h10 ;
			data[16774] <= 8'h10 ;
			data[16775] <= 8'h10 ;
			data[16776] <= 8'h10 ;
			data[16777] <= 8'h10 ;
			data[16778] <= 8'h10 ;
			data[16779] <= 8'h10 ;
			data[16780] <= 8'h10 ;
			data[16781] <= 8'h10 ;
			data[16782] <= 8'h10 ;
			data[16783] <= 8'h10 ;
			data[16784] <= 8'h10 ;
			data[16785] <= 8'h10 ;
			data[16786] <= 8'h10 ;
			data[16787] <= 8'h10 ;
			data[16788] <= 8'h10 ;
			data[16789] <= 8'h10 ;
			data[16790] <= 8'h10 ;
			data[16791] <= 8'h10 ;
			data[16792] <= 8'h10 ;
			data[16793] <= 8'h10 ;
			data[16794] <= 8'h10 ;
			data[16795] <= 8'h10 ;
			data[16796] <= 8'h10 ;
			data[16797] <= 8'h10 ;
			data[16798] <= 8'h10 ;
			data[16799] <= 8'h10 ;
			data[16800] <= 8'h10 ;
			data[16801] <= 8'h10 ;
			data[16802] <= 8'h10 ;
			data[16803] <= 8'h10 ;
			data[16804] <= 8'h10 ;
			data[16805] <= 8'h10 ;
			data[16806] <= 8'h10 ;
			data[16807] <= 8'h10 ;
			data[16808] <= 8'h10 ;
			data[16809] <= 8'h10 ;
			data[16810] <= 8'h10 ;
			data[16811] <= 8'h10 ;
			data[16812] <= 8'h10 ;
			data[16813] <= 8'h10 ;
			data[16814] <= 8'h10 ;
			data[16815] <= 8'h10 ;
			data[16816] <= 8'h10 ;
			data[16817] <= 8'h10 ;
			data[16818] <= 8'h10 ;
			data[16819] <= 8'h10 ;
			data[16820] <= 8'h10 ;
			data[16821] <= 8'h10 ;
			data[16822] <= 8'h10 ;
			data[16823] <= 8'h10 ;
			data[16824] <= 8'h10 ;
			data[16825] <= 8'h10 ;
			data[16826] <= 8'h10 ;
			data[16827] <= 8'h10 ;
			data[16828] <= 8'h10 ;
			data[16829] <= 8'h10 ;
			data[16830] <= 8'h10 ;
			data[16831] <= 8'h10 ;
			data[16832] <= 8'h10 ;
			data[16833] <= 8'h10 ;
			data[16834] <= 8'h10 ;
			data[16835] <= 8'h10 ;
			data[16836] <= 8'h10 ;
			data[16837] <= 8'h10 ;
			data[16838] <= 8'h10 ;
			data[16839] <= 8'h10 ;
			data[16840] <= 8'h10 ;
			data[16841] <= 8'h10 ;
			data[16842] <= 8'h10 ;
			data[16843] <= 8'h10 ;
			data[16844] <= 8'h10 ;
			data[16845] <= 8'h10 ;
			data[16846] <= 8'h10 ;
			data[16847] <= 8'h10 ;
			data[16848] <= 8'h10 ;
			data[16849] <= 8'h10 ;
			data[16850] <= 8'h10 ;
			data[16851] <= 8'h10 ;
			data[16852] <= 8'h10 ;
			data[16853] <= 8'h10 ;
			data[16854] <= 8'h10 ;
			data[16855] <= 8'h10 ;
			data[16856] <= 8'h10 ;
			data[16857] <= 8'h10 ;
			data[16858] <= 8'h10 ;
			data[16859] <= 8'h10 ;
			data[16860] <= 8'h10 ;
			data[16861] <= 8'h10 ;
			data[16862] <= 8'h10 ;
			data[16863] <= 8'h10 ;
			data[16864] <= 8'h10 ;
			data[16865] <= 8'h10 ;
			data[16866] <= 8'h10 ;
			data[16867] <= 8'h10 ;
			data[16868] <= 8'h10 ;
			data[16869] <= 8'h10 ;
			data[16870] <= 8'h10 ;
			data[16871] <= 8'h10 ;
			data[16872] <= 8'h10 ;
			data[16873] <= 8'h10 ;
			data[16874] <= 8'h10 ;
			data[16875] <= 8'h10 ;
			data[16876] <= 8'h10 ;
			data[16877] <= 8'h10 ;
			data[16878] <= 8'h10 ;
			data[16879] <= 8'h10 ;
			data[16880] <= 8'h10 ;
			data[16881] <= 8'h10 ;
			data[16882] <= 8'h10 ;
			data[16883] <= 8'h10 ;
			data[16884] <= 8'h10 ;
			data[16885] <= 8'h10 ;
			data[16886] <= 8'h10 ;
			data[16887] <= 8'h10 ;
			data[16888] <= 8'h10 ;
			data[16889] <= 8'h10 ;
			data[16890] <= 8'h10 ;
			data[16891] <= 8'h10 ;
			data[16892] <= 8'h10 ;
			data[16893] <= 8'h10 ;
			data[16894] <= 8'h10 ;
			data[16895] <= 8'h10 ;
			data[16896] <= 8'h10 ;
			data[16897] <= 8'h10 ;
			data[16898] <= 8'h10 ;
			data[16899] <= 8'h10 ;
			data[16900] <= 8'h10 ;
			data[16901] <= 8'h10 ;
			data[16902] <= 8'h10 ;
			data[16903] <= 8'h10 ;
			data[16904] <= 8'h10 ;
			data[16905] <= 8'h10 ;
			data[16906] <= 8'h10 ;
			data[16907] <= 8'h10 ;
			data[16908] <= 8'h10 ;
			data[16909] <= 8'h10 ;
			data[16910] <= 8'h10 ;
			data[16911] <= 8'h10 ;
			data[16912] <= 8'h10 ;
			data[16913] <= 8'h10 ;
			data[16914] <= 8'h10 ;
			data[16915] <= 8'h10 ;
			data[16916] <= 8'h10 ;
			data[16917] <= 8'h10 ;
			data[16918] <= 8'h10 ;
			data[16919] <= 8'h10 ;
			data[16920] <= 8'h10 ;
			data[16921] <= 8'h10 ;
			data[16922] <= 8'h10 ;
			data[16923] <= 8'h10 ;
			data[16924] <= 8'h10 ;
			data[16925] <= 8'h10 ;
			data[16926] <= 8'h10 ;
			data[16927] <= 8'h10 ;
			data[16928] <= 8'h10 ;
			data[16929] <= 8'h10 ;
			data[16930] <= 8'h10 ;
			data[16931] <= 8'h10 ;
			data[16932] <= 8'h10 ;
			data[16933] <= 8'h10 ;
			data[16934] <= 8'h10 ;
			data[16935] <= 8'h10 ;
			data[16936] <= 8'h10 ;
			data[16937] <= 8'h10 ;
			data[16938] <= 8'h10 ;
			data[16939] <= 8'h10 ;
			data[16940] <= 8'h10 ;
			data[16941] <= 8'h10 ;
			data[16942] <= 8'h10 ;
			data[16943] <= 8'h10 ;
			data[16944] <= 8'h10 ;
			data[16945] <= 8'h10 ;
			data[16946] <= 8'h10 ;
			data[16947] <= 8'h10 ;
			data[16948] <= 8'h10 ;
			data[16949] <= 8'h10 ;
			data[16950] <= 8'h10 ;
			data[16951] <= 8'h10 ;
			data[16952] <= 8'h10 ;
			data[16953] <= 8'h10 ;
			data[16954] <= 8'h10 ;
			data[16955] <= 8'h10 ;
			data[16956] <= 8'h10 ;
			data[16957] <= 8'h10 ;
			data[16958] <= 8'h10 ;
			data[16959] <= 8'h10 ;
			data[16960] <= 8'h10 ;
			data[16961] <= 8'h10 ;
			data[16962] <= 8'h10 ;
			data[16963] <= 8'h10 ;
			data[16964] <= 8'h10 ;
			data[16965] <= 8'h10 ;
			data[16966] <= 8'h10 ;
			data[16967] <= 8'h10 ;
			data[16968] <= 8'h10 ;
			data[16969] <= 8'h10 ;
			data[16970] <= 8'h10 ;
			data[16971] <= 8'h10 ;
			data[16972] <= 8'h10 ;
			data[16973] <= 8'h10 ;
			data[16974] <= 8'h10 ;
			data[16975] <= 8'h10 ;
			data[16976] <= 8'h10 ;
			data[16977] <= 8'h10 ;
			data[16978] <= 8'h10 ;
			data[16979] <= 8'h10 ;
			data[16980] <= 8'h10 ;
			data[16981] <= 8'h10 ;
			data[16982] <= 8'h10 ;
			data[16983] <= 8'h10 ;
			data[16984] <= 8'h10 ;
			data[16985] <= 8'h10 ;
			data[16986] <= 8'h10 ;
			data[16987] <= 8'h10 ;
			data[16988] <= 8'h10 ;
			data[16989] <= 8'h10 ;
			data[16990] <= 8'h10 ;
			data[16991] <= 8'h10 ;
			data[16992] <= 8'h10 ;
			data[16993] <= 8'h10 ;
			data[16994] <= 8'h10 ;
			data[16995] <= 8'h10 ;
			data[16996] <= 8'h10 ;
			data[16997] <= 8'h10 ;
			data[16998] <= 8'h10 ;
			data[16999] <= 8'h10 ;
			data[17000] <= 8'h10 ;
			data[17001] <= 8'h10 ;
			data[17002] <= 8'h10 ;
			data[17003] <= 8'h10 ;
			data[17004] <= 8'h10 ;
			data[17005] <= 8'h10 ;
			data[17006] <= 8'h10 ;
			data[17007] <= 8'h10 ;
			data[17008] <= 8'h10 ;
			data[17009] <= 8'h10 ;
			data[17010] <= 8'h10 ;
			data[17011] <= 8'h10 ;
			data[17012] <= 8'h10 ;
			data[17013] <= 8'h10 ;
			data[17014] <= 8'h10 ;
			data[17015] <= 8'h10 ;
			data[17016] <= 8'h10 ;
			data[17017] <= 8'h10 ;
			data[17018] <= 8'h10 ;
			data[17019] <= 8'h10 ;
			data[17020] <= 8'h10 ;
			data[17021] <= 8'h10 ;
			data[17022] <= 8'h10 ;
			data[17023] <= 8'h10 ;
			data[17024] <= 8'h10 ;
			data[17025] <= 8'h10 ;
			data[17026] <= 8'h10 ;
			data[17027] <= 8'h10 ;
			data[17028] <= 8'h10 ;
			data[17029] <= 8'h10 ;
			data[17030] <= 8'h10 ;
			data[17031] <= 8'h10 ;
			data[17032] <= 8'h10 ;
			data[17033] <= 8'h10 ;
			data[17034] <= 8'h10 ;
			data[17035] <= 8'h10 ;
			data[17036] <= 8'h10 ;
			data[17037] <= 8'h10 ;
			data[17038] <= 8'h10 ;
			data[17039] <= 8'h10 ;
			data[17040] <= 8'h10 ;
			data[17041] <= 8'h10 ;
			data[17042] <= 8'h10 ;
			data[17043] <= 8'h10 ;
			data[17044] <= 8'h10 ;
			data[17045] <= 8'h10 ;
			data[17046] <= 8'h10 ;
			data[17047] <= 8'h10 ;
			data[17048] <= 8'h10 ;
			data[17049] <= 8'h10 ;
			data[17050] <= 8'h10 ;
			data[17051] <= 8'h10 ;
			data[17052] <= 8'h10 ;
			data[17053] <= 8'h10 ;
			data[17054] <= 8'h10 ;
			data[17055] <= 8'h10 ;
			data[17056] <= 8'h10 ;
			data[17057] <= 8'h10 ;
			data[17058] <= 8'h10 ;
			data[17059] <= 8'h10 ;
			data[17060] <= 8'h10 ;
			data[17061] <= 8'h10 ;
			data[17062] <= 8'h10 ;
			data[17063] <= 8'h10 ;
			data[17064] <= 8'h10 ;
			data[17065] <= 8'h10 ;
			data[17066] <= 8'h10 ;
			data[17067] <= 8'h10 ;
			data[17068] <= 8'h10 ;
			data[17069] <= 8'h10 ;
			data[17070] <= 8'h10 ;
			data[17071] <= 8'h10 ;
			data[17072] <= 8'h10 ;
			data[17073] <= 8'h10 ;
			data[17074] <= 8'h10 ;
			data[17075] <= 8'h10 ;
			data[17076] <= 8'h10 ;
			data[17077] <= 8'h10 ;
			data[17078] <= 8'h10 ;
			data[17079] <= 8'h10 ;
			data[17080] <= 8'h10 ;
			data[17081] <= 8'h10 ;
			data[17082] <= 8'h10 ;
			data[17083] <= 8'h10 ;
			data[17084] <= 8'h10 ;
			data[17085] <= 8'h10 ;
			data[17086] <= 8'h10 ;
			data[17087] <= 8'h10 ;
			data[17088] <= 8'h10 ;
			data[17089] <= 8'h10 ;
			data[17090] <= 8'h10 ;
			data[17091] <= 8'h10 ;
			data[17092] <= 8'h10 ;
			data[17093] <= 8'h10 ;
			data[17094] <= 8'h10 ;
			data[17095] <= 8'h10 ;
			data[17096] <= 8'h10 ;
			data[17097] <= 8'h10 ;
			data[17098] <= 8'h10 ;
			data[17099] <= 8'h10 ;
			data[17100] <= 8'h10 ;
			data[17101] <= 8'h10 ;
			data[17102] <= 8'h10 ;
			data[17103] <= 8'h10 ;
			data[17104] <= 8'h10 ;
			data[17105] <= 8'h10 ;
			data[17106] <= 8'h10 ;
			data[17107] <= 8'h10 ;
			data[17108] <= 8'h10 ;
			data[17109] <= 8'h10 ;
			data[17110] <= 8'h10 ;
			data[17111] <= 8'h10 ;
			data[17112] <= 8'h10 ;
			data[17113] <= 8'h10 ;
			data[17114] <= 8'h10 ;
			data[17115] <= 8'h10 ;
			data[17116] <= 8'h10 ;
			data[17117] <= 8'h10 ;
			data[17118] <= 8'h10 ;
			data[17119] <= 8'h10 ;
			data[17120] <= 8'h10 ;
			data[17121] <= 8'h10 ;
			data[17122] <= 8'h10 ;
			data[17123] <= 8'h10 ;
			data[17124] <= 8'h10 ;
			data[17125] <= 8'h10 ;
			data[17126] <= 8'h10 ;
			data[17127] <= 8'h10 ;
			data[17128] <= 8'h10 ;
			data[17129] <= 8'h10 ;
			data[17130] <= 8'h10 ;
			data[17131] <= 8'h10 ;
			data[17132] <= 8'h10 ;
			data[17133] <= 8'h10 ;
			data[17134] <= 8'h10 ;
			data[17135] <= 8'h10 ;
			data[17136] <= 8'h10 ;
			data[17137] <= 8'h10 ;
			data[17138] <= 8'h10 ;
			data[17139] <= 8'h10 ;
			data[17140] <= 8'h10 ;
			data[17141] <= 8'h10 ;
			data[17142] <= 8'h10 ;
			data[17143] <= 8'h10 ;
			data[17144] <= 8'h10 ;
			data[17145] <= 8'h10 ;
			data[17146] <= 8'h10 ;
			data[17147] <= 8'h10 ;
			data[17148] <= 8'h10 ;
			data[17149] <= 8'h10 ;
			data[17150] <= 8'h10 ;
			data[17151] <= 8'h10 ;
			data[17152] <= 8'h10 ;
			data[17153] <= 8'h10 ;
			data[17154] <= 8'h10 ;
			data[17155] <= 8'h10 ;
			data[17156] <= 8'h10 ;
			data[17157] <= 8'h10 ;
			data[17158] <= 8'h10 ;
			data[17159] <= 8'h10 ;
			data[17160] <= 8'h10 ;
			data[17161] <= 8'h10 ;
			data[17162] <= 8'h10 ;
			data[17163] <= 8'h10 ;
			data[17164] <= 8'h10 ;
			data[17165] <= 8'h10 ;
			data[17166] <= 8'h10 ;
			data[17167] <= 8'h10 ;
			data[17168] <= 8'h10 ;
			data[17169] <= 8'h10 ;
			data[17170] <= 8'h10 ;
			data[17171] <= 8'h10 ;
			data[17172] <= 8'h10 ;
			data[17173] <= 8'h10 ;
			data[17174] <= 8'h10 ;
			data[17175] <= 8'h10 ;
			data[17176] <= 8'h10 ;
			data[17177] <= 8'h10 ;
			data[17178] <= 8'h10 ;
			data[17179] <= 8'h10 ;
			data[17180] <= 8'h10 ;
			data[17181] <= 8'h10 ;
			data[17182] <= 8'h10 ;
			data[17183] <= 8'h10 ;
			data[17184] <= 8'h10 ;
			data[17185] <= 8'h10 ;
			data[17186] <= 8'h10 ;
			data[17187] <= 8'h10 ;
			data[17188] <= 8'h10 ;
			data[17189] <= 8'h10 ;
			data[17190] <= 8'h10 ;
			data[17191] <= 8'h10 ;
			data[17192] <= 8'h10 ;
			data[17193] <= 8'h10 ;
			data[17194] <= 8'h10 ;
			data[17195] <= 8'h10 ;
			data[17196] <= 8'h10 ;
			data[17197] <= 8'h10 ;
			data[17198] <= 8'h10 ;
			data[17199] <= 8'h10 ;
			data[17200] <= 8'h10 ;
			data[17201] <= 8'h10 ;
			data[17202] <= 8'h10 ;
			data[17203] <= 8'h10 ;
			data[17204] <= 8'h10 ;
			data[17205] <= 8'h10 ;
			data[17206] <= 8'h10 ;
			data[17207] <= 8'h10 ;
			data[17208] <= 8'h10 ;
			data[17209] <= 8'h10 ;
			data[17210] <= 8'h10 ;
			data[17211] <= 8'h10 ;
			data[17212] <= 8'h10 ;
			data[17213] <= 8'h10 ;
			data[17214] <= 8'h10 ;
			data[17215] <= 8'h10 ;
			data[17216] <= 8'h10 ;
			data[17217] <= 8'h10 ;
			data[17218] <= 8'h10 ;
			data[17219] <= 8'h10 ;
			data[17220] <= 8'h10 ;
			data[17221] <= 8'h10 ;
			data[17222] <= 8'h10 ;
			data[17223] <= 8'h10 ;
			data[17224] <= 8'h10 ;
			data[17225] <= 8'h10 ;
			data[17226] <= 8'h10 ;
			data[17227] <= 8'h10 ;
			data[17228] <= 8'h10 ;
			data[17229] <= 8'h10 ;
			data[17230] <= 8'h10 ;
			data[17231] <= 8'h10 ;
			data[17232] <= 8'h10 ;
			data[17233] <= 8'h10 ;
			data[17234] <= 8'h10 ;
			data[17235] <= 8'h10 ;
			data[17236] <= 8'h10 ;
			data[17237] <= 8'h10 ;
			data[17238] <= 8'h10 ;
			data[17239] <= 8'h10 ;
			data[17240] <= 8'h10 ;
			data[17241] <= 8'h10 ;
			data[17242] <= 8'h10 ;
			data[17243] <= 8'h10 ;
			data[17244] <= 8'h10 ;
			data[17245] <= 8'h10 ;
			data[17246] <= 8'h10 ;
			data[17247] <= 8'h10 ;
			data[17248] <= 8'h10 ;
			data[17249] <= 8'h10 ;
			data[17250] <= 8'h10 ;
			data[17251] <= 8'h10 ;
			data[17252] <= 8'h10 ;
			data[17253] <= 8'h10 ;
			data[17254] <= 8'h10 ;
			data[17255] <= 8'h10 ;
			data[17256] <= 8'h10 ;
			data[17257] <= 8'h10 ;
			data[17258] <= 8'h10 ;
			data[17259] <= 8'h10 ;
			data[17260] <= 8'h10 ;
			data[17261] <= 8'h10 ;
			data[17262] <= 8'h10 ;
			data[17263] <= 8'h10 ;
			data[17264] <= 8'h10 ;
			data[17265] <= 8'h10 ;
			data[17266] <= 8'h10 ;
			data[17267] <= 8'h10 ;
			data[17268] <= 8'h10 ;
			data[17269] <= 8'h10 ;
			data[17270] <= 8'h10 ;
			data[17271] <= 8'h10 ;
			data[17272] <= 8'h10 ;
			data[17273] <= 8'h10 ;
			data[17274] <= 8'h10 ;
			data[17275] <= 8'h10 ;
			data[17276] <= 8'h10 ;
			data[17277] <= 8'h10 ;
			data[17278] <= 8'h10 ;
			data[17279] <= 8'h10 ;
			data[17280] <= 8'h10 ;
			data[17281] <= 8'h10 ;
			data[17282] <= 8'h10 ;
			data[17283] <= 8'h10 ;
			data[17284] <= 8'h10 ;
			data[17285] <= 8'h10 ;
			data[17286] <= 8'h10 ;
			data[17287] <= 8'h10 ;
			data[17288] <= 8'h10 ;
			data[17289] <= 8'h10 ;
			data[17290] <= 8'h10 ;
			data[17291] <= 8'h10 ;
			data[17292] <= 8'h10 ;
			data[17293] <= 8'h10 ;
			data[17294] <= 8'h10 ;
			data[17295] <= 8'h10 ;
			data[17296] <= 8'h10 ;
			data[17297] <= 8'h10 ;
			data[17298] <= 8'h10 ;
			data[17299] <= 8'h10 ;
			data[17300] <= 8'h10 ;
			data[17301] <= 8'h10 ;
			data[17302] <= 8'h10 ;
			data[17303] <= 8'h10 ;
			data[17304] <= 8'h10 ;
			data[17305] <= 8'h10 ;
			data[17306] <= 8'h10 ;
			data[17307] <= 8'h10 ;
			data[17308] <= 8'h10 ;
			data[17309] <= 8'h10 ;
			data[17310] <= 8'h10 ;
			data[17311] <= 8'h10 ;
			data[17312] <= 8'h10 ;
			data[17313] <= 8'h10 ;
			data[17314] <= 8'h10 ;
			data[17315] <= 8'h10 ;
			data[17316] <= 8'h10 ;
			data[17317] <= 8'h10 ;
			data[17318] <= 8'h10 ;
			data[17319] <= 8'h10 ;
			data[17320] <= 8'h10 ;
			data[17321] <= 8'h10 ;
			data[17322] <= 8'h10 ;
			data[17323] <= 8'h10 ;
			data[17324] <= 8'h10 ;
			data[17325] <= 8'h10 ;
			data[17326] <= 8'h10 ;
			data[17327] <= 8'h10 ;
			data[17328] <= 8'h10 ;
			data[17329] <= 8'h10 ;
			data[17330] <= 8'h10 ;
			data[17331] <= 8'h10 ;
			data[17332] <= 8'h10 ;
			data[17333] <= 8'h10 ;
			data[17334] <= 8'h10 ;
			data[17335] <= 8'h10 ;
			data[17336] <= 8'h10 ;
			data[17337] <= 8'h10 ;
			data[17338] <= 8'h10 ;
			data[17339] <= 8'h10 ;
			data[17340] <= 8'h10 ;
			data[17341] <= 8'h10 ;
			data[17342] <= 8'h10 ;
			data[17343] <= 8'h10 ;
			data[17344] <= 8'h10 ;
			data[17345] <= 8'h10 ;
			data[17346] <= 8'h10 ;
			data[17347] <= 8'h10 ;
			data[17348] <= 8'h10 ;
			data[17349] <= 8'h10 ;
			data[17350] <= 8'h10 ;
			data[17351] <= 8'h10 ;
			data[17352] <= 8'h10 ;
			data[17353] <= 8'h10 ;
			data[17354] <= 8'h10 ;
			data[17355] <= 8'h10 ;
			data[17356] <= 8'h10 ;
			data[17357] <= 8'h10 ;
			data[17358] <= 8'h10 ;
			data[17359] <= 8'h10 ;
			data[17360] <= 8'h10 ;
			data[17361] <= 8'h10 ;
			data[17362] <= 8'h10 ;
			data[17363] <= 8'h10 ;
			data[17364] <= 8'h10 ;
			data[17365] <= 8'h10 ;
			data[17366] <= 8'h10 ;
			data[17367] <= 8'h10 ;
			data[17368] <= 8'h10 ;
			data[17369] <= 8'h10 ;
			data[17370] <= 8'h10 ;
			data[17371] <= 8'h10 ;
			data[17372] <= 8'h10 ;
			data[17373] <= 8'h10 ;
			data[17374] <= 8'h10 ;
			data[17375] <= 8'h10 ;
			data[17376] <= 8'h10 ;
			data[17377] <= 8'h10 ;
			data[17378] <= 8'h10 ;
			data[17379] <= 8'h10 ;
			data[17380] <= 8'h10 ;
			data[17381] <= 8'h10 ;
			data[17382] <= 8'h10 ;
			data[17383] <= 8'h10 ;
			data[17384] <= 8'h10 ;
			data[17385] <= 8'h10 ;
			data[17386] <= 8'h10 ;
			data[17387] <= 8'h10 ;
			data[17388] <= 8'h10 ;
			data[17389] <= 8'h10 ;
			data[17390] <= 8'h10 ;
			data[17391] <= 8'h10 ;
			data[17392] <= 8'h10 ;
			data[17393] <= 8'h10 ;
			data[17394] <= 8'h10 ;
			data[17395] <= 8'h10 ;
			data[17396] <= 8'h10 ;
			data[17397] <= 8'h10 ;
			data[17398] <= 8'h10 ;
			data[17399] <= 8'h10 ;
			data[17400] <= 8'h10 ;
			data[17401] <= 8'h10 ;
			data[17402] <= 8'h10 ;
			data[17403] <= 8'h10 ;
			data[17404] <= 8'h10 ;
			data[17405] <= 8'h10 ;
			data[17406] <= 8'h10 ;
			data[17407] <= 8'h10 ;
			data[17408] <= 8'h10 ;
			data[17409] <= 8'h10 ;
			data[17410] <= 8'h10 ;
			data[17411] <= 8'h10 ;
			data[17412] <= 8'h10 ;
			data[17413] <= 8'h10 ;
			data[17414] <= 8'h10 ;
			data[17415] <= 8'h10 ;
			data[17416] <= 8'h10 ;
			data[17417] <= 8'h10 ;
			data[17418] <= 8'h10 ;
			data[17419] <= 8'h10 ;
			data[17420] <= 8'h10 ;
			data[17421] <= 8'h10 ;
			data[17422] <= 8'h10 ;
			data[17423] <= 8'h10 ;
			data[17424] <= 8'h10 ;
			data[17425] <= 8'h10 ;
			data[17426] <= 8'h10 ;
			data[17427] <= 8'h10 ;
			data[17428] <= 8'h10 ;
			data[17429] <= 8'h10 ;
			data[17430] <= 8'h10 ;
			data[17431] <= 8'h10 ;
			data[17432] <= 8'h10 ;
			data[17433] <= 8'h10 ;
			data[17434] <= 8'h10 ;
			data[17435] <= 8'h10 ;
			data[17436] <= 8'h10 ;
			data[17437] <= 8'h10 ;
			data[17438] <= 8'h10 ;
			data[17439] <= 8'h10 ;
			data[17440] <= 8'h10 ;
			data[17441] <= 8'h10 ;
			data[17442] <= 8'h10 ;
			data[17443] <= 8'h10 ;
			data[17444] <= 8'h10 ;
			data[17445] <= 8'h10 ;
			data[17446] <= 8'h10 ;
			data[17447] <= 8'h10 ;
			data[17448] <= 8'h10 ;
			data[17449] <= 8'h10 ;
			data[17450] <= 8'h10 ;
			data[17451] <= 8'h10 ;
			data[17452] <= 8'h10 ;
			data[17453] <= 8'h10 ;
			data[17454] <= 8'h10 ;
			data[17455] <= 8'h10 ;
			data[17456] <= 8'h10 ;
			data[17457] <= 8'h10 ;
			data[17458] <= 8'h10 ;
			data[17459] <= 8'h10 ;
			data[17460] <= 8'h10 ;
			data[17461] <= 8'h10 ;
			data[17462] <= 8'h10 ;
			data[17463] <= 8'h10 ;
			data[17464] <= 8'h10 ;
			data[17465] <= 8'h10 ;
			data[17466] <= 8'h10 ;
			data[17467] <= 8'h10 ;
			data[17468] <= 8'h10 ;
			data[17469] <= 8'h10 ;
			data[17470] <= 8'h10 ;
			data[17471] <= 8'h10 ;
			data[17472] <= 8'h10 ;
			data[17473] <= 8'h10 ;
			data[17474] <= 8'h10 ;
			data[17475] <= 8'h10 ;
			data[17476] <= 8'h10 ;
			data[17477] <= 8'h10 ;
			data[17478] <= 8'h10 ;
			data[17479] <= 8'h10 ;
			data[17480] <= 8'h10 ;
			data[17481] <= 8'h10 ;
			data[17482] <= 8'h10 ;
			data[17483] <= 8'h10 ;
			data[17484] <= 8'h10 ;
			data[17485] <= 8'h10 ;
			data[17486] <= 8'h10 ;
			data[17487] <= 8'h10 ;
			data[17488] <= 8'h10 ;
			data[17489] <= 8'h10 ;
			data[17490] <= 8'h10 ;
			data[17491] <= 8'h10 ;
			data[17492] <= 8'h10 ;
			data[17493] <= 8'h10 ;
			data[17494] <= 8'h10 ;
			data[17495] <= 8'h10 ;
			data[17496] <= 8'h10 ;
			data[17497] <= 8'h10 ;
			data[17498] <= 8'h10 ;
			data[17499] <= 8'h10 ;
			data[17500] <= 8'h10 ;
			data[17501] <= 8'h10 ;
			data[17502] <= 8'h10 ;
			data[17503] <= 8'h10 ;
			data[17504] <= 8'h10 ;
			data[17505] <= 8'h10 ;
			data[17506] <= 8'h10 ;
			data[17507] <= 8'h10 ;
			data[17508] <= 8'h10 ;
			data[17509] <= 8'h10 ;
			data[17510] <= 8'h10 ;
			data[17511] <= 8'h10 ;
			data[17512] <= 8'h10 ;
			data[17513] <= 8'h10 ;
			data[17514] <= 8'h10 ;
			data[17515] <= 8'h10 ;
			data[17516] <= 8'h10 ;
			data[17517] <= 8'h10 ;
			data[17518] <= 8'h10 ;
			data[17519] <= 8'h10 ;
			data[17520] <= 8'h10 ;
			data[17521] <= 8'h10 ;
			data[17522] <= 8'h10 ;
			data[17523] <= 8'h10 ;
			data[17524] <= 8'h10 ;
			data[17525] <= 8'h10 ;
			data[17526] <= 8'h10 ;
			data[17527] <= 8'h10 ;
			data[17528] <= 8'h10 ;
			data[17529] <= 8'h10 ;
			data[17530] <= 8'h10 ;
			data[17531] <= 8'h10 ;
			data[17532] <= 8'h10 ;
			data[17533] <= 8'h10 ;
			data[17534] <= 8'h10 ;
			data[17535] <= 8'h10 ;
			data[17536] <= 8'h10 ;
			data[17537] <= 8'h10 ;
			data[17538] <= 8'h10 ;
			data[17539] <= 8'h10 ;
			data[17540] <= 8'h10 ;
			data[17541] <= 8'h10 ;
			data[17542] <= 8'h10 ;
			data[17543] <= 8'h10 ;
			data[17544] <= 8'h10 ;
			data[17545] <= 8'h10 ;
			data[17546] <= 8'h10 ;
			data[17547] <= 8'h10 ;
			data[17548] <= 8'h10 ;
			data[17549] <= 8'h10 ;
			data[17550] <= 8'h10 ;
			data[17551] <= 8'h10 ;
			data[17552] <= 8'h10 ;
			data[17553] <= 8'h10 ;
			data[17554] <= 8'h10 ;
			data[17555] <= 8'h10 ;
			data[17556] <= 8'h10 ;
			data[17557] <= 8'h10 ;
			data[17558] <= 8'h10 ;
			data[17559] <= 8'h10 ;
			data[17560] <= 8'h10 ;
			data[17561] <= 8'h10 ;
			data[17562] <= 8'h10 ;
			data[17563] <= 8'h10 ;
			data[17564] <= 8'h10 ;
			data[17565] <= 8'h10 ;
			data[17566] <= 8'h10 ;
			data[17567] <= 8'h10 ;
			data[17568] <= 8'h10 ;
			data[17569] <= 8'h10 ;
			data[17570] <= 8'h10 ;
			data[17571] <= 8'h10 ;
			data[17572] <= 8'h10 ;
			data[17573] <= 8'h10 ;
			data[17574] <= 8'h10 ;
			data[17575] <= 8'h10 ;
			data[17576] <= 8'h10 ;
			data[17577] <= 8'h10 ;
			data[17578] <= 8'h10 ;
			data[17579] <= 8'h10 ;
			data[17580] <= 8'h10 ;
			data[17581] <= 8'h10 ;
			data[17582] <= 8'h10 ;
			data[17583] <= 8'h10 ;
			data[17584] <= 8'h10 ;
			data[17585] <= 8'h10 ;
			data[17586] <= 8'h10 ;
			data[17587] <= 8'h10 ;
			data[17588] <= 8'h10 ;
			data[17589] <= 8'h10 ;
			data[17590] <= 8'h10 ;
			data[17591] <= 8'h10 ;
			data[17592] <= 8'h10 ;
			data[17593] <= 8'h10 ;
			data[17594] <= 8'h10 ;
			data[17595] <= 8'h10 ;
			data[17596] <= 8'h10 ;
			data[17597] <= 8'h10 ;
			data[17598] <= 8'h10 ;
			data[17599] <= 8'h10 ;
			data[17600] <= 8'h10 ;
			data[17601] <= 8'h10 ;
			data[17602] <= 8'h10 ;
			data[17603] <= 8'h10 ;
			data[17604] <= 8'h10 ;
			data[17605] <= 8'h10 ;
			data[17606] <= 8'h10 ;
			data[17607] <= 8'h10 ;
			data[17608] <= 8'h10 ;
			data[17609] <= 8'h10 ;
			data[17610] <= 8'h10 ;
			data[17611] <= 8'h10 ;
			data[17612] <= 8'h10 ;
			data[17613] <= 8'h10 ;
			data[17614] <= 8'h10 ;
			data[17615] <= 8'h10 ;
			data[17616] <= 8'h10 ;
			data[17617] <= 8'h10 ;
			data[17618] <= 8'h10 ;
			data[17619] <= 8'h10 ;
			data[17620] <= 8'h10 ;
			data[17621] <= 8'h10 ;
			data[17622] <= 8'h10 ;
			data[17623] <= 8'h10 ;
			data[17624] <= 8'h10 ;
			data[17625] <= 8'h10 ;
			data[17626] <= 8'h10 ;
			data[17627] <= 8'h10 ;
			data[17628] <= 8'h10 ;
			data[17629] <= 8'h10 ;
			data[17630] <= 8'h10 ;
			data[17631] <= 8'h10 ;
			data[17632] <= 8'h10 ;
			data[17633] <= 8'h10 ;
			data[17634] <= 8'h10 ;
			data[17635] <= 8'h10 ;
			data[17636] <= 8'h10 ;
			data[17637] <= 8'h10 ;
			data[17638] <= 8'h10 ;
			data[17639] <= 8'h10 ;
			data[17640] <= 8'h10 ;
			data[17641] <= 8'h10 ;
			data[17642] <= 8'h10 ;
			data[17643] <= 8'h10 ;
			data[17644] <= 8'h10 ;
			data[17645] <= 8'h10 ;
			data[17646] <= 8'h10 ;
			data[17647] <= 8'h10 ;
			data[17648] <= 8'h10 ;
			data[17649] <= 8'h10 ;
			data[17650] <= 8'h10 ;
			data[17651] <= 8'h10 ;
			data[17652] <= 8'h10 ;
			data[17653] <= 8'h10 ;
			data[17654] <= 8'h10 ;
			data[17655] <= 8'h10 ;
			data[17656] <= 8'h10 ;
			data[17657] <= 8'h10 ;
			data[17658] <= 8'h10 ;
			data[17659] <= 8'h10 ;
			data[17660] <= 8'h10 ;
			data[17661] <= 8'h10 ;
			data[17662] <= 8'h10 ;
			data[17663] <= 8'h10 ;
			data[17664] <= 8'h10 ;
			data[17665] <= 8'h10 ;
			data[17666] <= 8'h10 ;
			data[17667] <= 8'h10 ;
			data[17668] <= 8'h10 ;
			data[17669] <= 8'h10 ;
			data[17670] <= 8'h10 ;
			data[17671] <= 8'h10 ;
			data[17672] <= 8'h10 ;
			data[17673] <= 8'h10 ;
			data[17674] <= 8'h10 ;
			data[17675] <= 8'h10 ;
			data[17676] <= 8'h10 ;
			data[17677] <= 8'h10 ;
			data[17678] <= 8'h10 ;
			data[17679] <= 8'h10 ;
			data[17680] <= 8'h10 ;
			data[17681] <= 8'h10 ;
			data[17682] <= 8'h10 ;
			data[17683] <= 8'h10 ;
			data[17684] <= 8'h10 ;
			data[17685] <= 8'h10 ;
			data[17686] <= 8'h10 ;
			data[17687] <= 8'h10 ;
			data[17688] <= 8'h10 ;
			data[17689] <= 8'h10 ;
			data[17690] <= 8'h10 ;
			data[17691] <= 8'h10 ;
			data[17692] <= 8'h10 ;
			data[17693] <= 8'h10 ;
			data[17694] <= 8'h10 ;
			data[17695] <= 8'h10 ;
			data[17696] <= 8'h10 ;
			data[17697] <= 8'h10 ;
			data[17698] <= 8'h10 ;
			data[17699] <= 8'h10 ;
			data[17700] <= 8'h10 ;
			data[17701] <= 8'h10 ;
			data[17702] <= 8'h10 ;
			data[17703] <= 8'h10 ;
			data[17704] <= 8'h10 ;
			data[17705] <= 8'h10 ;
			data[17706] <= 8'h10 ;
			data[17707] <= 8'h10 ;
			data[17708] <= 8'h10 ;
			data[17709] <= 8'h10 ;
			data[17710] <= 8'h10 ;
			data[17711] <= 8'h10 ;
			data[17712] <= 8'h10 ;
			data[17713] <= 8'h10 ;
			data[17714] <= 8'h10 ;
			data[17715] <= 8'h10 ;
			data[17716] <= 8'h10 ;
			data[17717] <= 8'h10 ;
			data[17718] <= 8'h10 ;
			data[17719] <= 8'h10 ;
			data[17720] <= 8'h10 ;
			data[17721] <= 8'h10 ;
			data[17722] <= 8'h10 ;
			data[17723] <= 8'h10 ;
			data[17724] <= 8'h10 ;
			data[17725] <= 8'h10 ;
			data[17726] <= 8'h10 ;
			data[17727] <= 8'h10 ;
			data[17728] <= 8'h10 ;
			data[17729] <= 8'h10 ;
			data[17730] <= 8'h10 ;
			data[17731] <= 8'h10 ;
			data[17732] <= 8'h10 ;
			data[17733] <= 8'h10 ;
			data[17734] <= 8'h10 ;
			data[17735] <= 8'h10 ;
			data[17736] <= 8'h10 ;
			data[17737] <= 8'h10 ;
			data[17738] <= 8'h10 ;
			data[17739] <= 8'h10 ;
			data[17740] <= 8'h10 ;
			data[17741] <= 8'h10 ;
			data[17742] <= 8'h10 ;
			data[17743] <= 8'h10 ;
			data[17744] <= 8'h10 ;
			data[17745] <= 8'h10 ;
			data[17746] <= 8'h10 ;
			data[17747] <= 8'h10 ;
			data[17748] <= 8'h10 ;
			data[17749] <= 8'h10 ;
			data[17750] <= 8'h10 ;
			data[17751] <= 8'h10 ;
			data[17752] <= 8'h10 ;
			data[17753] <= 8'h10 ;
			data[17754] <= 8'h10 ;
			data[17755] <= 8'h10 ;
			data[17756] <= 8'h10 ;
			data[17757] <= 8'h10 ;
			data[17758] <= 8'h10 ;
			data[17759] <= 8'h10 ;
			data[17760] <= 8'h10 ;
			data[17761] <= 8'h10 ;
			data[17762] <= 8'h10 ;
			data[17763] <= 8'h10 ;
			data[17764] <= 8'h10 ;
			data[17765] <= 8'h10 ;
			data[17766] <= 8'h10 ;
			data[17767] <= 8'h10 ;
			data[17768] <= 8'h10 ;
			data[17769] <= 8'h10 ;
			data[17770] <= 8'h10 ;
			data[17771] <= 8'h10 ;
			data[17772] <= 8'h10 ;
			data[17773] <= 8'h10 ;
			data[17774] <= 8'h10 ;
			data[17775] <= 8'h10 ;
			data[17776] <= 8'h10 ;
			data[17777] <= 8'h10 ;
			data[17778] <= 8'h10 ;
			data[17779] <= 8'h10 ;
			data[17780] <= 8'h10 ;
			data[17781] <= 8'h10 ;
			data[17782] <= 8'h10 ;
			data[17783] <= 8'h10 ;
			data[17784] <= 8'h10 ;
			data[17785] <= 8'h10 ;
			data[17786] <= 8'h10 ;
			data[17787] <= 8'h10 ;
			data[17788] <= 8'h10 ;
			data[17789] <= 8'h10 ;
			data[17790] <= 8'h10 ;
			data[17791] <= 8'h10 ;
			data[17792] <= 8'h10 ;
			data[17793] <= 8'h10 ;
			data[17794] <= 8'h10 ;
			data[17795] <= 8'h10 ;
			data[17796] <= 8'h10 ;
			data[17797] <= 8'h10 ;
			data[17798] <= 8'h10 ;
			data[17799] <= 8'h10 ;
			data[17800] <= 8'h10 ;
			data[17801] <= 8'h10 ;
			data[17802] <= 8'h10 ;
			data[17803] <= 8'h10 ;
			data[17804] <= 8'h10 ;
			data[17805] <= 8'h10 ;
			data[17806] <= 8'h10 ;
			data[17807] <= 8'h10 ;
			data[17808] <= 8'h10 ;
			data[17809] <= 8'h10 ;
			data[17810] <= 8'h10 ;
			data[17811] <= 8'h10 ;
			data[17812] <= 8'h10 ;
			data[17813] <= 8'h10 ;
			data[17814] <= 8'h10 ;
			data[17815] <= 8'h10 ;
			data[17816] <= 8'h10 ;
			data[17817] <= 8'h10 ;
			data[17818] <= 8'h10 ;
			data[17819] <= 8'h10 ;
			data[17820] <= 8'h10 ;
			data[17821] <= 8'h10 ;
			data[17822] <= 8'h10 ;
			data[17823] <= 8'h10 ;
			data[17824] <= 8'h10 ;
			data[17825] <= 8'h10 ;
			data[17826] <= 8'h10 ;
			data[17827] <= 8'h10 ;
			data[17828] <= 8'h10 ;
			data[17829] <= 8'h10 ;
			data[17830] <= 8'h10 ;
			data[17831] <= 8'h10 ;
			data[17832] <= 8'h10 ;
			data[17833] <= 8'h10 ;
			data[17834] <= 8'h10 ;
			data[17835] <= 8'h10 ;
			data[17836] <= 8'h10 ;
			data[17837] <= 8'h10 ;
			data[17838] <= 8'h10 ;
			data[17839] <= 8'h10 ;
			data[17840] <= 8'h10 ;
			data[17841] <= 8'h10 ;
			data[17842] <= 8'h10 ;
			data[17843] <= 8'h10 ;
			data[17844] <= 8'h10 ;
			data[17845] <= 8'h10 ;
			data[17846] <= 8'h10 ;
			data[17847] <= 8'h10 ;
			data[17848] <= 8'h10 ;
			data[17849] <= 8'h10 ;
			data[17850] <= 8'h10 ;
			data[17851] <= 8'h10 ;
			data[17852] <= 8'h10 ;
			data[17853] <= 8'h10 ;
			data[17854] <= 8'h10 ;
			data[17855] <= 8'h10 ;
			data[17856] <= 8'h10 ;
			data[17857] <= 8'h10 ;
			data[17858] <= 8'h10 ;
			data[17859] <= 8'h10 ;
			data[17860] <= 8'h10 ;
			data[17861] <= 8'h10 ;
			data[17862] <= 8'h10 ;
			data[17863] <= 8'h10 ;
			data[17864] <= 8'h10 ;
			data[17865] <= 8'h10 ;
			data[17866] <= 8'h10 ;
			data[17867] <= 8'h10 ;
			data[17868] <= 8'h10 ;
			data[17869] <= 8'h10 ;
			data[17870] <= 8'h10 ;
			data[17871] <= 8'h10 ;
			data[17872] <= 8'h10 ;
			data[17873] <= 8'h10 ;
			data[17874] <= 8'h10 ;
			data[17875] <= 8'h10 ;
			data[17876] <= 8'h10 ;
			data[17877] <= 8'h10 ;
			data[17878] <= 8'h10 ;
			data[17879] <= 8'h10 ;
			data[17880] <= 8'h10 ;
			data[17881] <= 8'h10 ;
			data[17882] <= 8'h10 ;
			data[17883] <= 8'h10 ;
			data[17884] <= 8'h10 ;
			data[17885] <= 8'h10 ;
			data[17886] <= 8'h10 ;
			data[17887] <= 8'h10 ;
			data[17888] <= 8'h10 ;
			data[17889] <= 8'h10 ;
			data[17890] <= 8'h10 ;
			data[17891] <= 8'h10 ;
			data[17892] <= 8'h10 ;
			data[17893] <= 8'h10 ;
			data[17894] <= 8'h10 ;
			data[17895] <= 8'h10 ;
			data[17896] <= 8'h10 ;
			data[17897] <= 8'h10 ;
			data[17898] <= 8'h10 ;
			data[17899] <= 8'h10 ;
			data[17900] <= 8'h10 ;
			data[17901] <= 8'h10 ;
			data[17902] <= 8'h10 ;
			data[17903] <= 8'h10 ;
			data[17904] <= 8'h10 ;
			data[17905] <= 8'h10 ;
			data[17906] <= 8'h10 ;
			data[17907] <= 8'h10 ;
			data[17908] <= 8'h10 ;
			data[17909] <= 8'h10 ;
			data[17910] <= 8'h10 ;
			data[17911] <= 8'h10 ;
			data[17912] <= 8'h10 ;
			data[17913] <= 8'h10 ;
			data[17914] <= 8'h10 ;
			data[17915] <= 8'h10 ;
			data[17916] <= 8'h10 ;
			data[17917] <= 8'h10 ;
			data[17918] <= 8'h10 ;
			data[17919] <= 8'h10 ;
			data[17920] <= 8'h10 ;
			data[17921] <= 8'h10 ;
			data[17922] <= 8'h10 ;
			data[17923] <= 8'h10 ;
			data[17924] <= 8'h10 ;
			data[17925] <= 8'h10 ;
			data[17926] <= 8'h10 ;
			data[17927] <= 8'h10 ;
			data[17928] <= 8'h10 ;
			data[17929] <= 8'h10 ;
			data[17930] <= 8'h10 ;
			data[17931] <= 8'h10 ;
			data[17932] <= 8'h10 ;
			data[17933] <= 8'h10 ;
			data[17934] <= 8'h10 ;
			data[17935] <= 8'h10 ;
			data[17936] <= 8'h10 ;
			data[17937] <= 8'h10 ;
			data[17938] <= 8'h10 ;
			data[17939] <= 8'h10 ;
			data[17940] <= 8'h10 ;
			data[17941] <= 8'h10 ;
			data[17942] <= 8'h10 ;
			data[17943] <= 8'h10 ;
			data[17944] <= 8'h10 ;
			data[17945] <= 8'h10 ;
			data[17946] <= 8'h10 ;
			data[17947] <= 8'h10 ;
			data[17948] <= 8'h10 ;
			data[17949] <= 8'h10 ;
			data[17950] <= 8'h10 ;
			data[17951] <= 8'h10 ;
			data[17952] <= 8'h10 ;
			data[17953] <= 8'h10 ;
			data[17954] <= 8'h10 ;
			data[17955] <= 8'h10 ;
			data[17956] <= 8'h10 ;
			data[17957] <= 8'h10 ;
			data[17958] <= 8'h10 ;
			data[17959] <= 8'h10 ;
			data[17960] <= 8'h10 ;
			data[17961] <= 8'h10 ;
			data[17962] <= 8'h10 ;
			data[17963] <= 8'h10 ;
			data[17964] <= 8'h10 ;
			data[17965] <= 8'h10 ;
			data[17966] <= 8'h10 ;
			data[17967] <= 8'h10 ;
			data[17968] <= 8'h10 ;
			data[17969] <= 8'h10 ;
			data[17970] <= 8'h10 ;
			data[17971] <= 8'h10 ;
			data[17972] <= 8'h10 ;
			data[17973] <= 8'h10 ;
			data[17974] <= 8'h10 ;
			data[17975] <= 8'h10 ;
			data[17976] <= 8'h10 ;
			data[17977] <= 8'h10 ;
			data[17978] <= 8'h10 ;
			data[17979] <= 8'h10 ;
			data[17980] <= 8'h10 ;
			data[17981] <= 8'h10 ;
			data[17982] <= 8'h10 ;
			data[17983] <= 8'h10 ;
			data[17984] <= 8'h10 ;
			data[17985] <= 8'h10 ;
			data[17986] <= 8'h10 ;
			data[17987] <= 8'h10 ;
			data[17988] <= 8'h10 ;
			data[17989] <= 8'h10 ;
			data[17990] <= 8'h10 ;
			data[17991] <= 8'h10 ;
			data[17992] <= 8'h10 ;
			data[17993] <= 8'h10 ;
			data[17994] <= 8'h10 ;
			data[17995] <= 8'h10 ;
			data[17996] <= 8'h10 ;
			data[17997] <= 8'h10 ;
			data[17998] <= 8'h10 ;
			data[17999] <= 8'h10 ;
			data[18000] <= 8'h10 ;
			data[18001] <= 8'h10 ;
			data[18002] <= 8'h10 ;
			data[18003] <= 8'h10 ;
			data[18004] <= 8'h10 ;
			data[18005] <= 8'h10 ;
			data[18006] <= 8'h10 ;
			data[18007] <= 8'h10 ;
			data[18008] <= 8'h10 ;
			data[18009] <= 8'h10 ;
			data[18010] <= 8'h10 ;
			data[18011] <= 8'h10 ;
			data[18012] <= 8'h10 ;
			data[18013] <= 8'h10 ;
			data[18014] <= 8'h10 ;
			data[18015] <= 8'h10 ;
			data[18016] <= 8'h10 ;
			data[18017] <= 8'h10 ;
			data[18018] <= 8'h10 ;
			data[18019] <= 8'h10 ;
			data[18020] <= 8'h10 ;
			data[18021] <= 8'h10 ;
			data[18022] <= 8'h10 ;
			data[18023] <= 8'h10 ;
			data[18024] <= 8'h10 ;
			data[18025] <= 8'h10 ;
			data[18026] <= 8'h10 ;
			data[18027] <= 8'h10 ;
			data[18028] <= 8'h10 ;
			data[18029] <= 8'h10 ;
			data[18030] <= 8'h10 ;
			data[18031] <= 8'h10 ;
			data[18032] <= 8'h10 ;
			data[18033] <= 8'h10 ;
			data[18034] <= 8'h10 ;
			data[18035] <= 8'h10 ;
			data[18036] <= 8'h10 ;
			data[18037] <= 8'h10 ;
			data[18038] <= 8'h10 ;
			data[18039] <= 8'h10 ;
			data[18040] <= 8'h10 ;
			data[18041] <= 8'h10 ;
			data[18042] <= 8'h10 ;
			data[18043] <= 8'h10 ;
			data[18044] <= 8'h10 ;
			data[18045] <= 8'h10 ;
			data[18046] <= 8'h10 ;
			data[18047] <= 8'h10 ;
			data[18048] <= 8'h10 ;
			data[18049] <= 8'h10 ;
			data[18050] <= 8'h10 ;
			data[18051] <= 8'h10 ;
			data[18052] <= 8'h10 ;
			data[18053] <= 8'h10 ;
			data[18054] <= 8'h10 ;
			data[18055] <= 8'h10 ;
			data[18056] <= 8'h10 ;
			data[18057] <= 8'h10 ;
			data[18058] <= 8'h10 ;
			data[18059] <= 8'h10 ;
			data[18060] <= 8'h10 ;
			data[18061] <= 8'h10 ;
			data[18062] <= 8'h10 ;
			data[18063] <= 8'h10 ;
			data[18064] <= 8'h10 ;
			data[18065] <= 8'h10 ;
			data[18066] <= 8'h10 ;
			data[18067] <= 8'h10 ;
			data[18068] <= 8'h10 ;
			data[18069] <= 8'h10 ;
			data[18070] <= 8'h10 ;
			data[18071] <= 8'h10 ;
			data[18072] <= 8'h10 ;
			data[18073] <= 8'h10 ;
			data[18074] <= 8'h10 ;
			data[18075] <= 8'h10 ;
			data[18076] <= 8'h10 ;
			data[18077] <= 8'h10 ;
			data[18078] <= 8'h10 ;
			data[18079] <= 8'h10 ;
			data[18080] <= 8'h10 ;
			data[18081] <= 8'h10 ;
			data[18082] <= 8'h10 ;
			data[18083] <= 8'h10 ;
			data[18084] <= 8'h10 ;
			data[18085] <= 8'h10 ;
			data[18086] <= 8'h10 ;
			data[18087] <= 8'h10 ;
			data[18088] <= 8'h10 ;
			data[18089] <= 8'h10 ;
			data[18090] <= 8'h10 ;
			data[18091] <= 8'h10 ;
			data[18092] <= 8'h10 ;
			data[18093] <= 8'h10 ;
			data[18094] <= 8'h10 ;
			data[18095] <= 8'h10 ;
			data[18096] <= 8'h10 ;
			data[18097] <= 8'h10 ;
			data[18098] <= 8'h10 ;
			data[18099] <= 8'h10 ;
			data[18100] <= 8'h10 ;
			data[18101] <= 8'h10 ;
			data[18102] <= 8'h10 ;
			data[18103] <= 8'h10 ;
			data[18104] <= 8'h10 ;
			data[18105] <= 8'h10 ;
			data[18106] <= 8'h10 ;
			data[18107] <= 8'h10 ;
			data[18108] <= 8'h10 ;
			data[18109] <= 8'h10 ;
			data[18110] <= 8'h10 ;
			data[18111] <= 8'h10 ;
			data[18112] <= 8'h10 ;
			data[18113] <= 8'h10 ;
			data[18114] <= 8'h10 ;
			data[18115] <= 8'h10 ;
			data[18116] <= 8'h10 ;
			data[18117] <= 8'h10 ;
			data[18118] <= 8'h10 ;
			data[18119] <= 8'h10 ;
			data[18120] <= 8'h10 ;
			data[18121] <= 8'h10 ;
			data[18122] <= 8'h10 ;
			data[18123] <= 8'h10 ;
			data[18124] <= 8'h10 ;
			data[18125] <= 8'h10 ;
			data[18126] <= 8'h10 ;
			data[18127] <= 8'h10 ;
			data[18128] <= 8'h10 ;
			data[18129] <= 8'h10 ;
			data[18130] <= 8'h10 ;
			data[18131] <= 8'h10 ;
			data[18132] <= 8'h10 ;
			data[18133] <= 8'h10 ;
			data[18134] <= 8'h10 ;
			data[18135] <= 8'h10 ;
			data[18136] <= 8'h10 ;
			data[18137] <= 8'h10 ;
			data[18138] <= 8'h10 ;
			data[18139] <= 8'h10 ;
			data[18140] <= 8'h10 ;
			data[18141] <= 8'h10 ;
			data[18142] <= 8'h10 ;
			data[18143] <= 8'h10 ;
			data[18144] <= 8'h10 ;
			data[18145] <= 8'h10 ;
			data[18146] <= 8'h10 ;
			data[18147] <= 8'h10 ;
			data[18148] <= 8'h10 ;
			data[18149] <= 8'h10 ;
			data[18150] <= 8'h10 ;
			data[18151] <= 8'h10 ;
			data[18152] <= 8'h10 ;
			data[18153] <= 8'h10 ;
			data[18154] <= 8'h10 ;
			data[18155] <= 8'h10 ;
			data[18156] <= 8'h10 ;
			data[18157] <= 8'h10 ;
			data[18158] <= 8'h10 ;
			data[18159] <= 8'h10 ;
			data[18160] <= 8'h10 ;
			data[18161] <= 8'h10 ;
			data[18162] <= 8'h10 ;
			data[18163] <= 8'h10 ;
			data[18164] <= 8'h10 ;
			data[18165] <= 8'h10 ;
			data[18166] <= 8'h10 ;
			data[18167] <= 8'h10 ;
			data[18168] <= 8'h10 ;
			data[18169] <= 8'h10 ;
			data[18170] <= 8'h10 ;
			data[18171] <= 8'h10 ;
			data[18172] <= 8'h10 ;
			data[18173] <= 8'h10 ;
			data[18174] <= 8'h10 ;
			data[18175] <= 8'h10 ;
			data[18176] <= 8'h10 ;
			data[18177] <= 8'h10 ;
			data[18178] <= 8'h10 ;
			data[18179] <= 8'h10 ;
			data[18180] <= 8'h10 ;
			data[18181] <= 8'h10 ;
			data[18182] <= 8'h10 ;
			data[18183] <= 8'h10 ;
			data[18184] <= 8'h10 ;
			data[18185] <= 8'h10 ;
			data[18186] <= 8'h10 ;
			data[18187] <= 8'h10 ;
			data[18188] <= 8'h10 ;
			data[18189] <= 8'h10 ;
			data[18190] <= 8'h10 ;
			data[18191] <= 8'h10 ;
			data[18192] <= 8'h10 ;
			data[18193] <= 8'h10 ;
			data[18194] <= 8'h10 ;
			data[18195] <= 8'h10 ;
			data[18196] <= 8'h10 ;
			data[18197] <= 8'h10 ;
			data[18198] <= 8'h10 ;
			data[18199] <= 8'h10 ;
			data[18200] <= 8'h10 ;
			data[18201] <= 8'h10 ;
			data[18202] <= 8'h10 ;
			data[18203] <= 8'h10 ;
			data[18204] <= 8'h10 ;
			data[18205] <= 8'h10 ;
			data[18206] <= 8'h10 ;
			data[18207] <= 8'h10 ;
			data[18208] <= 8'h10 ;
			data[18209] <= 8'h10 ;
			data[18210] <= 8'h10 ;
			data[18211] <= 8'h10 ;
			data[18212] <= 8'h10 ;
			data[18213] <= 8'h10 ;
			data[18214] <= 8'h10 ;
			data[18215] <= 8'h10 ;
			data[18216] <= 8'h10 ;
			data[18217] <= 8'h10 ;
			data[18218] <= 8'h10 ;
			data[18219] <= 8'h10 ;
			data[18220] <= 8'h10 ;
			data[18221] <= 8'h10 ;
			data[18222] <= 8'h10 ;
			data[18223] <= 8'h10 ;
			data[18224] <= 8'h10 ;
			data[18225] <= 8'h10 ;
			data[18226] <= 8'h10 ;
			data[18227] <= 8'h10 ;
			data[18228] <= 8'h10 ;
			data[18229] <= 8'h10 ;
			data[18230] <= 8'h10 ;
			data[18231] <= 8'h10 ;
			data[18232] <= 8'h10 ;
			data[18233] <= 8'h10 ;
			data[18234] <= 8'h10 ;
			data[18235] <= 8'h10 ;
			data[18236] <= 8'h10 ;
			data[18237] <= 8'h10 ;
			data[18238] <= 8'h10 ;
			data[18239] <= 8'h10 ;
			data[18240] <= 8'h10 ;
			data[18241] <= 8'h10 ;
			data[18242] <= 8'h10 ;
			data[18243] <= 8'h10 ;
			data[18244] <= 8'h10 ;
			data[18245] <= 8'h10 ;
			data[18246] <= 8'h10 ;
			data[18247] <= 8'h10 ;
			data[18248] <= 8'h10 ;
			data[18249] <= 8'h10 ;
			data[18250] <= 8'h10 ;
			data[18251] <= 8'h10 ;
			data[18252] <= 8'h10 ;
			data[18253] <= 8'h10 ;
			data[18254] <= 8'h10 ;
			data[18255] <= 8'h10 ;
			data[18256] <= 8'h10 ;
			data[18257] <= 8'h10 ;
			data[18258] <= 8'h10 ;
			data[18259] <= 8'h10 ;
			data[18260] <= 8'h10 ;
			data[18261] <= 8'h10 ;
			data[18262] <= 8'h10 ;
			data[18263] <= 8'h10 ;
			data[18264] <= 8'h10 ;
			data[18265] <= 8'h10 ;
			data[18266] <= 8'h10 ;
			data[18267] <= 8'h10 ;
			data[18268] <= 8'h10 ;
			data[18269] <= 8'h10 ;
			data[18270] <= 8'h10 ;
			data[18271] <= 8'h10 ;
			data[18272] <= 8'h10 ;
			data[18273] <= 8'h10 ;
			data[18274] <= 8'h10 ;
			data[18275] <= 8'h10 ;
			data[18276] <= 8'h10 ;
			data[18277] <= 8'h10 ;
			data[18278] <= 8'h10 ;
			data[18279] <= 8'h10 ;
			data[18280] <= 8'h10 ;
			data[18281] <= 8'h10 ;
			data[18282] <= 8'h10 ;
			data[18283] <= 8'h10 ;
			data[18284] <= 8'h10 ;
			data[18285] <= 8'h10 ;
			data[18286] <= 8'h10 ;
			data[18287] <= 8'h10 ;
			data[18288] <= 8'h10 ;
			data[18289] <= 8'h10 ;
			data[18290] <= 8'h10 ;
			data[18291] <= 8'h10 ;
			data[18292] <= 8'h10 ;
			data[18293] <= 8'h10 ;
			data[18294] <= 8'h10 ;
			data[18295] <= 8'h10 ;
			data[18296] <= 8'h10 ;
			data[18297] <= 8'h10 ;
			data[18298] <= 8'h10 ;
			data[18299] <= 8'h10 ;
			data[18300] <= 8'h10 ;
			data[18301] <= 8'h10 ;
			data[18302] <= 8'h10 ;
			data[18303] <= 8'h10 ;
			data[18304] <= 8'h10 ;
			data[18305] <= 8'h10 ;
			data[18306] <= 8'h10 ;
			data[18307] <= 8'h10 ;
			data[18308] <= 8'h10 ;
			data[18309] <= 8'h10 ;
			data[18310] <= 8'h10 ;
			data[18311] <= 8'h10 ;
			data[18312] <= 8'h10 ;
			data[18313] <= 8'h10 ;
			data[18314] <= 8'h10 ;
			data[18315] <= 8'h10 ;
			data[18316] <= 8'h10 ;
			data[18317] <= 8'h10 ;
			data[18318] <= 8'h10 ;
			data[18319] <= 8'h10 ;
			data[18320] <= 8'h10 ;
			data[18321] <= 8'h10 ;
			data[18322] <= 8'h10 ;
			data[18323] <= 8'h10 ;
			data[18324] <= 8'h10 ;
			data[18325] <= 8'h10 ;
			data[18326] <= 8'h10 ;
			data[18327] <= 8'h10 ;
			data[18328] <= 8'h10 ;
			data[18329] <= 8'h10 ;
			data[18330] <= 8'h10 ;
			data[18331] <= 8'h10 ;
			data[18332] <= 8'h10 ;
			data[18333] <= 8'h10 ;
			data[18334] <= 8'h10 ;
			data[18335] <= 8'h10 ;
			data[18336] <= 8'h10 ;
			data[18337] <= 8'h10 ;
			data[18338] <= 8'h10 ;
			data[18339] <= 8'h10 ;
			data[18340] <= 8'h10 ;
			data[18341] <= 8'h10 ;
			data[18342] <= 8'h10 ;
			data[18343] <= 8'h10 ;
			data[18344] <= 8'h10 ;
			data[18345] <= 8'h10 ;
			data[18346] <= 8'h10 ;
			data[18347] <= 8'h10 ;
			data[18348] <= 8'h10 ;
			data[18349] <= 8'h10 ;
			data[18350] <= 8'h10 ;
			data[18351] <= 8'h10 ;
			data[18352] <= 8'h10 ;
			data[18353] <= 8'h10 ;
			data[18354] <= 8'h10 ;
			data[18355] <= 8'h10 ;
			data[18356] <= 8'h10 ;
			data[18357] <= 8'h10 ;
			data[18358] <= 8'h10 ;
			data[18359] <= 8'h10 ;
			data[18360] <= 8'h10 ;
			data[18361] <= 8'h10 ;
			data[18362] <= 8'h10 ;
			data[18363] <= 8'h10 ;
			data[18364] <= 8'h10 ;
			data[18365] <= 8'h10 ;
			data[18366] <= 8'h10 ;
			data[18367] <= 8'h10 ;
			data[18368] <= 8'h10 ;
			data[18369] <= 8'h10 ;
			data[18370] <= 8'h10 ;
			data[18371] <= 8'h10 ;
			data[18372] <= 8'h10 ;
			data[18373] <= 8'h10 ;
			data[18374] <= 8'h10 ;
			data[18375] <= 8'h10 ;
			data[18376] <= 8'h10 ;
			data[18377] <= 8'h10 ;
			data[18378] <= 8'h10 ;
			data[18379] <= 8'h10 ;
			data[18380] <= 8'h10 ;
			data[18381] <= 8'h10 ;
			data[18382] <= 8'h10 ;
			data[18383] <= 8'h10 ;
			data[18384] <= 8'h10 ;
			data[18385] <= 8'h10 ;
			data[18386] <= 8'h10 ;
			data[18387] <= 8'h10 ;
			data[18388] <= 8'h10 ;
			data[18389] <= 8'h10 ;
			data[18390] <= 8'h10 ;
			data[18391] <= 8'h10 ;
			data[18392] <= 8'h10 ;
			data[18393] <= 8'h10 ;
			data[18394] <= 8'h10 ;
			data[18395] <= 8'h10 ;
			data[18396] <= 8'h10 ;
			data[18397] <= 8'h10 ;
			data[18398] <= 8'h10 ;
			data[18399] <= 8'h10 ;
			data[18400] <= 8'h10 ;
			data[18401] <= 8'h10 ;
			data[18402] <= 8'h10 ;
			data[18403] <= 8'h10 ;
			data[18404] <= 8'h10 ;
			data[18405] <= 8'h10 ;
			data[18406] <= 8'h10 ;
			data[18407] <= 8'h10 ;
			data[18408] <= 8'h10 ;
			data[18409] <= 8'h10 ;
			data[18410] <= 8'h10 ;
			data[18411] <= 8'h10 ;
			data[18412] <= 8'h10 ;
			data[18413] <= 8'h10 ;
			data[18414] <= 8'h10 ;
			data[18415] <= 8'h10 ;
			data[18416] <= 8'h10 ;
			data[18417] <= 8'h10 ;
			data[18418] <= 8'h10 ;
			data[18419] <= 8'h10 ;
			data[18420] <= 8'h10 ;
			data[18421] <= 8'h10 ;
			data[18422] <= 8'h10 ;
			data[18423] <= 8'h10 ;
			data[18424] <= 8'h10 ;
			data[18425] <= 8'h10 ;
			data[18426] <= 8'h10 ;
			data[18427] <= 8'h10 ;
			data[18428] <= 8'h10 ;
			data[18429] <= 8'h10 ;
			data[18430] <= 8'h10 ;
			data[18431] <= 8'h10 ;
			data[18432] <= 8'h10 ;
			data[18433] <= 8'h10 ;
			data[18434] <= 8'h10 ;
			data[18435] <= 8'h10 ;
			data[18436] <= 8'h10 ;
			data[18437] <= 8'h10 ;
			data[18438] <= 8'h10 ;
			data[18439] <= 8'h10 ;
			data[18440] <= 8'h10 ;
			data[18441] <= 8'h10 ;
			data[18442] <= 8'h10 ;
			data[18443] <= 8'h10 ;
			data[18444] <= 8'h10 ;
			data[18445] <= 8'h10 ;
			data[18446] <= 8'h10 ;
			data[18447] <= 8'h10 ;
			data[18448] <= 8'h10 ;
			data[18449] <= 8'h10 ;
			data[18450] <= 8'h10 ;
			data[18451] <= 8'h10 ;
			data[18452] <= 8'h10 ;
			data[18453] <= 8'h10 ;
			data[18454] <= 8'h10 ;
			data[18455] <= 8'h10 ;
			data[18456] <= 8'h10 ;
			data[18457] <= 8'h10 ;
			data[18458] <= 8'h10 ;
			data[18459] <= 8'h10 ;
			data[18460] <= 8'h10 ;
			data[18461] <= 8'h10 ;
			data[18462] <= 8'h10 ;
			data[18463] <= 8'h10 ;
			data[18464] <= 8'h10 ;
			data[18465] <= 8'h10 ;
			data[18466] <= 8'h10 ;
			data[18467] <= 8'h10 ;
			data[18468] <= 8'h10 ;
			data[18469] <= 8'h10 ;
			data[18470] <= 8'h10 ;
			data[18471] <= 8'h10 ;
			data[18472] <= 8'h10 ;
			data[18473] <= 8'h10 ;
			data[18474] <= 8'h10 ;
			data[18475] <= 8'h10 ;
			data[18476] <= 8'h10 ;
			data[18477] <= 8'h10 ;
			data[18478] <= 8'h10 ;
			data[18479] <= 8'h10 ;
			data[18480] <= 8'h10 ;
			data[18481] <= 8'h10 ;
			data[18482] <= 8'h10 ;
			data[18483] <= 8'h10 ;
			data[18484] <= 8'h10 ;
			data[18485] <= 8'h10 ;
			data[18486] <= 8'h10 ;
			data[18487] <= 8'h10 ;
			data[18488] <= 8'h10 ;
			data[18489] <= 8'h10 ;
			data[18490] <= 8'h10 ;
			data[18491] <= 8'h10 ;
			data[18492] <= 8'h10 ;
			data[18493] <= 8'h10 ;
			data[18494] <= 8'h10 ;
			data[18495] <= 8'h10 ;
			data[18496] <= 8'h10 ;
			data[18497] <= 8'h10 ;
			data[18498] <= 8'h10 ;
			data[18499] <= 8'h10 ;
			data[18500] <= 8'h10 ;
			data[18501] <= 8'h10 ;
			data[18502] <= 8'h10 ;
			data[18503] <= 8'h10 ;
			data[18504] <= 8'h10 ;
			data[18505] <= 8'h10 ;
			data[18506] <= 8'h10 ;
			data[18507] <= 8'h10 ;
			data[18508] <= 8'h10 ;
			data[18509] <= 8'h10 ;
			data[18510] <= 8'h10 ;
			data[18511] <= 8'h10 ;
			data[18512] <= 8'h10 ;
			data[18513] <= 8'h10 ;
			data[18514] <= 8'h10 ;
			data[18515] <= 8'h10 ;
			data[18516] <= 8'h10 ;
			data[18517] <= 8'h10 ;
			data[18518] <= 8'h10 ;
			data[18519] <= 8'h10 ;
			data[18520] <= 8'h10 ;
			data[18521] <= 8'h10 ;
			data[18522] <= 8'h10 ;
			data[18523] <= 8'h10 ;
			data[18524] <= 8'h10 ;
			data[18525] <= 8'h10 ;
			data[18526] <= 8'h10 ;
			data[18527] <= 8'h10 ;
			data[18528] <= 8'h10 ;
			data[18529] <= 8'h10 ;
			data[18530] <= 8'h10 ;
			data[18531] <= 8'h10 ;
			data[18532] <= 8'h10 ;
			data[18533] <= 8'h10 ;
			data[18534] <= 8'h10 ;
			data[18535] <= 8'h10 ;
			data[18536] <= 8'h10 ;
			data[18537] <= 8'h10 ;
			data[18538] <= 8'h10 ;
			data[18539] <= 8'h10 ;
			data[18540] <= 8'h10 ;
			data[18541] <= 8'h10 ;
			data[18542] <= 8'h10 ;
			data[18543] <= 8'h10 ;
			data[18544] <= 8'h10 ;
			data[18545] <= 8'h10 ;
			data[18546] <= 8'h10 ;
			data[18547] <= 8'h10 ;
			data[18548] <= 8'h10 ;
			data[18549] <= 8'h10 ;
			data[18550] <= 8'h10 ;
			data[18551] <= 8'h10 ;
			data[18552] <= 8'h10 ;
			data[18553] <= 8'h10 ;
			data[18554] <= 8'h10 ;
			data[18555] <= 8'h10 ;
			data[18556] <= 8'h10 ;
			data[18557] <= 8'h10 ;
			data[18558] <= 8'h10 ;
			data[18559] <= 8'h10 ;
			data[18560] <= 8'h10 ;
			data[18561] <= 8'h10 ;
			data[18562] <= 8'h10 ;
			data[18563] <= 8'h10 ;
			data[18564] <= 8'h10 ;
			data[18565] <= 8'h10 ;
			data[18566] <= 8'h10 ;
			data[18567] <= 8'h10 ;
			data[18568] <= 8'h10 ;
			data[18569] <= 8'h10 ;
			data[18570] <= 8'h10 ;
			data[18571] <= 8'h10 ;
			data[18572] <= 8'h10 ;
			data[18573] <= 8'h10 ;
			data[18574] <= 8'h10 ;
			data[18575] <= 8'h10 ;
			data[18576] <= 8'h10 ;
			data[18577] <= 8'h10 ;
			data[18578] <= 8'h10 ;
			data[18579] <= 8'h10 ;
			data[18580] <= 8'h10 ;
			data[18581] <= 8'h10 ;
			data[18582] <= 8'h10 ;
			data[18583] <= 8'h10 ;
			data[18584] <= 8'h10 ;
			data[18585] <= 8'h10 ;
			data[18586] <= 8'h10 ;
			data[18587] <= 8'h10 ;
			data[18588] <= 8'h10 ;
			data[18589] <= 8'h10 ;
			data[18590] <= 8'h10 ;
			data[18591] <= 8'h10 ;
			data[18592] <= 8'h10 ;
			data[18593] <= 8'h10 ;
			data[18594] <= 8'h10 ;
			data[18595] <= 8'h10 ;
			data[18596] <= 8'h10 ;
			data[18597] <= 8'h10 ;
			data[18598] <= 8'h10 ;
			data[18599] <= 8'h10 ;
			data[18600] <= 8'h10 ;
			data[18601] <= 8'h10 ;
			data[18602] <= 8'h10 ;
			data[18603] <= 8'h10 ;
			data[18604] <= 8'h10 ;
			data[18605] <= 8'h10 ;
			data[18606] <= 8'h10 ;
			data[18607] <= 8'h10 ;
			data[18608] <= 8'h10 ;
			data[18609] <= 8'h10 ;
			data[18610] <= 8'h10 ;
			data[18611] <= 8'h10 ;
			data[18612] <= 8'h10 ;
			data[18613] <= 8'h10 ;
			data[18614] <= 8'h10 ;
			data[18615] <= 8'h10 ;
			data[18616] <= 8'h10 ;
			data[18617] <= 8'h10 ;
			data[18618] <= 8'h10 ;
			data[18619] <= 8'h10 ;
			data[18620] <= 8'h10 ;
			data[18621] <= 8'h10 ;
			data[18622] <= 8'h10 ;
			data[18623] <= 8'h10 ;
			data[18624] <= 8'h10 ;
			data[18625] <= 8'h10 ;
			data[18626] <= 8'h10 ;
			data[18627] <= 8'h10 ;
			data[18628] <= 8'h10 ;
			data[18629] <= 8'h10 ;
			data[18630] <= 8'h10 ;
			data[18631] <= 8'h10 ;
			data[18632] <= 8'h10 ;
			data[18633] <= 8'h10 ;
			data[18634] <= 8'h10 ;
			data[18635] <= 8'h10 ;
			data[18636] <= 8'h10 ;
			data[18637] <= 8'h10 ;
			data[18638] <= 8'h10 ;
			data[18639] <= 8'h10 ;
			data[18640] <= 8'h10 ;
			data[18641] <= 8'h10 ;
			data[18642] <= 8'h10 ;
			data[18643] <= 8'h10 ;
			data[18644] <= 8'h10 ;
			data[18645] <= 8'h10 ;
			data[18646] <= 8'h10 ;
			data[18647] <= 8'h10 ;
			data[18648] <= 8'h10 ;
			data[18649] <= 8'h10 ;
			data[18650] <= 8'h10 ;
			data[18651] <= 8'h10 ;
			data[18652] <= 8'h10 ;
			data[18653] <= 8'h10 ;
			data[18654] <= 8'h10 ;
			data[18655] <= 8'h10 ;
			data[18656] <= 8'h10 ;
			data[18657] <= 8'h10 ;
			data[18658] <= 8'h10 ;
			data[18659] <= 8'h10 ;
			data[18660] <= 8'h10 ;
			data[18661] <= 8'h10 ;
			data[18662] <= 8'h10 ;
			data[18663] <= 8'h10 ;
			data[18664] <= 8'h10 ;
			data[18665] <= 8'h10 ;
			data[18666] <= 8'h10 ;
			data[18667] <= 8'h10 ;
			data[18668] <= 8'h10 ;
			data[18669] <= 8'h10 ;
			data[18670] <= 8'h10 ;
			data[18671] <= 8'h10 ;
			data[18672] <= 8'h10 ;
			data[18673] <= 8'h10 ;
			data[18674] <= 8'h10 ;
			data[18675] <= 8'h10 ;
			data[18676] <= 8'h10 ;
			data[18677] <= 8'h10 ;
			data[18678] <= 8'h10 ;
			data[18679] <= 8'h10 ;
			data[18680] <= 8'h10 ;
			data[18681] <= 8'h10 ;
			data[18682] <= 8'h10 ;
			data[18683] <= 8'h10 ;
			data[18684] <= 8'h10 ;
			data[18685] <= 8'h10 ;
			data[18686] <= 8'h10 ;
			data[18687] <= 8'h10 ;
			data[18688] <= 8'h10 ;
			data[18689] <= 8'h10 ;
			data[18690] <= 8'h10 ;
			data[18691] <= 8'h10 ;
			data[18692] <= 8'h10 ;
			data[18693] <= 8'h10 ;
			data[18694] <= 8'h10 ;
			data[18695] <= 8'h10 ;
			data[18696] <= 8'h10 ;
			data[18697] <= 8'h10 ;
			data[18698] <= 8'h10 ;
			data[18699] <= 8'h10 ;
			data[18700] <= 8'h10 ;
			data[18701] <= 8'h10 ;
			data[18702] <= 8'h10 ;
			data[18703] <= 8'h10 ;
			data[18704] <= 8'h10 ;
			data[18705] <= 8'h10 ;
			data[18706] <= 8'h10 ;
			data[18707] <= 8'h10 ;
			data[18708] <= 8'h10 ;
			data[18709] <= 8'h10 ;
			data[18710] <= 8'h10 ;
			data[18711] <= 8'h10 ;
			data[18712] <= 8'h10 ;
			data[18713] <= 8'h10 ;
			data[18714] <= 8'h10 ;
			data[18715] <= 8'h10 ;
			data[18716] <= 8'h10 ;
			data[18717] <= 8'h10 ;
			data[18718] <= 8'h10 ;
			data[18719] <= 8'h10 ;
			data[18720] <= 8'h10 ;
			data[18721] <= 8'h10 ;
			data[18722] <= 8'h10 ;
			data[18723] <= 8'h10 ;
			data[18724] <= 8'h10 ;
			data[18725] <= 8'h10 ;
			data[18726] <= 8'h10 ;
			data[18727] <= 8'h10 ;
			data[18728] <= 8'h10 ;
			data[18729] <= 8'h10 ;
			data[18730] <= 8'h10 ;
			data[18731] <= 8'h10 ;
			data[18732] <= 8'h10 ;
			data[18733] <= 8'h10 ;
			data[18734] <= 8'h10 ;
			data[18735] <= 8'h10 ;
			data[18736] <= 8'h10 ;
			data[18737] <= 8'h10 ;
			data[18738] <= 8'h10 ;
			data[18739] <= 8'h10 ;
			data[18740] <= 8'h10 ;
			data[18741] <= 8'h10 ;
			data[18742] <= 8'h10 ;
			data[18743] <= 8'h10 ;
			data[18744] <= 8'h10 ;
			data[18745] <= 8'h10 ;
			data[18746] <= 8'h10 ;
			data[18747] <= 8'h10 ;
			data[18748] <= 8'h10 ;
			data[18749] <= 8'h10 ;
			data[18750] <= 8'h10 ;
			data[18751] <= 8'h10 ;
			data[18752] <= 8'h10 ;
			data[18753] <= 8'h10 ;
			data[18754] <= 8'h10 ;
			data[18755] <= 8'h10 ;
			data[18756] <= 8'h10 ;
			data[18757] <= 8'h10 ;
			data[18758] <= 8'h10 ;
			data[18759] <= 8'h10 ;
			data[18760] <= 8'h10 ;
			data[18761] <= 8'h10 ;
			data[18762] <= 8'h10 ;
			data[18763] <= 8'h10 ;
			data[18764] <= 8'h10 ;
			data[18765] <= 8'h10 ;
			data[18766] <= 8'h10 ;
			data[18767] <= 8'h10 ;
			data[18768] <= 8'h10 ;
			data[18769] <= 8'h10 ;
			data[18770] <= 8'h10 ;
			data[18771] <= 8'h10 ;
			data[18772] <= 8'h10 ;
			data[18773] <= 8'h10 ;
			data[18774] <= 8'h10 ;
			data[18775] <= 8'h10 ;
			data[18776] <= 8'h10 ;
			data[18777] <= 8'h10 ;
			data[18778] <= 8'h10 ;
			data[18779] <= 8'h10 ;
			data[18780] <= 8'h10 ;
			data[18781] <= 8'h10 ;
			data[18782] <= 8'h10 ;
			data[18783] <= 8'h10 ;
			data[18784] <= 8'h10 ;
			data[18785] <= 8'h10 ;
			data[18786] <= 8'h10 ;
			data[18787] <= 8'h10 ;
			data[18788] <= 8'h10 ;
			data[18789] <= 8'h10 ;
			data[18790] <= 8'h10 ;
			data[18791] <= 8'h10 ;
			data[18792] <= 8'h10 ;
			data[18793] <= 8'h10 ;
			data[18794] <= 8'h10 ;
			data[18795] <= 8'h10 ;
			data[18796] <= 8'h10 ;
			data[18797] <= 8'h10 ;
			data[18798] <= 8'h10 ;
			data[18799] <= 8'h10 ;
			data[18800] <= 8'h10 ;
			data[18801] <= 8'h10 ;
			data[18802] <= 8'h10 ;
			data[18803] <= 8'h10 ;
			data[18804] <= 8'h10 ;
			data[18805] <= 8'h10 ;
			data[18806] <= 8'h10 ;
			data[18807] <= 8'h10 ;
			data[18808] <= 8'h10 ;
			data[18809] <= 8'h10 ;
			data[18810] <= 8'h10 ;
			data[18811] <= 8'h10 ;
			data[18812] <= 8'h10 ;
			data[18813] <= 8'h10 ;
			data[18814] <= 8'h10 ;
			data[18815] <= 8'h10 ;
			data[18816] <= 8'h10 ;
			data[18817] <= 8'h10 ;
			data[18818] <= 8'h10 ;
			data[18819] <= 8'h10 ;
			data[18820] <= 8'h10 ;
			data[18821] <= 8'h10 ;
			data[18822] <= 8'h10 ;
			data[18823] <= 8'h10 ;
			data[18824] <= 8'h10 ;
			data[18825] <= 8'h10 ;
			data[18826] <= 8'h10 ;
			data[18827] <= 8'h10 ;
			data[18828] <= 8'h10 ;
			data[18829] <= 8'h10 ;
			data[18830] <= 8'h10 ;
			data[18831] <= 8'h10 ;
			data[18832] <= 8'h10 ;
			data[18833] <= 8'h10 ;
			data[18834] <= 8'h10 ;
			data[18835] <= 8'h10 ;
			data[18836] <= 8'h10 ;
			data[18837] <= 8'h10 ;
			data[18838] <= 8'h10 ;
			data[18839] <= 8'h10 ;
			data[18840] <= 8'h10 ;
			data[18841] <= 8'h10 ;
			data[18842] <= 8'h10 ;
			data[18843] <= 8'h10 ;
			data[18844] <= 8'h10 ;
			data[18845] <= 8'h10 ;
			data[18846] <= 8'h10 ;
			data[18847] <= 8'h10 ;
			data[18848] <= 8'h10 ;
			data[18849] <= 8'h10 ;
			data[18850] <= 8'h10 ;
			data[18851] <= 8'h10 ;
			data[18852] <= 8'h10 ;
			data[18853] <= 8'h10 ;
			data[18854] <= 8'h10 ;
			data[18855] <= 8'h10 ;
			data[18856] <= 8'h10 ;
			data[18857] <= 8'h10 ;
			data[18858] <= 8'h10 ;
			data[18859] <= 8'h10 ;
			data[18860] <= 8'h10 ;
			data[18861] <= 8'h10 ;
			data[18862] <= 8'h10 ;
			data[18863] <= 8'h10 ;
			data[18864] <= 8'h10 ;
			data[18865] <= 8'h10 ;
			data[18866] <= 8'h10 ;
			data[18867] <= 8'h10 ;
			data[18868] <= 8'h10 ;
			data[18869] <= 8'h10 ;
			data[18870] <= 8'h10 ;
			data[18871] <= 8'h10 ;
			data[18872] <= 8'h10 ;
			data[18873] <= 8'h10 ;
			data[18874] <= 8'h10 ;
			data[18875] <= 8'h10 ;
			data[18876] <= 8'h10 ;
			data[18877] <= 8'h10 ;
			data[18878] <= 8'h10 ;
			data[18879] <= 8'h10 ;
			data[18880] <= 8'h10 ;
			data[18881] <= 8'h10 ;
			data[18882] <= 8'h10 ;
			data[18883] <= 8'h10 ;
			data[18884] <= 8'h10 ;
			data[18885] <= 8'h10 ;
			data[18886] <= 8'h10 ;
			data[18887] <= 8'h10 ;
			data[18888] <= 8'h10 ;
			data[18889] <= 8'h10 ;
			data[18890] <= 8'h10 ;
			data[18891] <= 8'h10 ;
			data[18892] <= 8'h10 ;
			data[18893] <= 8'h10 ;
			data[18894] <= 8'h10 ;
			data[18895] <= 8'h10 ;
			data[18896] <= 8'h10 ;
			data[18897] <= 8'h10 ;
			data[18898] <= 8'h10 ;
			data[18899] <= 8'h10 ;
			data[18900] <= 8'h10 ;
			data[18901] <= 8'h10 ;
			data[18902] <= 8'h10 ;
			data[18903] <= 8'h10 ;
			data[18904] <= 8'h10 ;
			data[18905] <= 8'h10 ;
			data[18906] <= 8'h10 ;
			data[18907] <= 8'h10 ;
			data[18908] <= 8'h10 ;
			data[18909] <= 8'h10 ;
			data[18910] <= 8'h10 ;
			data[18911] <= 8'h10 ;
			data[18912] <= 8'h10 ;
			data[18913] <= 8'h10 ;
			data[18914] <= 8'h10 ;
			data[18915] <= 8'h10 ;
			data[18916] <= 8'h10 ;
			data[18917] <= 8'h10 ;
			data[18918] <= 8'h10 ;
			data[18919] <= 8'h10 ;
			data[18920] <= 8'h10 ;
			data[18921] <= 8'h10 ;
			data[18922] <= 8'h10 ;
			data[18923] <= 8'h10 ;
			data[18924] <= 8'h10 ;
			data[18925] <= 8'h10 ;
			data[18926] <= 8'h10 ;
			data[18927] <= 8'h10 ;
			data[18928] <= 8'h10 ;
			data[18929] <= 8'h10 ;
			data[18930] <= 8'h10 ;
			data[18931] <= 8'h10 ;
			data[18932] <= 8'h10 ;
			data[18933] <= 8'h10 ;
			data[18934] <= 8'h10 ;
			data[18935] <= 8'h10 ;
			data[18936] <= 8'h10 ;
			data[18937] <= 8'h10 ;
			data[18938] <= 8'h10 ;
			data[18939] <= 8'h10 ;
			data[18940] <= 8'h10 ;
			data[18941] <= 8'h10 ;
			data[18942] <= 8'h10 ;
			data[18943] <= 8'h10 ;
			data[18944] <= 8'h10 ;
			data[18945] <= 8'h10 ;
			data[18946] <= 8'h10 ;
			data[18947] <= 8'h10 ;
			data[18948] <= 8'h10 ;
			data[18949] <= 8'h10 ;
			data[18950] <= 8'h10 ;
			data[18951] <= 8'h10 ;
			data[18952] <= 8'h10 ;
			data[18953] <= 8'h10 ;
			data[18954] <= 8'h10 ;
			data[18955] <= 8'h10 ;
			data[18956] <= 8'h10 ;
			data[18957] <= 8'h10 ;
			data[18958] <= 8'h10 ;
			data[18959] <= 8'h10 ;
			data[18960] <= 8'h10 ;
			data[18961] <= 8'h10 ;
			data[18962] <= 8'h10 ;
			data[18963] <= 8'h10 ;
			data[18964] <= 8'h10 ;
			data[18965] <= 8'h10 ;
			data[18966] <= 8'h10 ;
			data[18967] <= 8'h10 ;
			data[18968] <= 8'h10 ;
			data[18969] <= 8'h10 ;
			data[18970] <= 8'h10 ;
			data[18971] <= 8'h10 ;
			data[18972] <= 8'h10 ;
			data[18973] <= 8'h10 ;
			data[18974] <= 8'h10 ;
			data[18975] <= 8'h10 ;
			data[18976] <= 8'h10 ;
			data[18977] <= 8'h10 ;
			data[18978] <= 8'h10 ;
			data[18979] <= 8'h10 ;
			data[18980] <= 8'h10 ;
			data[18981] <= 8'h10 ;
			data[18982] <= 8'h10 ;
			data[18983] <= 8'h10 ;
			data[18984] <= 8'h10 ;
			data[18985] <= 8'h10 ;
			data[18986] <= 8'h10 ;
			data[18987] <= 8'h10 ;
			data[18988] <= 8'h10 ;
			data[18989] <= 8'h10 ;
			data[18990] <= 8'h10 ;
			data[18991] <= 8'h10 ;
			data[18992] <= 8'h10 ;
			data[18993] <= 8'h10 ;
			data[18994] <= 8'h10 ;
			data[18995] <= 8'h10 ;
			data[18996] <= 8'h10 ;
			data[18997] <= 8'h10 ;
			data[18998] <= 8'h10 ;
			data[18999] <= 8'h10 ;
			data[19000] <= 8'h10 ;
			data[19001] <= 8'h10 ;
			data[19002] <= 8'h10 ;
			data[19003] <= 8'h10 ;
			data[19004] <= 8'h10 ;
			data[19005] <= 8'h10 ;
			data[19006] <= 8'h10 ;
			data[19007] <= 8'h10 ;
			data[19008] <= 8'h10 ;
			data[19009] <= 8'h10 ;
			data[19010] <= 8'h10 ;
			data[19011] <= 8'h10 ;
			data[19012] <= 8'h10 ;
			data[19013] <= 8'h10 ;
			data[19014] <= 8'h10 ;
			data[19015] <= 8'h10 ;
			data[19016] <= 8'h10 ;
			data[19017] <= 8'h10 ;
			data[19018] <= 8'h10 ;
			data[19019] <= 8'h10 ;
			data[19020] <= 8'h10 ;
			data[19021] <= 8'h10 ;
			data[19022] <= 8'h10 ;
			data[19023] <= 8'h10 ;
			data[19024] <= 8'h10 ;
			data[19025] <= 8'h10 ;
			data[19026] <= 8'h10 ;
			data[19027] <= 8'h10 ;
			data[19028] <= 8'h10 ;
			data[19029] <= 8'h10 ;
			data[19030] <= 8'h10 ;
			data[19031] <= 8'h10 ;
			data[19032] <= 8'h10 ;
			data[19033] <= 8'h10 ;
			data[19034] <= 8'h10 ;
			data[19035] <= 8'h10 ;
			data[19036] <= 8'h10 ;
			data[19037] <= 8'h10 ;
			data[19038] <= 8'h10 ;
			data[19039] <= 8'h10 ;
			data[19040] <= 8'h10 ;
			data[19041] <= 8'h10 ;
			data[19042] <= 8'h10 ;
			data[19043] <= 8'h10 ;
			data[19044] <= 8'h10 ;
			data[19045] <= 8'h10 ;
			data[19046] <= 8'h10 ;
			data[19047] <= 8'h10 ;
			data[19048] <= 8'h10 ;
			data[19049] <= 8'h10 ;
			data[19050] <= 8'h10 ;
			data[19051] <= 8'h10 ;
			data[19052] <= 8'h10 ;
			data[19053] <= 8'h10 ;
			data[19054] <= 8'h10 ;
			data[19055] <= 8'h10 ;
			data[19056] <= 8'h10 ;
			data[19057] <= 8'h10 ;
			data[19058] <= 8'h10 ;
			data[19059] <= 8'h10 ;
			data[19060] <= 8'h10 ;
			data[19061] <= 8'h10 ;
			data[19062] <= 8'h10 ;
			data[19063] <= 8'h10 ;
			data[19064] <= 8'h10 ;
			data[19065] <= 8'h10 ;
			data[19066] <= 8'h10 ;
			data[19067] <= 8'h10 ;
			data[19068] <= 8'h10 ;
			data[19069] <= 8'h10 ;
			data[19070] <= 8'h10 ;
			data[19071] <= 8'h10 ;
			data[19072] <= 8'h10 ;
			data[19073] <= 8'h10 ;
			data[19074] <= 8'h10 ;
			data[19075] <= 8'h10 ;
			data[19076] <= 8'h10 ;
			data[19077] <= 8'h10 ;
			data[19078] <= 8'h10 ;
			data[19079] <= 8'h10 ;
			data[19080] <= 8'h10 ;
			data[19081] <= 8'h10 ;
			data[19082] <= 8'h10 ;
			data[19083] <= 8'h10 ;
			data[19084] <= 8'h10 ;
			data[19085] <= 8'h10 ;
			data[19086] <= 8'h10 ;
			data[19087] <= 8'h10 ;
			data[19088] <= 8'h10 ;
			data[19089] <= 8'h10 ;
			data[19090] <= 8'h10 ;
			data[19091] <= 8'h10 ;
			data[19092] <= 8'h10 ;
			data[19093] <= 8'h10 ;
			data[19094] <= 8'h10 ;
			data[19095] <= 8'h10 ;
			data[19096] <= 8'h10 ;
			data[19097] <= 8'h10 ;
			data[19098] <= 8'h10 ;
			data[19099] <= 8'h10 ;
			data[19100] <= 8'h10 ;
			data[19101] <= 8'h10 ;
			data[19102] <= 8'h10 ;
			data[19103] <= 8'h10 ;
			data[19104] <= 8'h10 ;
			data[19105] <= 8'h10 ;
			data[19106] <= 8'h10 ;
			data[19107] <= 8'h10 ;
			data[19108] <= 8'h10 ;
			data[19109] <= 8'h10 ;
			data[19110] <= 8'h10 ;
			data[19111] <= 8'h10 ;
			data[19112] <= 8'h10 ;
			data[19113] <= 8'h10 ;
			data[19114] <= 8'h10 ;
			data[19115] <= 8'h10 ;
			data[19116] <= 8'h10 ;
			data[19117] <= 8'h10 ;
			data[19118] <= 8'h10 ;
			data[19119] <= 8'h10 ;
			data[19120] <= 8'h10 ;
			data[19121] <= 8'h10 ;
			data[19122] <= 8'h10 ;
			data[19123] <= 8'h10 ;
			data[19124] <= 8'h10 ;
			data[19125] <= 8'h10 ;
			data[19126] <= 8'h10 ;
			data[19127] <= 8'h10 ;
			data[19128] <= 8'h10 ;
			data[19129] <= 8'h10 ;
			data[19130] <= 8'h10 ;
			data[19131] <= 8'h10 ;
			data[19132] <= 8'h10 ;
			data[19133] <= 8'h10 ;
			data[19134] <= 8'h10 ;
			data[19135] <= 8'h10 ;
			data[19136] <= 8'h10 ;
			data[19137] <= 8'h10 ;
			data[19138] <= 8'h10 ;
			data[19139] <= 8'h10 ;
			data[19140] <= 8'h10 ;
			data[19141] <= 8'h10 ;
			data[19142] <= 8'h10 ;
			data[19143] <= 8'h10 ;
			data[19144] <= 8'h10 ;
			data[19145] <= 8'h10 ;
			data[19146] <= 8'h10 ;
			data[19147] <= 8'h10 ;
			data[19148] <= 8'h10 ;
			data[19149] <= 8'h10 ;
			data[19150] <= 8'h10 ;
			data[19151] <= 8'h10 ;
			data[19152] <= 8'h10 ;
			data[19153] <= 8'h10 ;
			data[19154] <= 8'h10 ;
			data[19155] <= 8'h10 ;
			data[19156] <= 8'h10 ;
			data[19157] <= 8'h10 ;
			data[19158] <= 8'h10 ;
			data[19159] <= 8'h10 ;
			data[19160] <= 8'h10 ;
			data[19161] <= 8'h10 ;
			data[19162] <= 8'h10 ;
			data[19163] <= 8'h10 ;
			data[19164] <= 8'h10 ;
			data[19165] <= 8'h10 ;
			data[19166] <= 8'h10 ;
			data[19167] <= 8'h10 ;
			data[19168] <= 8'h10 ;
			data[19169] <= 8'h10 ;
			data[19170] <= 8'h10 ;
			data[19171] <= 8'h10 ;
			data[19172] <= 8'h10 ;
			data[19173] <= 8'h10 ;
			data[19174] <= 8'h10 ;
			data[19175] <= 8'h10 ;
			data[19176] <= 8'h10 ;
			data[19177] <= 8'h10 ;
			data[19178] <= 8'h10 ;
			data[19179] <= 8'h10 ;
			data[19180] <= 8'h10 ;
			data[19181] <= 8'h10 ;
			data[19182] <= 8'h10 ;
			data[19183] <= 8'h10 ;
			data[19184] <= 8'h10 ;
			data[19185] <= 8'h10 ;
			data[19186] <= 8'h10 ;
			data[19187] <= 8'h10 ;
			data[19188] <= 8'h10 ;
			data[19189] <= 8'h10 ;
			data[19190] <= 8'h10 ;
			data[19191] <= 8'h10 ;
			data[19192] <= 8'h10 ;
			data[19193] <= 8'h10 ;
			data[19194] <= 8'h10 ;
			data[19195] <= 8'h10 ;
			data[19196] <= 8'h10 ;
			data[19197] <= 8'h10 ;
			data[19198] <= 8'h10 ;
			data[19199] <= 8'h10 ;
			data[19200] <= 8'h10 ;
			data[19201] <= 8'h10 ;
			data[19202] <= 8'h10 ;
			data[19203] <= 8'h10 ;
			data[19204] <= 8'h10 ;
			data[19205] <= 8'h10 ;
			data[19206] <= 8'h10 ;
			data[19207] <= 8'h10 ;
			data[19208] <= 8'h10 ;
			data[19209] <= 8'h10 ;
			data[19210] <= 8'h10 ;
			data[19211] <= 8'h10 ;
			data[19212] <= 8'h10 ;
			data[19213] <= 8'h10 ;
			data[19214] <= 8'h10 ;
			data[19215] <= 8'h10 ;
			data[19216] <= 8'h10 ;
			data[19217] <= 8'h10 ;
			data[19218] <= 8'h10 ;
			data[19219] <= 8'h10 ;
			data[19220] <= 8'h10 ;
			data[19221] <= 8'h10 ;
			data[19222] <= 8'h10 ;
			data[19223] <= 8'h10 ;
			data[19224] <= 8'h10 ;
			data[19225] <= 8'h10 ;
			data[19226] <= 8'h10 ;
			data[19227] <= 8'h10 ;
			data[19228] <= 8'h10 ;
			data[19229] <= 8'h10 ;
			data[19230] <= 8'h10 ;
			data[19231] <= 8'h10 ;
			data[19232] <= 8'h10 ;
			data[19233] <= 8'h10 ;
			data[19234] <= 8'h10 ;
			data[19235] <= 8'h10 ;
			data[19236] <= 8'h10 ;
			data[19237] <= 8'h10 ;
			data[19238] <= 8'h10 ;
			data[19239] <= 8'h10 ;
			data[19240] <= 8'h10 ;
			data[19241] <= 8'h10 ;
			data[19242] <= 8'h10 ;
			data[19243] <= 8'h10 ;
			data[19244] <= 8'h10 ;
			data[19245] <= 8'h10 ;
			data[19246] <= 8'h10 ;
			data[19247] <= 8'h10 ;
			data[19248] <= 8'h10 ;
			data[19249] <= 8'h10 ;
			data[19250] <= 8'h10 ;
			data[19251] <= 8'h10 ;
			data[19252] <= 8'h10 ;
			data[19253] <= 8'h10 ;
			data[19254] <= 8'h10 ;
			data[19255] <= 8'h10 ;
			data[19256] <= 8'h10 ;
			data[19257] <= 8'h10 ;
			data[19258] <= 8'h10 ;
			data[19259] <= 8'h10 ;
			data[19260] <= 8'h10 ;
			data[19261] <= 8'h10 ;
			data[19262] <= 8'h10 ;
			data[19263] <= 8'h10 ;
			data[19264] <= 8'h10 ;
			data[19265] <= 8'h10 ;
			data[19266] <= 8'h10 ;
			data[19267] <= 8'h10 ;
			data[19268] <= 8'h10 ;
			data[19269] <= 8'h10 ;
			data[19270] <= 8'h10 ;
			data[19271] <= 8'h10 ;
			data[19272] <= 8'h10 ;
			data[19273] <= 8'h10 ;
			data[19274] <= 8'h10 ;
			data[19275] <= 8'h10 ;
			data[19276] <= 8'h10 ;
			data[19277] <= 8'h10 ;
			data[19278] <= 8'h10 ;
			data[19279] <= 8'h10 ;
			data[19280] <= 8'h10 ;
			data[19281] <= 8'h10 ;
			data[19282] <= 8'h10 ;
			data[19283] <= 8'h10 ;
			data[19284] <= 8'h10 ;
			data[19285] <= 8'h10 ;
			data[19286] <= 8'h10 ;
			data[19287] <= 8'h10 ;
			data[19288] <= 8'h10 ;
			data[19289] <= 8'h10 ;
			data[19290] <= 8'h10 ;
			data[19291] <= 8'h10 ;
			data[19292] <= 8'h10 ;
			data[19293] <= 8'h10 ;
			data[19294] <= 8'h10 ;
			data[19295] <= 8'h10 ;
			data[19296] <= 8'h10 ;
			data[19297] <= 8'h10 ;
			data[19298] <= 8'h10 ;
			data[19299] <= 8'h10 ;
			data[19300] <= 8'h10 ;
			data[19301] <= 8'h10 ;
			data[19302] <= 8'h10 ;
			data[19303] <= 8'h10 ;
			data[19304] <= 8'h10 ;
			data[19305] <= 8'h10 ;
			data[19306] <= 8'h10 ;
			data[19307] <= 8'h10 ;
			data[19308] <= 8'h10 ;
			data[19309] <= 8'h10 ;
			data[19310] <= 8'h10 ;
			data[19311] <= 8'h10 ;
			data[19312] <= 8'h10 ;
			data[19313] <= 8'h10 ;
			data[19314] <= 8'h10 ;
			data[19315] <= 8'h10 ;
			data[19316] <= 8'h10 ;
			data[19317] <= 8'h10 ;
			data[19318] <= 8'h10 ;
			data[19319] <= 8'h10 ;
			data[19320] <= 8'h10 ;
			data[19321] <= 8'h10 ;
			data[19322] <= 8'h10 ;
			data[19323] <= 8'h10 ;
			data[19324] <= 8'h10 ;
			data[19325] <= 8'h10 ;
			data[19326] <= 8'h10 ;
			data[19327] <= 8'h10 ;
			data[19328] <= 8'h10 ;
			data[19329] <= 8'h10 ;
			data[19330] <= 8'h10 ;
			data[19331] <= 8'h10 ;
			data[19332] <= 8'h10 ;
			data[19333] <= 8'h10 ;
			data[19334] <= 8'h10 ;
			data[19335] <= 8'h10 ;
			data[19336] <= 8'h10 ;
			data[19337] <= 8'h10 ;
			data[19338] <= 8'h10 ;
			data[19339] <= 8'h10 ;
			data[19340] <= 8'h10 ;
			data[19341] <= 8'h10 ;
			data[19342] <= 8'h10 ;
			data[19343] <= 8'h10 ;
			data[19344] <= 8'h10 ;
			data[19345] <= 8'h10 ;
			data[19346] <= 8'h10 ;
			data[19347] <= 8'h10 ;
			data[19348] <= 8'h10 ;
			data[19349] <= 8'h10 ;
			data[19350] <= 8'h10 ;
			data[19351] <= 8'h10 ;
			data[19352] <= 8'h10 ;
			data[19353] <= 8'h10 ;
			data[19354] <= 8'h10 ;
			data[19355] <= 8'h10 ;
			data[19356] <= 8'h10 ;
			data[19357] <= 8'h10 ;
			data[19358] <= 8'h10 ;
			data[19359] <= 8'h10 ;
			data[19360] <= 8'h10 ;
			data[19361] <= 8'h10 ;
			data[19362] <= 8'h10 ;
			data[19363] <= 8'h10 ;
			data[19364] <= 8'h10 ;
			data[19365] <= 8'h10 ;
			data[19366] <= 8'h10 ;
			data[19367] <= 8'h10 ;
			data[19368] <= 8'h10 ;
			data[19369] <= 8'h10 ;
			data[19370] <= 8'h10 ;
			data[19371] <= 8'h10 ;
			data[19372] <= 8'h10 ;
			data[19373] <= 8'h10 ;
			data[19374] <= 8'h10 ;
			data[19375] <= 8'h10 ;
			data[19376] <= 8'h10 ;
			data[19377] <= 8'h10 ;
			data[19378] <= 8'h10 ;
			data[19379] <= 8'h10 ;
			data[19380] <= 8'h10 ;
			data[19381] <= 8'h10 ;
			data[19382] <= 8'h10 ;
			data[19383] <= 8'h10 ;
			data[19384] <= 8'h10 ;
			data[19385] <= 8'h10 ;
			data[19386] <= 8'h10 ;
			data[19387] <= 8'h10 ;
			data[19388] <= 8'h10 ;
			data[19389] <= 8'h10 ;
			data[19390] <= 8'h10 ;
			data[19391] <= 8'h10 ;
			data[19392] <= 8'h10 ;
			data[19393] <= 8'h10 ;
			data[19394] <= 8'h10 ;
			data[19395] <= 8'h10 ;
			data[19396] <= 8'h10 ;
			data[19397] <= 8'h10 ;
			data[19398] <= 8'h10 ;
			data[19399] <= 8'h10 ;
			data[19400] <= 8'h10 ;
			data[19401] <= 8'h10 ;
			data[19402] <= 8'h10 ;
			data[19403] <= 8'h10 ;
			data[19404] <= 8'h10 ;
			data[19405] <= 8'h10 ;
			data[19406] <= 8'h10 ;
			data[19407] <= 8'h10 ;
			data[19408] <= 8'h10 ;
			data[19409] <= 8'h10 ;
			data[19410] <= 8'h10 ;
			data[19411] <= 8'h10 ;
			data[19412] <= 8'h10 ;
			data[19413] <= 8'h10 ;
			data[19414] <= 8'h10 ;
			data[19415] <= 8'h10 ;
			data[19416] <= 8'h10 ;
			data[19417] <= 8'h10 ;
			data[19418] <= 8'h10 ;
			data[19419] <= 8'h10 ;
			data[19420] <= 8'h10 ;
			data[19421] <= 8'h10 ;
			data[19422] <= 8'h10 ;
			data[19423] <= 8'h10 ;
			data[19424] <= 8'h10 ;
			data[19425] <= 8'h10 ;
			data[19426] <= 8'h10 ;
			data[19427] <= 8'h10 ;
			data[19428] <= 8'h10 ;
			data[19429] <= 8'h10 ;
			data[19430] <= 8'h10 ;
			data[19431] <= 8'h10 ;
			data[19432] <= 8'h10 ;
			data[19433] <= 8'h10 ;
			data[19434] <= 8'h10 ;
			data[19435] <= 8'h10 ;
			data[19436] <= 8'h10 ;
			data[19437] <= 8'h10 ;
			data[19438] <= 8'h10 ;
			data[19439] <= 8'h10 ;
			data[19440] <= 8'h10 ;
			data[19441] <= 8'h10 ;
			data[19442] <= 8'h10 ;
			data[19443] <= 8'h10 ;
			data[19444] <= 8'h10 ;
			data[19445] <= 8'h10 ;
			data[19446] <= 8'h10 ;
			data[19447] <= 8'h10 ;
			data[19448] <= 8'h10 ;
			data[19449] <= 8'h10 ;
			data[19450] <= 8'h10 ;
			data[19451] <= 8'h10 ;
			data[19452] <= 8'h10 ;
			data[19453] <= 8'h10 ;
			data[19454] <= 8'h10 ;
			data[19455] <= 8'h10 ;
			data[19456] <= 8'h10 ;
			data[19457] <= 8'h10 ;
			data[19458] <= 8'h10 ;
			data[19459] <= 8'h10 ;
			data[19460] <= 8'h10 ;
			data[19461] <= 8'h10 ;
			data[19462] <= 8'h10 ;
			data[19463] <= 8'h10 ;
			data[19464] <= 8'h10 ;
			data[19465] <= 8'h10 ;
			data[19466] <= 8'h10 ;
			data[19467] <= 8'h10 ;
			data[19468] <= 8'h10 ;
			data[19469] <= 8'h10 ;
			data[19470] <= 8'h10 ;
			data[19471] <= 8'h10 ;
			data[19472] <= 8'h10 ;
			data[19473] <= 8'h10 ;
			data[19474] <= 8'h10 ;
			data[19475] <= 8'h10 ;
			data[19476] <= 8'h10 ;
			data[19477] <= 8'h10 ;
			data[19478] <= 8'h10 ;
			data[19479] <= 8'h10 ;
			data[19480] <= 8'h10 ;
			data[19481] <= 8'h10 ;
			data[19482] <= 8'h10 ;
			data[19483] <= 8'h10 ;
			data[19484] <= 8'h10 ;
			data[19485] <= 8'h10 ;
			data[19486] <= 8'h10 ;
			data[19487] <= 8'h10 ;
			data[19488] <= 8'h10 ;
			data[19489] <= 8'h10 ;
			data[19490] <= 8'h10 ;
			data[19491] <= 8'h10 ;
			data[19492] <= 8'h10 ;
			data[19493] <= 8'h10 ;
			data[19494] <= 8'h10 ;
			data[19495] <= 8'h10 ;
			data[19496] <= 8'h10 ;
			data[19497] <= 8'h10 ;
			data[19498] <= 8'h10 ;
			data[19499] <= 8'h10 ;
			data[19500] <= 8'h10 ;
			data[19501] <= 8'h10 ;
			data[19502] <= 8'h10 ;
			data[19503] <= 8'h10 ;
			data[19504] <= 8'h10 ;
			data[19505] <= 8'h10 ;
			data[19506] <= 8'h10 ;
			data[19507] <= 8'h10 ;
			data[19508] <= 8'h10 ;
			data[19509] <= 8'h10 ;
			data[19510] <= 8'h10 ;
			data[19511] <= 8'h10 ;
			data[19512] <= 8'h10 ;
			data[19513] <= 8'h10 ;
			data[19514] <= 8'h10 ;
			data[19515] <= 8'h10 ;
			data[19516] <= 8'h10 ;
			data[19517] <= 8'h10 ;
			data[19518] <= 8'h10 ;
			data[19519] <= 8'h10 ;
			data[19520] <= 8'h10 ;
			data[19521] <= 8'h10 ;
			data[19522] <= 8'h10 ;
			data[19523] <= 8'h10 ;
			data[19524] <= 8'h10 ;
			data[19525] <= 8'h10 ;
			data[19526] <= 8'h10 ;
			data[19527] <= 8'h10 ;
			data[19528] <= 8'h10 ;
			data[19529] <= 8'h10 ;
			data[19530] <= 8'h10 ;
			data[19531] <= 8'h10 ;
			data[19532] <= 8'h10 ;
			data[19533] <= 8'h10 ;
			data[19534] <= 8'h10 ;
			data[19535] <= 8'h10 ;
			data[19536] <= 8'h10 ;
			data[19537] <= 8'h10 ;
			data[19538] <= 8'h10 ;
			data[19539] <= 8'h10 ;
			data[19540] <= 8'h10 ;
			data[19541] <= 8'h10 ;
			data[19542] <= 8'h10 ;
			data[19543] <= 8'h10 ;
			data[19544] <= 8'h10 ;
			data[19545] <= 8'h10 ;
			data[19546] <= 8'h10 ;
			data[19547] <= 8'h10 ;
			data[19548] <= 8'h10 ;
			data[19549] <= 8'h10 ;
			data[19550] <= 8'h10 ;
			data[19551] <= 8'h10 ;
			data[19552] <= 8'h10 ;
			data[19553] <= 8'h10 ;
			data[19554] <= 8'h10 ;
			data[19555] <= 8'h10 ;
			data[19556] <= 8'h10 ;
			data[19557] <= 8'h10 ;
			data[19558] <= 8'h10 ;
			data[19559] <= 8'h10 ;
			data[19560] <= 8'h10 ;
			data[19561] <= 8'h10 ;
			data[19562] <= 8'h10 ;
			data[19563] <= 8'h10 ;
			data[19564] <= 8'h10 ;
			data[19565] <= 8'h10 ;
			data[19566] <= 8'h10 ;
			data[19567] <= 8'h10 ;
			data[19568] <= 8'h10 ;
			data[19569] <= 8'h10 ;
			data[19570] <= 8'h10 ;
			data[19571] <= 8'h10 ;
			data[19572] <= 8'h10 ;
			data[19573] <= 8'h10 ;
			data[19574] <= 8'h10 ;
			data[19575] <= 8'h10 ;
			data[19576] <= 8'h10 ;
			data[19577] <= 8'h10 ;
			data[19578] <= 8'h10 ;
			data[19579] <= 8'h10 ;
			data[19580] <= 8'h10 ;
			data[19581] <= 8'h10 ;
			data[19582] <= 8'h10 ;
			data[19583] <= 8'h10 ;
			data[19584] <= 8'h10 ;
			data[19585] <= 8'h10 ;
			data[19586] <= 8'h10 ;
			data[19587] <= 8'h10 ;
			data[19588] <= 8'h10 ;
			data[19589] <= 8'h10 ;
			data[19590] <= 8'h10 ;
			data[19591] <= 8'h10 ;
			data[19592] <= 8'h10 ;
			data[19593] <= 8'h10 ;
			data[19594] <= 8'h10 ;
			data[19595] <= 8'h10 ;
			data[19596] <= 8'h10 ;
			data[19597] <= 8'h10 ;
			data[19598] <= 8'h10 ;
			data[19599] <= 8'h10 ;
			data[19600] <= 8'h10 ;
			data[19601] <= 8'h10 ;
			data[19602] <= 8'h10 ;
			data[19603] <= 8'h10 ;
			data[19604] <= 8'h10 ;
			data[19605] <= 8'h10 ;
			data[19606] <= 8'h10 ;
			data[19607] <= 8'h10 ;
			data[19608] <= 8'h10 ;
			data[19609] <= 8'h10 ;
			data[19610] <= 8'h10 ;
			data[19611] <= 8'h10 ;
			data[19612] <= 8'h10 ;
			data[19613] <= 8'h10 ;
			data[19614] <= 8'h10 ;
			data[19615] <= 8'h10 ;
			data[19616] <= 8'h10 ;
			data[19617] <= 8'h10 ;
			data[19618] <= 8'h10 ;
			data[19619] <= 8'h10 ;
			data[19620] <= 8'h10 ;
			data[19621] <= 8'h10 ;
			data[19622] <= 8'h10 ;
			data[19623] <= 8'h10 ;
			data[19624] <= 8'h10 ;
			data[19625] <= 8'h10 ;
			data[19626] <= 8'h10 ;
			data[19627] <= 8'h10 ;
			data[19628] <= 8'h10 ;
			data[19629] <= 8'h10 ;
			data[19630] <= 8'h10 ;
			data[19631] <= 8'h10 ;
			data[19632] <= 8'h10 ;
			data[19633] <= 8'h10 ;
			data[19634] <= 8'h10 ;
			data[19635] <= 8'h10 ;
			data[19636] <= 8'h10 ;
			data[19637] <= 8'h10 ;
			data[19638] <= 8'h10 ;
			data[19639] <= 8'h10 ;
			data[19640] <= 8'h10 ;
			data[19641] <= 8'h10 ;
			data[19642] <= 8'h10 ;
			data[19643] <= 8'h10 ;
			data[19644] <= 8'h10 ;
			data[19645] <= 8'h10 ;
			data[19646] <= 8'h10 ;
			data[19647] <= 8'h10 ;
			data[19648] <= 8'h10 ;
			data[19649] <= 8'h10 ;
			data[19650] <= 8'h10 ;
			data[19651] <= 8'h10 ;
			data[19652] <= 8'h10 ;
			data[19653] <= 8'h10 ;
			data[19654] <= 8'h10 ;
			data[19655] <= 8'h10 ;
			data[19656] <= 8'h10 ;
			data[19657] <= 8'h10 ;
			data[19658] <= 8'h10 ;
			data[19659] <= 8'h10 ;
			data[19660] <= 8'h10 ;
			data[19661] <= 8'h10 ;
			data[19662] <= 8'h10 ;
			data[19663] <= 8'h10 ;
			data[19664] <= 8'h10 ;
			data[19665] <= 8'h10 ;
			data[19666] <= 8'h10 ;
			data[19667] <= 8'h10 ;
			data[19668] <= 8'h10 ;
			data[19669] <= 8'h10 ;
			data[19670] <= 8'h10 ;
			data[19671] <= 8'h10 ;
			data[19672] <= 8'h10 ;
			data[19673] <= 8'h10 ;
			data[19674] <= 8'h10 ;
			data[19675] <= 8'h10 ;
			data[19676] <= 8'h10 ;
			data[19677] <= 8'h10 ;
			data[19678] <= 8'h10 ;
			data[19679] <= 8'h10 ;
			data[19680] <= 8'h10 ;
			data[19681] <= 8'h10 ;
			data[19682] <= 8'h10 ;
			data[19683] <= 8'h10 ;
			data[19684] <= 8'h10 ;
			data[19685] <= 8'h10 ;
			data[19686] <= 8'h10 ;
			data[19687] <= 8'h10 ;
			data[19688] <= 8'h10 ;
			data[19689] <= 8'h10 ;
			data[19690] <= 8'h10 ;
			data[19691] <= 8'h10 ;
			data[19692] <= 8'h10 ;
			data[19693] <= 8'h10 ;
			data[19694] <= 8'h10 ;
			data[19695] <= 8'h10 ;
			data[19696] <= 8'h10 ;
			data[19697] <= 8'h10 ;
			data[19698] <= 8'h10 ;
			data[19699] <= 8'h10 ;
			data[19700] <= 8'h10 ;
			data[19701] <= 8'h10 ;
			data[19702] <= 8'h10 ;
			data[19703] <= 8'h10 ;
			data[19704] <= 8'h10 ;
			data[19705] <= 8'h10 ;
			data[19706] <= 8'h10 ;
			data[19707] <= 8'h10 ;
			data[19708] <= 8'h10 ;
			data[19709] <= 8'h10 ;
			data[19710] <= 8'h10 ;
			data[19711] <= 8'h10 ;
			data[19712] <= 8'h10 ;
			data[19713] <= 8'h10 ;
			data[19714] <= 8'h10 ;
			data[19715] <= 8'h10 ;
			data[19716] <= 8'h10 ;
			data[19717] <= 8'h10 ;
			data[19718] <= 8'h10 ;
			data[19719] <= 8'h10 ;
			data[19720] <= 8'h10 ;
			data[19721] <= 8'h10 ;
			data[19722] <= 8'h10 ;
			data[19723] <= 8'h10 ;
			data[19724] <= 8'h10 ;
			data[19725] <= 8'h10 ;
			data[19726] <= 8'h10 ;
			data[19727] <= 8'h10 ;
			data[19728] <= 8'h10 ;
			data[19729] <= 8'h10 ;
			data[19730] <= 8'h10 ;
			data[19731] <= 8'h10 ;
			data[19732] <= 8'h10 ;
			data[19733] <= 8'h10 ;
			data[19734] <= 8'h10 ;
			data[19735] <= 8'h10 ;
			data[19736] <= 8'h10 ;
			data[19737] <= 8'h10 ;
			data[19738] <= 8'h10 ;
			data[19739] <= 8'h10 ;
			data[19740] <= 8'h10 ;
			data[19741] <= 8'h10 ;
			data[19742] <= 8'h10 ;
			data[19743] <= 8'h10 ;
			data[19744] <= 8'h10 ;
			data[19745] <= 8'h10 ;
			data[19746] <= 8'h10 ;
			data[19747] <= 8'h10 ;
			data[19748] <= 8'h10 ;
			data[19749] <= 8'h10 ;
			data[19750] <= 8'h10 ;
			data[19751] <= 8'h10 ;
			data[19752] <= 8'h10 ;
			data[19753] <= 8'h10 ;
			data[19754] <= 8'h10 ;
			data[19755] <= 8'h10 ;
			data[19756] <= 8'h10 ;
			data[19757] <= 8'h10 ;
			data[19758] <= 8'h10 ;
			data[19759] <= 8'h10 ;
			data[19760] <= 8'h10 ;
			data[19761] <= 8'h10 ;
			data[19762] <= 8'h10 ;
			data[19763] <= 8'h10 ;
			data[19764] <= 8'h10 ;
			data[19765] <= 8'h10 ;
			data[19766] <= 8'h10 ;
			data[19767] <= 8'h10 ;
			data[19768] <= 8'h10 ;
			data[19769] <= 8'h10 ;
			data[19770] <= 8'h10 ;
			data[19771] <= 8'h10 ;
			data[19772] <= 8'h10 ;
			data[19773] <= 8'h10 ;
			data[19774] <= 8'h10 ;
			data[19775] <= 8'h10 ;
			data[19776] <= 8'h10 ;
			data[19777] <= 8'h10 ;
			data[19778] <= 8'h10 ;
			data[19779] <= 8'h10 ;
			data[19780] <= 8'h10 ;
			data[19781] <= 8'h10 ;
			data[19782] <= 8'h10 ;
			data[19783] <= 8'h10 ;
			data[19784] <= 8'h10 ;
			data[19785] <= 8'h10 ;
			data[19786] <= 8'h10 ;
			data[19787] <= 8'h10 ;
			data[19788] <= 8'h10 ;
			data[19789] <= 8'h10 ;
			data[19790] <= 8'h10 ;
			data[19791] <= 8'h10 ;
			data[19792] <= 8'h10 ;
			data[19793] <= 8'h10 ;
			data[19794] <= 8'h10 ;
			data[19795] <= 8'h10 ;
			data[19796] <= 8'h10 ;
			data[19797] <= 8'h10 ;
			data[19798] <= 8'h10 ;
			data[19799] <= 8'h10 ;
			data[19800] <= 8'h10 ;
			data[19801] <= 8'h10 ;
			data[19802] <= 8'h10 ;
			data[19803] <= 8'h10 ;
			data[19804] <= 8'h10 ;
			data[19805] <= 8'h10 ;
			data[19806] <= 8'h10 ;
			data[19807] <= 8'h10 ;
			data[19808] <= 8'h10 ;
			data[19809] <= 8'h10 ;
			data[19810] <= 8'h10 ;
			data[19811] <= 8'h10 ;
			data[19812] <= 8'h10 ;
			data[19813] <= 8'h10 ;
			data[19814] <= 8'h10 ;
			data[19815] <= 8'h10 ;
			data[19816] <= 8'h10 ;
			data[19817] <= 8'h10 ;
			data[19818] <= 8'h10 ;
			data[19819] <= 8'h10 ;
			data[19820] <= 8'h10 ;
			data[19821] <= 8'h10 ;
			data[19822] <= 8'h10 ;
			data[19823] <= 8'h10 ;
			data[19824] <= 8'h10 ;
			data[19825] <= 8'h10 ;
			data[19826] <= 8'h10 ;
			data[19827] <= 8'h10 ;
			data[19828] <= 8'h10 ;
			data[19829] <= 8'h10 ;
			data[19830] <= 8'h10 ;
			data[19831] <= 8'h10 ;
			data[19832] <= 8'h10 ;
			data[19833] <= 8'h10 ;
			data[19834] <= 8'h10 ;
			data[19835] <= 8'h10 ;
			data[19836] <= 8'h10 ;
			data[19837] <= 8'h10 ;
			data[19838] <= 8'h10 ;
			data[19839] <= 8'h10 ;
			data[19840] <= 8'h10 ;
			data[19841] <= 8'h10 ;
			data[19842] <= 8'h10 ;
			data[19843] <= 8'h10 ;
			data[19844] <= 8'h10 ;
			data[19845] <= 8'h10 ;
			data[19846] <= 8'h10 ;
			data[19847] <= 8'h10 ;
			data[19848] <= 8'h10 ;
			data[19849] <= 8'h10 ;
			data[19850] <= 8'h10 ;
			data[19851] <= 8'h10 ;
			data[19852] <= 8'h10 ;
			data[19853] <= 8'h10 ;
			data[19854] <= 8'h10 ;
			data[19855] <= 8'h10 ;
			data[19856] <= 8'h10 ;
			data[19857] <= 8'h10 ;
			data[19858] <= 8'h10 ;
			data[19859] <= 8'h10 ;
			data[19860] <= 8'h10 ;
			data[19861] <= 8'h10 ;
			data[19862] <= 8'h10 ;
			data[19863] <= 8'h10 ;
			data[19864] <= 8'h10 ;
			data[19865] <= 8'h10 ;
			data[19866] <= 8'h10 ;
			data[19867] <= 8'h10 ;
			data[19868] <= 8'h10 ;
			data[19869] <= 8'h10 ;
			data[19870] <= 8'h10 ;
			data[19871] <= 8'h10 ;
			data[19872] <= 8'h10 ;
			data[19873] <= 8'h10 ;
			data[19874] <= 8'h10 ;
			data[19875] <= 8'h10 ;
			data[19876] <= 8'h10 ;
			data[19877] <= 8'h10 ;
			data[19878] <= 8'h10 ;
			data[19879] <= 8'h10 ;
			data[19880] <= 8'h10 ;
			data[19881] <= 8'h10 ;
			data[19882] <= 8'h10 ;
			data[19883] <= 8'h10 ;
			data[19884] <= 8'h10 ;
			data[19885] <= 8'h10 ;
			data[19886] <= 8'h10 ;
			data[19887] <= 8'h10 ;
			data[19888] <= 8'h10 ;
			data[19889] <= 8'h10 ;
			data[19890] <= 8'h10 ;
			data[19891] <= 8'h10 ;
			data[19892] <= 8'h10 ;
			data[19893] <= 8'h10 ;
			data[19894] <= 8'h10 ;
			data[19895] <= 8'h10 ;
			data[19896] <= 8'h10 ;
			data[19897] <= 8'h10 ;
			data[19898] <= 8'h10 ;
			data[19899] <= 8'h10 ;
			data[19900] <= 8'h10 ;
			data[19901] <= 8'h10 ;
			data[19902] <= 8'h10 ;
			data[19903] <= 8'h10 ;
			data[19904] <= 8'h10 ;
			data[19905] <= 8'h10 ;
			data[19906] <= 8'h10 ;
			data[19907] <= 8'h10 ;
			data[19908] <= 8'h10 ;
			data[19909] <= 8'h10 ;
			data[19910] <= 8'h10 ;
			data[19911] <= 8'h10 ;
			data[19912] <= 8'h10 ;
			data[19913] <= 8'h10 ;
			data[19914] <= 8'h10 ;
			data[19915] <= 8'h10 ;
			data[19916] <= 8'h10 ;
			data[19917] <= 8'h10 ;
			data[19918] <= 8'h10 ;
			data[19919] <= 8'h10 ;
			data[19920] <= 8'h10 ;
			data[19921] <= 8'h10 ;
			data[19922] <= 8'h10 ;
			data[19923] <= 8'h10 ;
			data[19924] <= 8'h10 ;
			data[19925] <= 8'h10 ;
			data[19926] <= 8'h10 ;
			data[19927] <= 8'h10 ;
			data[19928] <= 8'h10 ;
			data[19929] <= 8'h10 ;
			data[19930] <= 8'h10 ;
			data[19931] <= 8'h10 ;
			data[19932] <= 8'h10 ;
			data[19933] <= 8'h10 ;
			data[19934] <= 8'h10 ;
			data[19935] <= 8'h10 ;
			data[19936] <= 8'h10 ;
			data[19937] <= 8'h10 ;
			data[19938] <= 8'h10 ;
			data[19939] <= 8'h10 ;
			data[19940] <= 8'h10 ;
			data[19941] <= 8'h10 ;
			data[19942] <= 8'h10 ;
			data[19943] <= 8'h10 ;
			data[19944] <= 8'h10 ;
			data[19945] <= 8'h10 ;
			data[19946] <= 8'h10 ;
			data[19947] <= 8'h10 ;
			data[19948] <= 8'h10 ;
			data[19949] <= 8'h10 ;
			data[19950] <= 8'h10 ;
			data[19951] <= 8'h10 ;
			data[19952] <= 8'h10 ;
			data[19953] <= 8'h10 ;
			data[19954] <= 8'h10 ;
			data[19955] <= 8'h10 ;
			data[19956] <= 8'h10 ;
			data[19957] <= 8'h10 ;
			data[19958] <= 8'h10 ;
			data[19959] <= 8'h10 ;
			data[19960] <= 8'h10 ;
			data[19961] <= 8'h10 ;
			data[19962] <= 8'h10 ;
			data[19963] <= 8'h10 ;
			data[19964] <= 8'h10 ;
			data[19965] <= 8'h10 ;
			data[19966] <= 8'h10 ;
			data[19967] <= 8'h10 ;
			data[19968] <= 8'h10 ;
			data[19969] <= 8'h10 ;
			data[19970] <= 8'h10 ;
			data[19971] <= 8'h10 ;
			data[19972] <= 8'h10 ;
			data[19973] <= 8'h10 ;
			data[19974] <= 8'h10 ;
			data[19975] <= 8'h10 ;
			data[19976] <= 8'h10 ;
			data[19977] <= 8'h10 ;
			data[19978] <= 8'h10 ;
			data[19979] <= 8'h10 ;
			data[19980] <= 8'h10 ;
			data[19981] <= 8'h10 ;
			data[19982] <= 8'h10 ;
			data[19983] <= 8'h10 ;
			data[19984] <= 8'h10 ;
			data[19985] <= 8'h10 ;
			data[19986] <= 8'h10 ;
			data[19987] <= 8'h10 ;
			data[19988] <= 8'h10 ;
			data[19989] <= 8'h10 ;
			data[19990] <= 8'h10 ;
			data[19991] <= 8'h10 ;
			data[19992] <= 8'h10 ;
			data[19993] <= 8'h10 ;
			data[19994] <= 8'h10 ;
			data[19995] <= 8'h10 ;
			data[19996] <= 8'h10 ;
			data[19997] <= 8'h10 ;
			data[19998] <= 8'h10 ;
			data[19999] <= 8'h10 ;
			data[20000] <= 8'h10 ;
			data[20001] <= 8'h10 ;
			data[20002] <= 8'h10 ;
			data[20003] <= 8'h10 ;
			data[20004] <= 8'h10 ;
			data[20005] <= 8'h10 ;
			data[20006] <= 8'h10 ;
			data[20007] <= 8'h10 ;
			data[20008] <= 8'h10 ;
			data[20009] <= 8'h10 ;
			data[20010] <= 8'h10 ;
			data[20011] <= 8'h10 ;
			data[20012] <= 8'h10 ;
			data[20013] <= 8'h10 ;
			data[20014] <= 8'h10 ;
			data[20015] <= 8'h10 ;
			data[20016] <= 8'h10 ;
			data[20017] <= 8'h10 ;
			data[20018] <= 8'h10 ;
			data[20019] <= 8'h10 ;
			data[20020] <= 8'h10 ;
			data[20021] <= 8'h10 ;
			data[20022] <= 8'h10 ;
			data[20023] <= 8'h10 ;
			data[20024] <= 8'h10 ;
			data[20025] <= 8'h10 ;
			data[20026] <= 8'h10 ;
			data[20027] <= 8'h10 ;
			data[20028] <= 8'h10 ;
			data[20029] <= 8'h10 ;
			data[20030] <= 8'h10 ;
			data[20031] <= 8'h10 ;
			data[20032] <= 8'h10 ;
			data[20033] <= 8'h10 ;
			data[20034] <= 8'h10 ;
			data[20035] <= 8'h10 ;
			data[20036] <= 8'h10 ;
			data[20037] <= 8'h10 ;
			data[20038] <= 8'h10 ;
			data[20039] <= 8'h10 ;
			data[20040] <= 8'h10 ;
			data[20041] <= 8'h10 ;
			data[20042] <= 8'h10 ;
			data[20043] <= 8'h10 ;
			data[20044] <= 8'h10 ;
			data[20045] <= 8'h10 ;
			data[20046] <= 8'h10 ;
			data[20047] <= 8'h10 ;
			data[20048] <= 8'h10 ;
			data[20049] <= 8'h10 ;
			data[20050] <= 8'h10 ;
			data[20051] <= 8'h10 ;
			data[20052] <= 8'h10 ;
			data[20053] <= 8'h10 ;
			data[20054] <= 8'h10 ;
			data[20055] <= 8'h10 ;
			data[20056] <= 8'h10 ;
			data[20057] <= 8'h10 ;
			data[20058] <= 8'h10 ;
			data[20059] <= 8'h10 ;
			data[20060] <= 8'h10 ;
			data[20061] <= 8'h10 ;
			data[20062] <= 8'h10 ;
			data[20063] <= 8'h10 ;
			data[20064] <= 8'h10 ;
			data[20065] <= 8'h10 ;
			data[20066] <= 8'h10 ;
			data[20067] <= 8'h10 ;
			data[20068] <= 8'h10 ;
			data[20069] <= 8'h10 ;
			data[20070] <= 8'h10 ;
			data[20071] <= 8'h10 ;
			data[20072] <= 8'h10 ;
			data[20073] <= 8'h10 ;
			data[20074] <= 8'h10 ;
			data[20075] <= 8'h10 ;
			data[20076] <= 8'h10 ;
			data[20077] <= 8'h10 ;
			data[20078] <= 8'h10 ;
			data[20079] <= 8'h10 ;
			data[20080] <= 8'h10 ;
			data[20081] <= 8'h10 ;
			data[20082] <= 8'h10 ;
			data[20083] <= 8'h10 ;
			data[20084] <= 8'h10 ;
			data[20085] <= 8'h10 ;
			data[20086] <= 8'h10 ;
			data[20087] <= 8'h10 ;
			data[20088] <= 8'h10 ;
			data[20089] <= 8'h10 ;
			data[20090] <= 8'h10 ;
			data[20091] <= 8'h10 ;
			data[20092] <= 8'h10 ;
			data[20093] <= 8'h10 ;
			data[20094] <= 8'h10 ;
			data[20095] <= 8'h10 ;
			data[20096] <= 8'h10 ;
			data[20097] <= 8'h10 ;
			data[20098] <= 8'h10 ;
			data[20099] <= 8'h10 ;
			data[20100] <= 8'h10 ;
			data[20101] <= 8'h10 ;
			data[20102] <= 8'h10 ;
			data[20103] <= 8'h10 ;
			data[20104] <= 8'h10 ;
			data[20105] <= 8'h10 ;
			data[20106] <= 8'h10 ;
			data[20107] <= 8'h10 ;
			data[20108] <= 8'h10 ;
			data[20109] <= 8'h10 ;
			data[20110] <= 8'h10 ;
			data[20111] <= 8'h10 ;
			data[20112] <= 8'h10 ;
			data[20113] <= 8'h10 ;
			data[20114] <= 8'h10 ;
			data[20115] <= 8'h10 ;
			data[20116] <= 8'h10 ;
			data[20117] <= 8'h10 ;
			data[20118] <= 8'h10 ;
			data[20119] <= 8'h10 ;
			data[20120] <= 8'h10 ;
			data[20121] <= 8'h10 ;
			data[20122] <= 8'h10 ;
			data[20123] <= 8'h10 ;
			data[20124] <= 8'h10 ;
			data[20125] <= 8'h10 ;
			data[20126] <= 8'h10 ;
			data[20127] <= 8'h10 ;
			data[20128] <= 8'h10 ;
			data[20129] <= 8'h10 ;
			data[20130] <= 8'h10 ;
			data[20131] <= 8'h10 ;
			data[20132] <= 8'h10 ;
			data[20133] <= 8'h10 ;
			data[20134] <= 8'h10 ;
			data[20135] <= 8'h10 ;
			data[20136] <= 8'h10 ;
			data[20137] <= 8'h10 ;
			data[20138] <= 8'h10 ;
			data[20139] <= 8'h10 ;
			data[20140] <= 8'h10 ;
			data[20141] <= 8'h10 ;
			data[20142] <= 8'h10 ;
			data[20143] <= 8'h10 ;
			data[20144] <= 8'h10 ;
			data[20145] <= 8'h10 ;
			data[20146] <= 8'h10 ;
			data[20147] <= 8'h10 ;
			data[20148] <= 8'h10 ;
			data[20149] <= 8'h10 ;
			data[20150] <= 8'h10 ;
			data[20151] <= 8'h10 ;
			data[20152] <= 8'h10 ;
			data[20153] <= 8'h10 ;
			data[20154] <= 8'h10 ;
			data[20155] <= 8'h10 ;
			data[20156] <= 8'h10 ;
			data[20157] <= 8'h10 ;
			data[20158] <= 8'h10 ;
			data[20159] <= 8'h10 ;
			data[20160] <= 8'h10 ;
			data[20161] <= 8'h10 ;
			data[20162] <= 8'h10 ;
			data[20163] <= 8'h10 ;
			data[20164] <= 8'h10 ;
			data[20165] <= 8'h10 ;
			data[20166] <= 8'h10 ;
			data[20167] <= 8'h10 ;
			data[20168] <= 8'h10 ;
			data[20169] <= 8'h10 ;
			data[20170] <= 8'h10 ;
			data[20171] <= 8'h10 ;
			data[20172] <= 8'h10 ;
			data[20173] <= 8'h10 ;
			data[20174] <= 8'h10 ;
			data[20175] <= 8'h10 ;
			data[20176] <= 8'h10 ;
			data[20177] <= 8'h10 ;
			data[20178] <= 8'h10 ;
			data[20179] <= 8'h10 ;
			data[20180] <= 8'h10 ;
			data[20181] <= 8'h10 ;
			data[20182] <= 8'h10 ;
			data[20183] <= 8'h10 ;
			data[20184] <= 8'h10 ;
			data[20185] <= 8'h10 ;
			data[20186] <= 8'h10 ;
			data[20187] <= 8'h10 ;
			data[20188] <= 8'h10 ;
			data[20189] <= 8'h10 ;
			data[20190] <= 8'h10 ;
			data[20191] <= 8'h10 ;
			data[20192] <= 8'h10 ;
			data[20193] <= 8'h10 ;
			data[20194] <= 8'h10 ;
			data[20195] <= 8'h10 ;
			data[20196] <= 8'h10 ;
			data[20197] <= 8'h10 ;
			data[20198] <= 8'h10 ;
			data[20199] <= 8'h10 ;
			data[20200] <= 8'h10 ;
			data[20201] <= 8'h10 ;
			data[20202] <= 8'h10 ;
			data[20203] <= 8'h10 ;
			data[20204] <= 8'h10 ;
			data[20205] <= 8'h10 ;
			data[20206] <= 8'h10 ;
			data[20207] <= 8'h10 ;
			data[20208] <= 8'h10 ;
			data[20209] <= 8'h10 ;
			data[20210] <= 8'h10 ;
			data[20211] <= 8'h10 ;
			data[20212] <= 8'h10 ;
			data[20213] <= 8'h10 ;
			data[20214] <= 8'h10 ;
			data[20215] <= 8'h10 ;
			data[20216] <= 8'h10 ;
			data[20217] <= 8'h10 ;
			data[20218] <= 8'h10 ;
			data[20219] <= 8'h10 ;
			data[20220] <= 8'h10 ;
			data[20221] <= 8'h10 ;
			data[20222] <= 8'h10 ;
			data[20223] <= 8'h10 ;
			data[20224] <= 8'h10 ;
			data[20225] <= 8'h10 ;
			data[20226] <= 8'h10 ;
			data[20227] <= 8'h10 ;
			data[20228] <= 8'h10 ;
			data[20229] <= 8'h10 ;
			data[20230] <= 8'h10 ;
			data[20231] <= 8'h10 ;
			data[20232] <= 8'h10 ;
			data[20233] <= 8'h10 ;
			data[20234] <= 8'h10 ;
			data[20235] <= 8'h10 ;
			data[20236] <= 8'h10 ;
			data[20237] <= 8'h10 ;
			data[20238] <= 8'h10 ;
			data[20239] <= 8'h10 ;
			data[20240] <= 8'h10 ;
			data[20241] <= 8'h10 ;
			data[20242] <= 8'h10 ;
			data[20243] <= 8'h10 ;
			data[20244] <= 8'h10 ;
			data[20245] <= 8'h10 ;
			data[20246] <= 8'h10 ;
			data[20247] <= 8'h10 ;
			data[20248] <= 8'h10 ;
			data[20249] <= 8'h10 ;
			data[20250] <= 8'h10 ;
			data[20251] <= 8'h10 ;
			data[20252] <= 8'h10 ;
			data[20253] <= 8'h10 ;
			data[20254] <= 8'h10 ;
			data[20255] <= 8'h10 ;
			data[20256] <= 8'h10 ;
			data[20257] <= 8'h10 ;
			data[20258] <= 8'h10 ;
			data[20259] <= 8'h10 ;
			data[20260] <= 8'h10 ;
			data[20261] <= 8'h10 ;
			data[20262] <= 8'h10 ;
			data[20263] <= 8'h10 ;
			data[20264] <= 8'h10 ;
			data[20265] <= 8'h10 ;
			data[20266] <= 8'h10 ;
			data[20267] <= 8'h10 ;
			data[20268] <= 8'h10 ;
			data[20269] <= 8'h10 ;
			data[20270] <= 8'h10 ;
			data[20271] <= 8'h10 ;
			data[20272] <= 8'h10 ;
			data[20273] <= 8'h10 ;
			data[20274] <= 8'h10 ;
			data[20275] <= 8'h10 ;
			data[20276] <= 8'h10 ;
			data[20277] <= 8'h10 ;
			data[20278] <= 8'h10 ;
			data[20279] <= 8'h10 ;
			data[20280] <= 8'h10 ;
			data[20281] <= 8'h10 ;
			data[20282] <= 8'h10 ;
			data[20283] <= 8'h10 ;
			data[20284] <= 8'h10 ;
			data[20285] <= 8'h10 ;
			data[20286] <= 8'h10 ;
			data[20287] <= 8'h10 ;
			data[20288] <= 8'h10 ;
			data[20289] <= 8'h10 ;
			data[20290] <= 8'h10 ;
			data[20291] <= 8'h10 ;
			data[20292] <= 8'h10 ;
			data[20293] <= 8'h10 ;
			data[20294] <= 8'h10 ;
			data[20295] <= 8'h10 ;
			data[20296] <= 8'h10 ;
			data[20297] <= 8'h10 ;
			data[20298] <= 8'h10 ;
			data[20299] <= 8'h10 ;
			data[20300] <= 8'h10 ;
			data[20301] <= 8'h10 ;
			data[20302] <= 8'h10 ;
			data[20303] <= 8'h10 ;
			data[20304] <= 8'h10 ;
			data[20305] <= 8'h10 ;
			data[20306] <= 8'h10 ;
			data[20307] <= 8'h10 ;
			data[20308] <= 8'h10 ;
			data[20309] <= 8'h10 ;
			data[20310] <= 8'h10 ;
			data[20311] <= 8'h10 ;
			data[20312] <= 8'h10 ;
			data[20313] <= 8'h10 ;
			data[20314] <= 8'h10 ;
			data[20315] <= 8'h10 ;
			data[20316] <= 8'h10 ;
			data[20317] <= 8'h10 ;
			data[20318] <= 8'h10 ;
			data[20319] <= 8'h10 ;
			data[20320] <= 8'h10 ;
			data[20321] <= 8'h10 ;
			data[20322] <= 8'h10 ;
			data[20323] <= 8'h10 ;
			data[20324] <= 8'h10 ;
			data[20325] <= 8'h10 ;
			data[20326] <= 8'h10 ;
			data[20327] <= 8'h10 ;
			data[20328] <= 8'h10 ;
			data[20329] <= 8'h10 ;
			data[20330] <= 8'h10 ;
			data[20331] <= 8'h10 ;
			data[20332] <= 8'h10 ;
			data[20333] <= 8'h10 ;
			data[20334] <= 8'h10 ;
			data[20335] <= 8'h10 ;
			data[20336] <= 8'h10 ;
			data[20337] <= 8'h10 ;
			data[20338] <= 8'h10 ;
			data[20339] <= 8'h10 ;
			data[20340] <= 8'h10 ;
			data[20341] <= 8'h10 ;
			data[20342] <= 8'h10 ;
			data[20343] <= 8'h10 ;
			data[20344] <= 8'h10 ;
			data[20345] <= 8'h10 ;
			data[20346] <= 8'h10 ;
			data[20347] <= 8'h10 ;
			data[20348] <= 8'h10 ;
			data[20349] <= 8'h10 ;
			data[20350] <= 8'h10 ;
			data[20351] <= 8'h10 ;
			data[20352] <= 8'h10 ;
			data[20353] <= 8'h10 ;
			data[20354] <= 8'h10 ;
			data[20355] <= 8'h10 ;
			data[20356] <= 8'h10 ;
			data[20357] <= 8'h10 ;
			data[20358] <= 8'h10 ;
			data[20359] <= 8'h10 ;
			data[20360] <= 8'h10 ;
			data[20361] <= 8'h10 ;
			data[20362] <= 8'h10 ;
			data[20363] <= 8'h10 ;
			data[20364] <= 8'h10 ;
			data[20365] <= 8'h10 ;
			data[20366] <= 8'h10 ;
			data[20367] <= 8'h10 ;
			data[20368] <= 8'h10 ;
			data[20369] <= 8'h10 ;
			data[20370] <= 8'h10 ;
			data[20371] <= 8'h10 ;
			data[20372] <= 8'h10 ;
			data[20373] <= 8'h10 ;
			data[20374] <= 8'h10 ;
			data[20375] <= 8'h10 ;
			data[20376] <= 8'h10 ;
			data[20377] <= 8'h10 ;
			data[20378] <= 8'h10 ;
			data[20379] <= 8'h10 ;
			data[20380] <= 8'h10 ;
			data[20381] <= 8'h10 ;
			data[20382] <= 8'h10 ;
			data[20383] <= 8'h10 ;
			data[20384] <= 8'h10 ;
			data[20385] <= 8'h10 ;
			data[20386] <= 8'h10 ;
			data[20387] <= 8'h10 ;
			data[20388] <= 8'h10 ;
			data[20389] <= 8'h10 ;
			data[20390] <= 8'h10 ;
			data[20391] <= 8'h10 ;
			data[20392] <= 8'h10 ;
			data[20393] <= 8'h10 ;
			data[20394] <= 8'h10 ;
			data[20395] <= 8'h10 ;
			data[20396] <= 8'h10 ;
			data[20397] <= 8'h10 ;
			data[20398] <= 8'h10 ;
			data[20399] <= 8'h10 ;
			data[20400] <= 8'h10 ;
			data[20401] <= 8'h10 ;
			data[20402] <= 8'h10 ;
			data[20403] <= 8'h10 ;
			data[20404] <= 8'h10 ;
			data[20405] <= 8'h10 ;
			data[20406] <= 8'h10 ;
			data[20407] <= 8'h10 ;
			data[20408] <= 8'h10 ;
			data[20409] <= 8'h10 ;
			data[20410] <= 8'h10 ;
			data[20411] <= 8'h10 ;
			data[20412] <= 8'h10 ;
			data[20413] <= 8'h10 ;
			data[20414] <= 8'h10 ;
			data[20415] <= 8'h10 ;
			data[20416] <= 8'h10 ;
			data[20417] <= 8'h10 ;
			data[20418] <= 8'h10 ;
			data[20419] <= 8'h10 ;
			data[20420] <= 8'h10 ;
			data[20421] <= 8'h10 ;
			data[20422] <= 8'h10 ;
			data[20423] <= 8'h10 ;
			data[20424] <= 8'h10 ;
			data[20425] <= 8'h10 ;
			data[20426] <= 8'h10 ;
			data[20427] <= 8'h10 ;
			data[20428] <= 8'h10 ;
			data[20429] <= 8'h10 ;
			data[20430] <= 8'h10 ;
			data[20431] <= 8'h10 ;
			data[20432] <= 8'h10 ;
			data[20433] <= 8'h10 ;
			data[20434] <= 8'h10 ;
			data[20435] <= 8'h10 ;
			data[20436] <= 8'h10 ;
			data[20437] <= 8'h10 ;
			data[20438] <= 8'h10 ;
			data[20439] <= 8'h10 ;
			data[20440] <= 8'h10 ;
			data[20441] <= 8'h10 ;
			data[20442] <= 8'h10 ;
			data[20443] <= 8'h10 ;
			data[20444] <= 8'h10 ;
			data[20445] <= 8'h10 ;
			data[20446] <= 8'h10 ;
			data[20447] <= 8'h10 ;
			data[20448] <= 8'h10 ;
			data[20449] <= 8'h10 ;
			data[20450] <= 8'h10 ;
			data[20451] <= 8'h10 ;
			data[20452] <= 8'h10 ;
			data[20453] <= 8'h10 ;
			data[20454] <= 8'h10 ;
			data[20455] <= 8'h10 ;
			data[20456] <= 8'h10 ;
			data[20457] <= 8'h10 ;
			data[20458] <= 8'h10 ;
			data[20459] <= 8'h10 ;
			data[20460] <= 8'h10 ;
			data[20461] <= 8'h10 ;
			data[20462] <= 8'h10 ;
			data[20463] <= 8'h10 ;
			data[20464] <= 8'h10 ;
			data[20465] <= 8'h10 ;
			data[20466] <= 8'h10 ;
			data[20467] <= 8'h10 ;
			data[20468] <= 8'h10 ;
			data[20469] <= 8'h10 ;
			data[20470] <= 8'h10 ;
			data[20471] <= 8'h10 ;
			data[20472] <= 8'h10 ;
			data[20473] <= 8'h10 ;
			data[20474] <= 8'h10 ;
			data[20475] <= 8'h10 ;
			data[20476] <= 8'h10 ;
			data[20477] <= 8'h10 ;
			data[20478] <= 8'h10 ;
			data[20479] <= 8'h10 ;
			data[20480] <= 8'h10 ;
			data[20481] <= 8'h10 ;
			data[20482] <= 8'h10 ;
			data[20483] <= 8'h10 ;
			data[20484] <= 8'h10 ;
			data[20485] <= 8'h10 ;
			data[20486] <= 8'h10 ;
			data[20487] <= 8'h10 ;
			data[20488] <= 8'h10 ;
			data[20489] <= 8'h10 ;
			data[20490] <= 8'h10 ;
			data[20491] <= 8'h10 ;
			data[20492] <= 8'h10 ;
			data[20493] <= 8'h10 ;
			data[20494] <= 8'h10 ;
			data[20495] <= 8'h10 ;
			data[20496] <= 8'h10 ;
			data[20497] <= 8'h10 ;
			data[20498] <= 8'h10 ;
			data[20499] <= 8'h10 ;
			data[20500] <= 8'h10 ;
			data[20501] <= 8'h10 ;
			data[20502] <= 8'h10 ;
			data[20503] <= 8'h10 ;
			data[20504] <= 8'h10 ;
			data[20505] <= 8'h10 ;
			data[20506] <= 8'h10 ;
			data[20507] <= 8'h10 ;
			data[20508] <= 8'h10 ;
			data[20509] <= 8'h10 ;
			data[20510] <= 8'h10 ;
			data[20511] <= 8'h10 ;
			data[20512] <= 8'h10 ;
			data[20513] <= 8'h10 ;
			data[20514] <= 8'h10 ;
			data[20515] <= 8'h10 ;
			data[20516] <= 8'h10 ;
			data[20517] <= 8'h10 ;
			data[20518] <= 8'h10 ;
			data[20519] <= 8'h10 ;
			data[20520] <= 8'h10 ;
			data[20521] <= 8'h10 ;
			data[20522] <= 8'h10 ;
			data[20523] <= 8'h10 ;
			data[20524] <= 8'h10 ;
			data[20525] <= 8'h10 ;
			data[20526] <= 8'h10 ;
			data[20527] <= 8'h10 ;
			data[20528] <= 8'h10 ;
			data[20529] <= 8'h10 ;
			data[20530] <= 8'h10 ;
			data[20531] <= 8'h10 ;
			data[20532] <= 8'h10 ;
			data[20533] <= 8'h10 ;
			data[20534] <= 8'h10 ;
			data[20535] <= 8'h10 ;
			data[20536] <= 8'h10 ;
			data[20537] <= 8'h10 ;
			data[20538] <= 8'h10 ;
			data[20539] <= 8'h10 ;
			data[20540] <= 8'h10 ;
			data[20541] <= 8'h10 ;
			data[20542] <= 8'h10 ;
			data[20543] <= 8'h10 ;
			data[20544] <= 8'h10 ;
			data[20545] <= 8'h10 ;
			data[20546] <= 8'h10 ;
			data[20547] <= 8'h10 ;
			data[20548] <= 8'h10 ;
			data[20549] <= 8'h10 ;
			data[20550] <= 8'h10 ;
			data[20551] <= 8'h10 ;
			data[20552] <= 8'h10 ;
			data[20553] <= 8'h10 ;
			data[20554] <= 8'h10 ;
			data[20555] <= 8'h10 ;
			data[20556] <= 8'h10 ;
			data[20557] <= 8'h10 ;
			data[20558] <= 8'h10 ;
			data[20559] <= 8'h10 ;
			data[20560] <= 8'h10 ;
			data[20561] <= 8'h10 ;
			data[20562] <= 8'h10 ;
			data[20563] <= 8'h10 ;
			data[20564] <= 8'h10 ;
			data[20565] <= 8'h10 ;
			data[20566] <= 8'h10 ;
			data[20567] <= 8'h10 ;
			data[20568] <= 8'h10 ;
			data[20569] <= 8'h10 ;
			data[20570] <= 8'h10 ;
			data[20571] <= 8'h10 ;
			data[20572] <= 8'h10 ;
			data[20573] <= 8'h10 ;
			data[20574] <= 8'h10 ;
			data[20575] <= 8'h10 ;
			data[20576] <= 8'h10 ;
			data[20577] <= 8'h10 ;
			data[20578] <= 8'h10 ;
			data[20579] <= 8'h10 ;
			data[20580] <= 8'h10 ;
			data[20581] <= 8'h10 ;
			data[20582] <= 8'h10 ;
			data[20583] <= 8'h10 ;
			data[20584] <= 8'h10 ;
			data[20585] <= 8'h10 ;
			data[20586] <= 8'h10 ;
			data[20587] <= 8'h10 ;
			data[20588] <= 8'h10 ;
			data[20589] <= 8'h10 ;
			data[20590] <= 8'h10 ;
			data[20591] <= 8'h10 ;
			data[20592] <= 8'h10 ;
			data[20593] <= 8'h10 ;
			data[20594] <= 8'h10 ;
			data[20595] <= 8'h10 ;
			data[20596] <= 8'h10 ;
			data[20597] <= 8'h10 ;
			data[20598] <= 8'h10 ;
			data[20599] <= 8'h10 ;
			data[20600] <= 8'h10 ;
			data[20601] <= 8'h10 ;
			data[20602] <= 8'h10 ;
			data[20603] <= 8'h10 ;
			data[20604] <= 8'h10 ;
			data[20605] <= 8'h10 ;
			data[20606] <= 8'h10 ;
			data[20607] <= 8'h10 ;
			data[20608] <= 8'h10 ;
			data[20609] <= 8'h10 ;
			data[20610] <= 8'h10 ;
			data[20611] <= 8'h10 ;
			data[20612] <= 8'h10 ;
			data[20613] <= 8'h10 ;
			data[20614] <= 8'h10 ;
			data[20615] <= 8'h10 ;
			data[20616] <= 8'h10 ;
			data[20617] <= 8'h10 ;
			data[20618] <= 8'h10 ;
			data[20619] <= 8'h10 ;
			data[20620] <= 8'h10 ;
			data[20621] <= 8'h10 ;
			data[20622] <= 8'h10 ;
			data[20623] <= 8'h10 ;
			data[20624] <= 8'h10 ;
			data[20625] <= 8'h10 ;
			data[20626] <= 8'h10 ;
			data[20627] <= 8'h10 ;
			data[20628] <= 8'h10 ;
			data[20629] <= 8'h10 ;
			data[20630] <= 8'h10 ;
			data[20631] <= 8'h10 ;
			data[20632] <= 8'h10 ;
			data[20633] <= 8'h10 ;
			data[20634] <= 8'h10 ;
			data[20635] <= 8'h10 ;
			data[20636] <= 8'h10 ;
			data[20637] <= 8'h10 ;
			data[20638] <= 8'h10 ;
			data[20639] <= 8'h10 ;
			data[20640] <= 8'h10 ;
			data[20641] <= 8'h10 ;
			data[20642] <= 8'h10 ;
			data[20643] <= 8'h10 ;
			data[20644] <= 8'h10 ;
			data[20645] <= 8'h10 ;
			data[20646] <= 8'h10 ;
			data[20647] <= 8'h10 ;
			data[20648] <= 8'h10 ;
			data[20649] <= 8'h10 ;
			data[20650] <= 8'h10 ;
			data[20651] <= 8'h10 ;
			data[20652] <= 8'h10 ;
			data[20653] <= 8'h10 ;
			data[20654] <= 8'h10 ;
			data[20655] <= 8'h10 ;
			data[20656] <= 8'h10 ;
			data[20657] <= 8'h10 ;
			data[20658] <= 8'h10 ;
			data[20659] <= 8'h10 ;
			data[20660] <= 8'h10 ;
			data[20661] <= 8'h10 ;
			data[20662] <= 8'h10 ;
			data[20663] <= 8'h10 ;
			data[20664] <= 8'h10 ;
			data[20665] <= 8'h10 ;
			data[20666] <= 8'h10 ;
			data[20667] <= 8'h10 ;
			data[20668] <= 8'h10 ;
			data[20669] <= 8'h10 ;
			data[20670] <= 8'h10 ;
			data[20671] <= 8'h10 ;
			data[20672] <= 8'h10 ;
			data[20673] <= 8'h10 ;
			data[20674] <= 8'h10 ;
			data[20675] <= 8'h10 ;
			data[20676] <= 8'h10 ;
			data[20677] <= 8'h10 ;
			data[20678] <= 8'h10 ;
			data[20679] <= 8'h10 ;
			data[20680] <= 8'h10 ;
			data[20681] <= 8'h10 ;
			data[20682] <= 8'h10 ;
			data[20683] <= 8'h10 ;
			data[20684] <= 8'h10 ;
			data[20685] <= 8'h10 ;
			data[20686] <= 8'h10 ;
			data[20687] <= 8'h10 ;
			data[20688] <= 8'h10 ;
			data[20689] <= 8'h10 ;
			data[20690] <= 8'h10 ;
			data[20691] <= 8'h10 ;
			data[20692] <= 8'h10 ;
			data[20693] <= 8'h10 ;
			data[20694] <= 8'h10 ;
			data[20695] <= 8'h10 ;
			data[20696] <= 8'h10 ;
			data[20697] <= 8'h10 ;
			data[20698] <= 8'h10 ;
			data[20699] <= 8'h10 ;
			data[20700] <= 8'h10 ;
			data[20701] <= 8'h10 ;
			data[20702] <= 8'h10 ;
			data[20703] <= 8'h10 ;
			data[20704] <= 8'h10 ;
			data[20705] <= 8'h10 ;
			data[20706] <= 8'h10 ;
			data[20707] <= 8'h10 ;
			data[20708] <= 8'h10 ;
			data[20709] <= 8'h10 ;
			data[20710] <= 8'h10 ;
			data[20711] <= 8'h10 ;
			data[20712] <= 8'h10 ;
			data[20713] <= 8'h10 ;
			data[20714] <= 8'h10 ;
			data[20715] <= 8'h10 ;
			data[20716] <= 8'h10 ;
			data[20717] <= 8'h10 ;
			data[20718] <= 8'h10 ;
			data[20719] <= 8'h10 ;
			data[20720] <= 8'h10 ;
			data[20721] <= 8'h10 ;
			data[20722] <= 8'h10 ;
			data[20723] <= 8'h10 ;
			data[20724] <= 8'h10 ;
			data[20725] <= 8'h10 ;
			data[20726] <= 8'h10 ;
			data[20727] <= 8'h10 ;
			data[20728] <= 8'h10 ;
			data[20729] <= 8'h10 ;
			data[20730] <= 8'h10 ;
			data[20731] <= 8'h10 ;
			data[20732] <= 8'h10 ;
			data[20733] <= 8'h10 ;
			data[20734] <= 8'h10 ;
			data[20735] <= 8'h10 ;
			data[20736] <= 8'h10 ;
			data[20737] <= 8'h10 ;
			data[20738] <= 8'h10 ;
			data[20739] <= 8'h10 ;
			data[20740] <= 8'h10 ;
			data[20741] <= 8'h10 ;
			data[20742] <= 8'h10 ;
			data[20743] <= 8'h10 ;
			data[20744] <= 8'h10 ;
			data[20745] <= 8'h10 ;
			data[20746] <= 8'h10 ;
			data[20747] <= 8'h10 ;
			data[20748] <= 8'h10 ;
			data[20749] <= 8'h10 ;
			data[20750] <= 8'h10 ;
			data[20751] <= 8'h10 ;
			data[20752] <= 8'h10 ;
			data[20753] <= 8'h10 ;
			data[20754] <= 8'h10 ;
			data[20755] <= 8'h10 ;
			data[20756] <= 8'h10 ;
			data[20757] <= 8'h10 ;
			data[20758] <= 8'h10 ;
			data[20759] <= 8'h10 ;
			data[20760] <= 8'h10 ;
			data[20761] <= 8'h10 ;
			data[20762] <= 8'h10 ;
			data[20763] <= 8'h10 ;
			data[20764] <= 8'h10 ;
			data[20765] <= 8'h10 ;
			data[20766] <= 8'h10 ;
			data[20767] <= 8'h10 ;
			data[20768] <= 8'h10 ;
			data[20769] <= 8'h10 ;
			data[20770] <= 8'h10 ;
			data[20771] <= 8'h10 ;
			data[20772] <= 8'h10 ;
			data[20773] <= 8'h10 ;
			data[20774] <= 8'h10 ;
			data[20775] <= 8'h10 ;
			data[20776] <= 8'h10 ;
			data[20777] <= 8'h10 ;
			data[20778] <= 8'h10 ;
			data[20779] <= 8'h10 ;
			data[20780] <= 8'h10 ;
			data[20781] <= 8'h10 ;
			data[20782] <= 8'h10 ;
			data[20783] <= 8'h10 ;
			data[20784] <= 8'h10 ;
			data[20785] <= 8'h10 ;
			data[20786] <= 8'h10 ;
			data[20787] <= 8'h10 ;
			data[20788] <= 8'h10 ;
			data[20789] <= 8'h10 ;
			data[20790] <= 8'h10 ;
			data[20791] <= 8'h10 ;
			data[20792] <= 8'h10 ;
			data[20793] <= 8'h10 ;
			data[20794] <= 8'h10 ;
			data[20795] <= 8'h10 ;
			data[20796] <= 8'h10 ;
			data[20797] <= 8'h10 ;
			data[20798] <= 8'h10 ;
			data[20799] <= 8'h10 ;
			data[20800] <= 8'h10 ;
			data[20801] <= 8'h10 ;
			data[20802] <= 8'h10 ;
			data[20803] <= 8'h10 ;
			data[20804] <= 8'h10 ;
			data[20805] <= 8'h10 ;
			data[20806] <= 8'h10 ;
			data[20807] <= 8'h10 ;
			data[20808] <= 8'h10 ;
			data[20809] <= 8'h10 ;
			data[20810] <= 8'h10 ;
			data[20811] <= 8'h10 ;
			data[20812] <= 8'h10 ;
			data[20813] <= 8'h10 ;
			data[20814] <= 8'h10 ;
			data[20815] <= 8'h10 ;
			data[20816] <= 8'h10 ;
			data[20817] <= 8'h10 ;
			data[20818] <= 8'h10 ;
			data[20819] <= 8'h10 ;
			data[20820] <= 8'h10 ;
			data[20821] <= 8'h10 ;
			data[20822] <= 8'h10 ;
			data[20823] <= 8'h10 ;
			data[20824] <= 8'h10 ;
			data[20825] <= 8'h10 ;
			data[20826] <= 8'h10 ;
			data[20827] <= 8'h10 ;
			data[20828] <= 8'h10 ;
			data[20829] <= 8'h10 ;
			data[20830] <= 8'h10 ;
			data[20831] <= 8'h10 ;
			data[20832] <= 8'h10 ;
			data[20833] <= 8'h10 ;
			data[20834] <= 8'h10 ;
			data[20835] <= 8'h10 ;
			data[20836] <= 8'h10 ;
			data[20837] <= 8'h10 ;
			data[20838] <= 8'h10 ;
			data[20839] <= 8'h10 ;
			data[20840] <= 8'h10 ;
			data[20841] <= 8'h10 ;
			data[20842] <= 8'h10 ;
			data[20843] <= 8'h10 ;
			data[20844] <= 8'h10 ;
			data[20845] <= 8'h10 ;
			data[20846] <= 8'h10 ;
			data[20847] <= 8'h10 ;
			data[20848] <= 8'h10 ;
			data[20849] <= 8'h10 ;
			data[20850] <= 8'h10 ;
			data[20851] <= 8'h10 ;
			data[20852] <= 8'h10 ;
			data[20853] <= 8'h10 ;
			data[20854] <= 8'h10 ;
			data[20855] <= 8'h10 ;
			data[20856] <= 8'h10 ;
			data[20857] <= 8'h10 ;
			data[20858] <= 8'h10 ;
			data[20859] <= 8'h10 ;
			data[20860] <= 8'h10 ;
			data[20861] <= 8'h10 ;
			data[20862] <= 8'h10 ;
			data[20863] <= 8'h10 ;
			data[20864] <= 8'h10 ;
			data[20865] <= 8'h10 ;
			data[20866] <= 8'h10 ;
			data[20867] <= 8'h10 ;
			data[20868] <= 8'h10 ;
			data[20869] <= 8'h10 ;
			data[20870] <= 8'h10 ;
			data[20871] <= 8'h10 ;
			data[20872] <= 8'h10 ;
			data[20873] <= 8'h10 ;
			data[20874] <= 8'h10 ;
			data[20875] <= 8'h10 ;
			data[20876] <= 8'h10 ;
			data[20877] <= 8'h10 ;
			data[20878] <= 8'h10 ;
			data[20879] <= 8'h10 ;
			data[20880] <= 8'h10 ;
			data[20881] <= 8'h10 ;
			data[20882] <= 8'h10 ;
			data[20883] <= 8'h10 ;
			data[20884] <= 8'h10 ;
			data[20885] <= 8'h10 ;
			data[20886] <= 8'h10 ;
			data[20887] <= 8'h10 ;
			data[20888] <= 8'h10 ;
			data[20889] <= 8'h10 ;
			data[20890] <= 8'h10 ;
			data[20891] <= 8'h10 ;
			data[20892] <= 8'h10 ;
			data[20893] <= 8'h10 ;
			data[20894] <= 8'h10 ;
			data[20895] <= 8'h10 ;
			data[20896] <= 8'h10 ;
			data[20897] <= 8'h10 ;
			data[20898] <= 8'h10 ;
			data[20899] <= 8'h10 ;
			data[20900] <= 8'h10 ;
			data[20901] <= 8'h10 ;
			data[20902] <= 8'h10 ;
			data[20903] <= 8'h10 ;
			data[20904] <= 8'h10 ;
			data[20905] <= 8'h10 ;
			data[20906] <= 8'h10 ;
			data[20907] <= 8'h10 ;
			data[20908] <= 8'h10 ;
			data[20909] <= 8'h10 ;
			data[20910] <= 8'h10 ;
			data[20911] <= 8'h10 ;
			data[20912] <= 8'h10 ;
			data[20913] <= 8'h10 ;
			data[20914] <= 8'h10 ;
			data[20915] <= 8'h10 ;
			data[20916] <= 8'h10 ;
			data[20917] <= 8'h10 ;
			data[20918] <= 8'h10 ;
			data[20919] <= 8'h10 ;
			data[20920] <= 8'h10 ;
			data[20921] <= 8'h10 ;
			data[20922] <= 8'h10 ;
			data[20923] <= 8'h10 ;
			data[20924] <= 8'h10 ;
			data[20925] <= 8'h10 ;
			data[20926] <= 8'h10 ;
			data[20927] <= 8'h10 ;
			data[20928] <= 8'h10 ;
			data[20929] <= 8'h10 ;
			data[20930] <= 8'h10 ;
			data[20931] <= 8'h10 ;
			data[20932] <= 8'h10 ;
			data[20933] <= 8'h10 ;
			data[20934] <= 8'h10 ;
			data[20935] <= 8'h10 ;
			data[20936] <= 8'h10 ;
			data[20937] <= 8'h10 ;
			data[20938] <= 8'h10 ;
			data[20939] <= 8'h10 ;
			data[20940] <= 8'h10 ;
			data[20941] <= 8'h10 ;
			data[20942] <= 8'h10 ;
			data[20943] <= 8'h10 ;
			data[20944] <= 8'h10 ;
			data[20945] <= 8'h10 ;
			data[20946] <= 8'h10 ;
			data[20947] <= 8'h10 ;
			data[20948] <= 8'h10 ;
			data[20949] <= 8'h10 ;
			data[20950] <= 8'h10 ;
			data[20951] <= 8'h10 ;
			data[20952] <= 8'h10 ;
			data[20953] <= 8'h10 ;
			data[20954] <= 8'h10 ;
			data[20955] <= 8'h10 ;
			data[20956] <= 8'h10 ;
			data[20957] <= 8'h10 ;
			data[20958] <= 8'h10 ;
			data[20959] <= 8'h10 ;
			data[20960] <= 8'h10 ;
			data[20961] <= 8'h10 ;
			data[20962] <= 8'h10 ;
			data[20963] <= 8'h10 ;
			data[20964] <= 8'h10 ;
			data[20965] <= 8'h10 ;
			data[20966] <= 8'h10 ;
			data[20967] <= 8'h10 ;
			data[20968] <= 8'h10 ;
			data[20969] <= 8'h10 ;
			data[20970] <= 8'h10 ;
			data[20971] <= 8'h10 ;
			data[20972] <= 8'h10 ;
			data[20973] <= 8'h10 ;
			data[20974] <= 8'h10 ;
			data[20975] <= 8'h10 ;
			data[20976] <= 8'h10 ;
			data[20977] <= 8'h10 ;
			data[20978] <= 8'h10 ;
			data[20979] <= 8'h10 ;
			data[20980] <= 8'h10 ;
			data[20981] <= 8'h10 ;
			data[20982] <= 8'h10 ;
			data[20983] <= 8'h10 ;
			data[20984] <= 8'h10 ;
			data[20985] <= 8'h10 ;
			data[20986] <= 8'h10 ;
			data[20987] <= 8'h10 ;
			data[20988] <= 8'h10 ;
			data[20989] <= 8'h10 ;
			data[20990] <= 8'h10 ;
			data[20991] <= 8'h10 ;
			data[20992] <= 8'h10 ;
			data[20993] <= 8'h10 ;
			data[20994] <= 8'h10 ;
			data[20995] <= 8'h10 ;
			data[20996] <= 8'h10 ;
			data[20997] <= 8'h10 ;
			data[20998] <= 8'h10 ;
			data[20999] <= 8'h10 ;
			data[21000] <= 8'h10 ;
			data[21001] <= 8'h10 ;
			data[21002] <= 8'h10 ;
			data[21003] <= 8'h10 ;
			data[21004] <= 8'h10 ;
			data[21005] <= 8'h10 ;
			data[21006] <= 8'h10 ;
			data[21007] <= 8'h10 ;
			data[21008] <= 8'h10 ;
			data[21009] <= 8'h10 ;
			data[21010] <= 8'h10 ;
			data[21011] <= 8'h10 ;
			data[21012] <= 8'h10 ;
			data[21013] <= 8'h10 ;
			data[21014] <= 8'h10 ;
			data[21015] <= 8'h10 ;
			data[21016] <= 8'h10 ;
			data[21017] <= 8'h10 ;
			data[21018] <= 8'h10 ;
			data[21019] <= 8'h10 ;
			data[21020] <= 8'h10 ;
			data[21021] <= 8'h10 ;
			data[21022] <= 8'h10 ;
			data[21023] <= 8'h10 ;
			data[21024] <= 8'h10 ;
			data[21025] <= 8'h10 ;
			data[21026] <= 8'h10 ;
			data[21027] <= 8'h10 ;
			data[21028] <= 8'h10 ;
			data[21029] <= 8'h10 ;
			data[21030] <= 8'h10 ;
			data[21031] <= 8'h10 ;
			data[21032] <= 8'h10 ;
			data[21033] <= 8'h10 ;
			data[21034] <= 8'h10 ;
			data[21035] <= 8'h10 ;
			data[21036] <= 8'h10 ;
			data[21037] <= 8'h10 ;
			data[21038] <= 8'h10 ;
			data[21039] <= 8'h10 ;
			data[21040] <= 8'h10 ;
			data[21041] <= 8'h10 ;
			data[21042] <= 8'h10 ;
			data[21043] <= 8'h10 ;
			data[21044] <= 8'h10 ;
			data[21045] <= 8'h10 ;
			data[21046] <= 8'h10 ;
			data[21047] <= 8'h10 ;
			data[21048] <= 8'h10 ;
			data[21049] <= 8'h10 ;
			data[21050] <= 8'h10 ;
			data[21051] <= 8'h10 ;
			data[21052] <= 8'h10 ;
			data[21053] <= 8'h10 ;
			data[21054] <= 8'h10 ;
			data[21055] <= 8'h10 ;
			data[21056] <= 8'h10 ;
			data[21057] <= 8'h10 ;
			data[21058] <= 8'h10 ;
			data[21059] <= 8'h10 ;
			data[21060] <= 8'h10 ;
			data[21061] <= 8'h10 ;
			data[21062] <= 8'h10 ;
			data[21063] <= 8'h10 ;
			data[21064] <= 8'h10 ;
			data[21065] <= 8'h10 ;
			data[21066] <= 8'h10 ;
			data[21067] <= 8'h10 ;
			data[21068] <= 8'h10 ;
			data[21069] <= 8'h10 ;
			data[21070] <= 8'h10 ;
			data[21071] <= 8'h10 ;
			data[21072] <= 8'h10 ;
			data[21073] <= 8'h10 ;
			data[21074] <= 8'h10 ;
			data[21075] <= 8'h10 ;
			data[21076] <= 8'h10 ;
			data[21077] <= 8'h10 ;
			data[21078] <= 8'h10 ;
			data[21079] <= 8'h10 ;
			data[21080] <= 8'h10 ;
			data[21081] <= 8'h10 ;
			data[21082] <= 8'h10 ;
			data[21083] <= 8'h10 ;
			data[21084] <= 8'h10 ;
			data[21085] <= 8'h10 ;
			data[21086] <= 8'h10 ;
			data[21087] <= 8'h10 ;
			data[21088] <= 8'h10 ;
			data[21089] <= 8'h10 ;
			data[21090] <= 8'h10 ;
			data[21091] <= 8'h10 ;
			data[21092] <= 8'h10 ;
			data[21093] <= 8'h10 ;
			data[21094] <= 8'h10 ;
			data[21095] <= 8'h10 ;
			data[21096] <= 8'h10 ;
			data[21097] <= 8'h10 ;
			data[21098] <= 8'h10 ;
			data[21099] <= 8'h10 ;
			data[21100] <= 8'h10 ;
			data[21101] <= 8'h10 ;
			data[21102] <= 8'h10 ;
			data[21103] <= 8'h10 ;
			data[21104] <= 8'h10 ;
			data[21105] <= 8'h10 ;
			data[21106] <= 8'h10 ;
			data[21107] <= 8'h10 ;
			data[21108] <= 8'h10 ;
			data[21109] <= 8'h10 ;
			data[21110] <= 8'h10 ;
			data[21111] <= 8'h10 ;
			data[21112] <= 8'h10 ;
			data[21113] <= 8'h10 ;
			data[21114] <= 8'h10 ;
			data[21115] <= 8'h10 ;
			data[21116] <= 8'h10 ;
			data[21117] <= 8'h10 ;
			data[21118] <= 8'h10 ;
			data[21119] <= 8'h10 ;
			data[21120] <= 8'h10 ;
			data[21121] <= 8'h10 ;
			data[21122] <= 8'h10 ;
			data[21123] <= 8'h10 ;
			data[21124] <= 8'h10 ;
			data[21125] <= 8'h10 ;
			data[21126] <= 8'h10 ;
			data[21127] <= 8'h10 ;
			data[21128] <= 8'h10 ;
			data[21129] <= 8'h10 ;
			data[21130] <= 8'h10 ;
			data[21131] <= 8'h10 ;
			data[21132] <= 8'h10 ;
			data[21133] <= 8'h10 ;
			data[21134] <= 8'h10 ;
			data[21135] <= 8'h10 ;
			data[21136] <= 8'h10 ;
			data[21137] <= 8'h10 ;
			data[21138] <= 8'h10 ;
			data[21139] <= 8'h10 ;
			data[21140] <= 8'h10 ;
			data[21141] <= 8'h10 ;
			data[21142] <= 8'h10 ;
			data[21143] <= 8'h10 ;
			data[21144] <= 8'h10 ;
			data[21145] <= 8'h10 ;
			data[21146] <= 8'h10 ;
			data[21147] <= 8'h10 ;
			data[21148] <= 8'h10 ;
			data[21149] <= 8'h10 ;
			data[21150] <= 8'h10 ;
			data[21151] <= 8'h10 ;
			data[21152] <= 8'h10 ;
			data[21153] <= 8'h10 ;
			data[21154] <= 8'h10 ;
			data[21155] <= 8'h10 ;
			data[21156] <= 8'h10 ;
			data[21157] <= 8'h10 ;
			data[21158] <= 8'h10 ;
			data[21159] <= 8'h10 ;
			data[21160] <= 8'h10 ;
			data[21161] <= 8'h10 ;
			data[21162] <= 8'h10 ;
			data[21163] <= 8'h10 ;
			data[21164] <= 8'h10 ;
			data[21165] <= 8'h10 ;
			data[21166] <= 8'h10 ;
			data[21167] <= 8'h10 ;
			data[21168] <= 8'h10 ;
			data[21169] <= 8'h10 ;
			data[21170] <= 8'h10 ;
			data[21171] <= 8'h10 ;
			data[21172] <= 8'h10 ;
			data[21173] <= 8'h10 ;
			data[21174] <= 8'h10 ;
			data[21175] <= 8'h10 ;
			data[21176] <= 8'h10 ;
			data[21177] <= 8'h10 ;
			data[21178] <= 8'h10 ;
			data[21179] <= 8'h10 ;
			data[21180] <= 8'h10 ;
			data[21181] <= 8'h10 ;
			data[21182] <= 8'h10 ;
			data[21183] <= 8'h10 ;
			data[21184] <= 8'h10 ;
			data[21185] <= 8'h10 ;
			data[21186] <= 8'h10 ;
			data[21187] <= 8'h10 ;
			data[21188] <= 8'h10 ;
			data[21189] <= 8'h10 ;
			data[21190] <= 8'h10 ;
			data[21191] <= 8'h10 ;
			data[21192] <= 8'h10 ;
			data[21193] <= 8'h10 ;
			data[21194] <= 8'h10 ;
			data[21195] <= 8'h10 ;
			data[21196] <= 8'h10 ;
			data[21197] <= 8'h10 ;
			data[21198] <= 8'h10 ;
			data[21199] <= 8'h10 ;
			data[21200] <= 8'h10 ;
			data[21201] <= 8'h10 ;
			data[21202] <= 8'h10 ;
			data[21203] <= 8'h10 ;
			data[21204] <= 8'h10 ;
			data[21205] <= 8'h10 ;
			data[21206] <= 8'h10 ;
			data[21207] <= 8'h10 ;
			data[21208] <= 8'h10 ;
			data[21209] <= 8'h10 ;
			data[21210] <= 8'h10 ;
			data[21211] <= 8'h10 ;
			data[21212] <= 8'h10 ;
			data[21213] <= 8'h10 ;
			data[21214] <= 8'h10 ;
			data[21215] <= 8'h10 ;
			data[21216] <= 8'h10 ;
			data[21217] <= 8'h10 ;
			data[21218] <= 8'h10 ;
			data[21219] <= 8'h10 ;
			data[21220] <= 8'h10 ;
			data[21221] <= 8'h10 ;
			data[21222] <= 8'h10 ;
			data[21223] <= 8'h10 ;
			data[21224] <= 8'h10 ;
			data[21225] <= 8'h10 ;
			data[21226] <= 8'h10 ;
			data[21227] <= 8'h10 ;
			data[21228] <= 8'h10 ;
			data[21229] <= 8'h10 ;
			data[21230] <= 8'h10 ;
			data[21231] <= 8'h10 ;
			data[21232] <= 8'h10 ;
			data[21233] <= 8'h10 ;
			data[21234] <= 8'h10 ;
			data[21235] <= 8'h10 ;
			data[21236] <= 8'h10 ;
			data[21237] <= 8'h10 ;
			data[21238] <= 8'h10 ;
			data[21239] <= 8'h10 ;
			data[21240] <= 8'h10 ;
			data[21241] <= 8'h10 ;
			data[21242] <= 8'h10 ;
			data[21243] <= 8'h10 ;
			data[21244] <= 8'h10 ;
			data[21245] <= 8'h10 ;
			data[21246] <= 8'h10 ;
			data[21247] <= 8'h10 ;
			data[21248] <= 8'h10 ;
			data[21249] <= 8'h10 ;
			data[21250] <= 8'h10 ;
			data[21251] <= 8'h10 ;
			data[21252] <= 8'h10 ;
			data[21253] <= 8'h10 ;
			data[21254] <= 8'h10 ;
			data[21255] <= 8'h10 ;
			data[21256] <= 8'h10 ;
			data[21257] <= 8'h10 ;
			data[21258] <= 8'h10 ;
			data[21259] <= 8'h10 ;
			data[21260] <= 8'h10 ;
			data[21261] <= 8'h10 ;
			data[21262] <= 8'h10 ;
			data[21263] <= 8'h10 ;
			data[21264] <= 8'h10 ;
			data[21265] <= 8'h10 ;
			data[21266] <= 8'h10 ;
			data[21267] <= 8'h10 ;
			data[21268] <= 8'h10 ;
			data[21269] <= 8'h10 ;
			data[21270] <= 8'h10 ;
			data[21271] <= 8'h10 ;
			data[21272] <= 8'h10 ;
			data[21273] <= 8'h10 ;
			data[21274] <= 8'h10 ;
			data[21275] <= 8'h10 ;
			data[21276] <= 8'h10 ;
			data[21277] <= 8'h10 ;
			data[21278] <= 8'h10 ;
			data[21279] <= 8'h10 ;
			data[21280] <= 8'h10 ;
			data[21281] <= 8'h10 ;
			data[21282] <= 8'h10 ;
			data[21283] <= 8'h10 ;
			data[21284] <= 8'h10 ;
			data[21285] <= 8'h10 ;
			data[21286] <= 8'h10 ;
			data[21287] <= 8'h10 ;
			data[21288] <= 8'h10 ;
			data[21289] <= 8'h10 ;
			data[21290] <= 8'h10 ;
			data[21291] <= 8'h10 ;
			data[21292] <= 8'h10 ;
			data[21293] <= 8'h10 ;
			data[21294] <= 8'h10 ;
			data[21295] <= 8'h10 ;
			data[21296] <= 8'h10 ;
			data[21297] <= 8'h10 ;
			data[21298] <= 8'h10 ;
			data[21299] <= 8'h10 ;
			data[21300] <= 8'h10 ;
			data[21301] <= 8'h10 ;
			data[21302] <= 8'h10 ;
			data[21303] <= 8'h10 ;
			data[21304] <= 8'h10 ;
			data[21305] <= 8'h10 ;
			data[21306] <= 8'h10 ;
			data[21307] <= 8'h10 ;
			data[21308] <= 8'h10 ;
			data[21309] <= 8'h10 ;
			data[21310] <= 8'h10 ;
			data[21311] <= 8'h10 ;
			data[21312] <= 8'h10 ;
			data[21313] <= 8'h10 ;
			data[21314] <= 8'h10 ;
			data[21315] <= 8'h10 ;
			data[21316] <= 8'h10 ;
			data[21317] <= 8'h10 ;
			data[21318] <= 8'h10 ;
			data[21319] <= 8'h10 ;
			data[21320] <= 8'h10 ;
			data[21321] <= 8'h10 ;
			data[21322] <= 8'h10 ;
			data[21323] <= 8'h10 ;
			data[21324] <= 8'h10 ;
			data[21325] <= 8'h10 ;
			data[21326] <= 8'h10 ;
			data[21327] <= 8'h10 ;
			data[21328] <= 8'h10 ;
			data[21329] <= 8'h10 ;
			data[21330] <= 8'h10 ;
			data[21331] <= 8'h10 ;
			data[21332] <= 8'h10 ;
			data[21333] <= 8'h10 ;
			data[21334] <= 8'h10 ;
			data[21335] <= 8'h10 ;
			data[21336] <= 8'h10 ;
			data[21337] <= 8'h10 ;
			data[21338] <= 8'h10 ;
			data[21339] <= 8'h10 ;
			data[21340] <= 8'h10 ;
			data[21341] <= 8'h10 ;
			data[21342] <= 8'h10 ;
			data[21343] <= 8'h10 ;
			data[21344] <= 8'h10 ;
			data[21345] <= 8'h10 ;
			data[21346] <= 8'h10 ;
			data[21347] <= 8'h10 ;
			data[21348] <= 8'h10 ;
			data[21349] <= 8'h10 ;
			data[21350] <= 8'h10 ;
			data[21351] <= 8'h10 ;
			data[21352] <= 8'h10 ;
			data[21353] <= 8'h10 ;
			data[21354] <= 8'h10 ;
			data[21355] <= 8'h10 ;
			data[21356] <= 8'h10 ;
			data[21357] <= 8'h10 ;
			data[21358] <= 8'h10 ;
			data[21359] <= 8'h10 ;
			data[21360] <= 8'h10 ;
			data[21361] <= 8'h10 ;
			data[21362] <= 8'h10 ;
			data[21363] <= 8'h10 ;
			data[21364] <= 8'h10 ;
			data[21365] <= 8'h10 ;
			data[21366] <= 8'h10 ;
			data[21367] <= 8'h10 ;
			data[21368] <= 8'h10 ;
			data[21369] <= 8'h10 ;
			data[21370] <= 8'h10 ;
			data[21371] <= 8'h10 ;
			data[21372] <= 8'h10 ;
			data[21373] <= 8'h10 ;
			data[21374] <= 8'h10 ;
			data[21375] <= 8'h10 ;
			data[21376] <= 8'h10 ;
			data[21377] <= 8'h10 ;
			data[21378] <= 8'h10 ;
			data[21379] <= 8'h10 ;
			data[21380] <= 8'h10 ;
			data[21381] <= 8'h10 ;
			data[21382] <= 8'h10 ;
			data[21383] <= 8'h10 ;
			data[21384] <= 8'h10 ;
			data[21385] <= 8'h10 ;
			data[21386] <= 8'h10 ;
			data[21387] <= 8'h10 ;
			data[21388] <= 8'h10 ;
			data[21389] <= 8'h10 ;
			data[21390] <= 8'h10 ;
			data[21391] <= 8'h10 ;
			data[21392] <= 8'h10 ;
			data[21393] <= 8'h10 ;
			data[21394] <= 8'h10 ;
			data[21395] <= 8'h10 ;
			data[21396] <= 8'h10 ;
			data[21397] <= 8'h10 ;
			data[21398] <= 8'h10 ;
			data[21399] <= 8'h10 ;
			data[21400] <= 8'h10 ;
			data[21401] <= 8'h10 ;
			data[21402] <= 8'h10 ;
			data[21403] <= 8'h10 ;
			data[21404] <= 8'h10 ;
			data[21405] <= 8'h10 ;
			data[21406] <= 8'h10 ;
			data[21407] <= 8'h10 ;
			data[21408] <= 8'h10 ;
			data[21409] <= 8'h10 ;
			data[21410] <= 8'h10 ;
			data[21411] <= 8'h10 ;
			data[21412] <= 8'h10 ;
			data[21413] <= 8'h10 ;
			data[21414] <= 8'h10 ;
			data[21415] <= 8'h10 ;
			data[21416] <= 8'h10 ;
			data[21417] <= 8'h10 ;
			data[21418] <= 8'h10 ;
			data[21419] <= 8'h10 ;
			data[21420] <= 8'h10 ;
			data[21421] <= 8'h10 ;
			data[21422] <= 8'h10 ;
			data[21423] <= 8'h10 ;
			data[21424] <= 8'h10 ;
			data[21425] <= 8'h10 ;
			data[21426] <= 8'h10 ;
			data[21427] <= 8'h10 ;
			data[21428] <= 8'h10 ;
			data[21429] <= 8'h10 ;
			data[21430] <= 8'h10 ;
			data[21431] <= 8'h10 ;
			data[21432] <= 8'h10 ;
			data[21433] <= 8'h10 ;
			data[21434] <= 8'h10 ;
			data[21435] <= 8'h10 ;
			data[21436] <= 8'h10 ;
			data[21437] <= 8'h10 ;
			data[21438] <= 8'h10 ;
			data[21439] <= 8'h10 ;
			data[21440] <= 8'h10 ;
			data[21441] <= 8'h10 ;
			data[21442] <= 8'h10 ;
			data[21443] <= 8'h10 ;
			data[21444] <= 8'h10 ;
			data[21445] <= 8'h10 ;
			data[21446] <= 8'h10 ;
			data[21447] <= 8'h10 ;
			data[21448] <= 8'h10 ;
			data[21449] <= 8'h10 ;
			data[21450] <= 8'h10 ;
			data[21451] <= 8'h10 ;
			data[21452] <= 8'h10 ;
			data[21453] <= 8'h10 ;
			data[21454] <= 8'h10 ;
			data[21455] <= 8'h10 ;
			data[21456] <= 8'h10 ;
			data[21457] <= 8'h10 ;
			data[21458] <= 8'h10 ;
			data[21459] <= 8'h10 ;
			data[21460] <= 8'h10 ;
			data[21461] <= 8'h10 ;
			data[21462] <= 8'h10 ;
			data[21463] <= 8'h10 ;
			data[21464] <= 8'h10 ;
			data[21465] <= 8'h10 ;
			data[21466] <= 8'h10 ;
			data[21467] <= 8'h10 ;
			data[21468] <= 8'h10 ;
			data[21469] <= 8'h10 ;
			data[21470] <= 8'h10 ;
			data[21471] <= 8'h10 ;
			data[21472] <= 8'h10 ;
			data[21473] <= 8'h10 ;
			data[21474] <= 8'h10 ;
			data[21475] <= 8'h10 ;
			data[21476] <= 8'h10 ;
			data[21477] <= 8'h10 ;
			data[21478] <= 8'h10 ;
			data[21479] <= 8'h10 ;
			data[21480] <= 8'h10 ;
			data[21481] <= 8'h10 ;
			data[21482] <= 8'h10 ;
			data[21483] <= 8'h10 ;
			data[21484] <= 8'h10 ;
			data[21485] <= 8'h10 ;
			data[21486] <= 8'h10 ;
			data[21487] <= 8'h10 ;
			data[21488] <= 8'h10 ;
			data[21489] <= 8'h10 ;
			data[21490] <= 8'h10 ;
			data[21491] <= 8'h10 ;
			data[21492] <= 8'h10 ;
			data[21493] <= 8'h10 ;
			data[21494] <= 8'h10 ;
			data[21495] <= 8'h10 ;
			data[21496] <= 8'h10 ;
			data[21497] <= 8'h10 ;
			data[21498] <= 8'h10 ;
			data[21499] <= 8'h10 ;
			data[21500] <= 8'h10 ;
			data[21501] <= 8'h10 ;
			data[21502] <= 8'h10 ;
			data[21503] <= 8'h10 ;
			data[21504] <= 8'h10 ;
			data[21505] <= 8'h10 ;
			data[21506] <= 8'h10 ;
			data[21507] <= 8'h10 ;
			data[21508] <= 8'h10 ;
			data[21509] <= 8'h10 ;
			data[21510] <= 8'h10 ;
			data[21511] <= 8'h10 ;
			data[21512] <= 8'h10 ;
			data[21513] <= 8'h10 ;
			data[21514] <= 8'h10 ;
			data[21515] <= 8'h10 ;
			data[21516] <= 8'h10 ;
			data[21517] <= 8'h10 ;
			data[21518] <= 8'h10 ;
			data[21519] <= 8'h10 ;
			data[21520] <= 8'h10 ;
			data[21521] <= 8'h10 ;
			data[21522] <= 8'h10 ;
			data[21523] <= 8'h10 ;
			data[21524] <= 8'h10 ;
			data[21525] <= 8'h10 ;
			data[21526] <= 8'h10 ;
			data[21527] <= 8'h10 ;
			data[21528] <= 8'h10 ;
			data[21529] <= 8'h10 ;
			data[21530] <= 8'h10 ;
			data[21531] <= 8'h10 ;
			data[21532] <= 8'h10 ;
			data[21533] <= 8'h10 ;
			data[21534] <= 8'h10 ;
			data[21535] <= 8'h10 ;
			data[21536] <= 8'h10 ;
			data[21537] <= 8'h10 ;
			data[21538] <= 8'h10 ;
			data[21539] <= 8'h10 ;
			data[21540] <= 8'h10 ;
			data[21541] <= 8'h10 ;
			data[21542] <= 8'h10 ;
			data[21543] <= 8'h10 ;
			data[21544] <= 8'h10 ;
			data[21545] <= 8'h10 ;
			data[21546] <= 8'h10 ;
			data[21547] <= 8'h10 ;
			data[21548] <= 8'h10 ;
			data[21549] <= 8'h10 ;
			data[21550] <= 8'h10 ;
			data[21551] <= 8'h10 ;
			data[21552] <= 8'h10 ;
			data[21553] <= 8'h10 ;
			data[21554] <= 8'h10 ;
			data[21555] <= 8'h10 ;
			data[21556] <= 8'h10 ;
			data[21557] <= 8'h10 ;
			data[21558] <= 8'h10 ;
			data[21559] <= 8'h10 ;
			data[21560] <= 8'h10 ;
			data[21561] <= 8'h10 ;
			data[21562] <= 8'h10 ;
			data[21563] <= 8'h10 ;
			data[21564] <= 8'h10 ;
			data[21565] <= 8'h10 ;
			data[21566] <= 8'h10 ;
			data[21567] <= 8'h10 ;
			data[21568] <= 8'h10 ;
			data[21569] <= 8'h10 ;
			data[21570] <= 8'h10 ;
			data[21571] <= 8'h10 ;
			data[21572] <= 8'h10 ;
			data[21573] <= 8'h10 ;
			data[21574] <= 8'h10 ;
			data[21575] <= 8'h10 ;
			data[21576] <= 8'h10 ;
			data[21577] <= 8'h10 ;
			data[21578] <= 8'h10 ;
			data[21579] <= 8'h10 ;
			data[21580] <= 8'h10 ;
			data[21581] <= 8'h10 ;
			data[21582] <= 8'h10 ;
			data[21583] <= 8'h10 ;
			data[21584] <= 8'h10 ;
			data[21585] <= 8'h10 ;
			data[21586] <= 8'h10 ;
			data[21587] <= 8'h10 ;
			data[21588] <= 8'h10 ;
			data[21589] <= 8'h10 ;
			data[21590] <= 8'h10 ;
			data[21591] <= 8'h10 ;
			data[21592] <= 8'h10 ;
			data[21593] <= 8'h10 ;
			data[21594] <= 8'h10 ;
			data[21595] <= 8'h10 ;
			data[21596] <= 8'h10 ;
			data[21597] <= 8'h10 ;
			data[21598] <= 8'h10 ;
			data[21599] <= 8'h10 ;
			data[21600] <= 8'h10 ;
			data[21601] <= 8'h10 ;
			data[21602] <= 8'h10 ;
			data[21603] <= 8'h10 ;
			data[21604] <= 8'h10 ;
			data[21605] <= 8'h10 ;
			data[21606] <= 8'h10 ;
			data[21607] <= 8'h10 ;
			data[21608] <= 8'h10 ;
			data[21609] <= 8'h10 ;
			data[21610] <= 8'h10 ;
			data[21611] <= 8'h10 ;
			data[21612] <= 8'h10 ;
			data[21613] <= 8'h10 ;
			data[21614] <= 8'h10 ;
			data[21615] <= 8'h10 ;
			data[21616] <= 8'h10 ;
			data[21617] <= 8'h10 ;
			data[21618] <= 8'h10 ;
			data[21619] <= 8'h10 ;
			data[21620] <= 8'h10 ;
			data[21621] <= 8'h10 ;
			data[21622] <= 8'h10 ;
			data[21623] <= 8'h10 ;
			data[21624] <= 8'h10 ;
			data[21625] <= 8'h10 ;
			data[21626] <= 8'h10 ;
			data[21627] <= 8'h10 ;
			data[21628] <= 8'h10 ;
			data[21629] <= 8'h10 ;
			data[21630] <= 8'h10 ;
			data[21631] <= 8'h10 ;
			data[21632] <= 8'h10 ;
			data[21633] <= 8'h10 ;
			data[21634] <= 8'h10 ;
			data[21635] <= 8'h10 ;
			data[21636] <= 8'h10 ;
			data[21637] <= 8'h10 ;
			data[21638] <= 8'h10 ;
			data[21639] <= 8'h10 ;
			data[21640] <= 8'h10 ;
			data[21641] <= 8'h10 ;
			data[21642] <= 8'h10 ;
			data[21643] <= 8'h10 ;
			data[21644] <= 8'h10 ;
			data[21645] <= 8'h10 ;
			data[21646] <= 8'h10 ;
			data[21647] <= 8'h10 ;
			data[21648] <= 8'h10 ;
			data[21649] <= 8'h10 ;
			data[21650] <= 8'h10 ;
			data[21651] <= 8'h10 ;
			data[21652] <= 8'h10 ;
			data[21653] <= 8'h10 ;
			data[21654] <= 8'h10 ;
			data[21655] <= 8'h10 ;
			data[21656] <= 8'h10 ;
			data[21657] <= 8'h10 ;
			data[21658] <= 8'h10 ;
			data[21659] <= 8'h10 ;
			data[21660] <= 8'h10 ;
			data[21661] <= 8'h10 ;
			data[21662] <= 8'h10 ;
			data[21663] <= 8'h10 ;
			data[21664] <= 8'h10 ;
			data[21665] <= 8'h10 ;
			data[21666] <= 8'h10 ;
			data[21667] <= 8'h10 ;
			data[21668] <= 8'h10 ;
			data[21669] <= 8'h10 ;
			data[21670] <= 8'h10 ;
			data[21671] <= 8'h10 ;
			data[21672] <= 8'h10 ;
			data[21673] <= 8'h10 ;
			data[21674] <= 8'h10 ;
			data[21675] <= 8'h10 ;
			data[21676] <= 8'h10 ;
			data[21677] <= 8'h10 ;
			data[21678] <= 8'h10 ;
			data[21679] <= 8'h10 ;
			data[21680] <= 8'h10 ;
			data[21681] <= 8'h10 ;
			data[21682] <= 8'h10 ;
			data[21683] <= 8'h10 ;
			data[21684] <= 8'h10 ;
			data[21685] <= 8'h10 ;
			data[21686] <= 8'h10 ;
			data[21687] <= 8'h10 ;
			data[21688] <= 8'h10 ;
			data[21689] <= 8'h10 ;
			data[21690] <= 8'h10 ;
			data[21691] <= 8'h10 ;
			data[21692] <= 8'h10 ;
			data[21693] <= 8'h10 ;
			data[21694] <= 8'h10 ;
			data[21695] <= 8'h10 ;
			data[21696] <= 8'h10 ;
			data[21697] <= 8'h10 ;
			data[21698] <= 8'h10 ;
			data[21699] <= 8'h10 ;
			data[21700] <= 8'h10 ;
			data[21701] <= 8'h10 ;
			data[21702] <= 8'h10 ;
			data[21703] <= 8'h10 ;
			data[21704] <= 8'h10 ;
			data[21705] <= 8'h10 ;
			data[21706] <= 8'h10 ;
			data[21707] <= 8'h10 ;
			data[21708] <= 8'h10 ;
			data[21709] <= 8'h10 ;
			data[21710] <= 8'h10 ;
			data[21711] <= 8'h10 ;
			data[21712] <= 8'h10 ;
			data[21713] <= 8'h10 ;
			data[21714] <= 8'h10 ;
			data[21715] <= 8'h10 ;
			data[21716] <= 8'h10 ;
			data[21717] <= 8'h10 ;
			data[21718] <= 8'h10 ;
			data[21719] <= 8'h10 ;
			data[21720] <= 8'h10 ;
			data[21721] <= 8'h10 ;
			data[21722] <= 8'h10 ;
			data[21723] <= 8'h10 ;
			data[21724] <= 8'h10 ;
			data[21725] <= 8'h10 ;
			data[21726] <= 8'h10 ;
			data[21727] <= 8'h10 ;
			data[21728] <= 8'h10 ;
			data[21729] <= 8'h10 ;
			data[21730] <= 8'h10 ;
			data[21731] <= 8'h10 ;
			data[21732] <= 8'h10 ;
			data[21733] <= 8'h10 ;
			data[21734] <= 8'h10 ;
			data[21735] <= 8'h10 ;
			data[21736] <= 8'h10 ;
			data[21737] <= 8'h10 ;
			data[21738] <= 8'h10 ;
			data[21739] <= 8'h10 ;
			data[21740] <= 8'h10 ;
			data[21741] <= 8'h10 ;
			data[21742] <= 8'h10 ;
			data[21743] <= 8'h10 ;
			data[21744] <= 8'h10 ;
			data[21745] <= 8'h10 ;
			data[21746] <= 8'h10 ;
			data[21747] <= 8'h10 ;
			data[21748] <= 8'h10 ;
			data[21749] <= 8'h10 ;
			data[21750] <= 8'h10 ;
			data[21751] <= 8'h10 ;
			data[21752] <= 8'h10 ;
			data[21753] <= 8'h10 ;
			data[21754] <= 8'h10 ;
			data[21755] <= 8'h10 ;
			data[21756] <= 8'h10 ;
			data[21757] <= 8'h10 ;
			data[21758] <= 8'h10 ;
			data[21759] <= 8'h10 ;
			data[21760] <= 8'h10 ;
			data[21761] <= 8'h10 ;
			data[21762] <= 8'h10 ;
			data[21763] <= 8'h10 ;
			data[21764] <= 8'h10 ;
			data[21765] <= 8'h10 ;
			data[21766] <= 8'h10 ;
			data[21767] <= 8'h10 ;
			data[21768] <= 8'h10 ;
			data[21769] <= 8'h10 ;
			data[21770] <= 8'h10 ;
			data[21771] <= 8'h10 ;
			data[21772] <= 8'h10 ;
			data[21773] <= 8'h10 ;
			data[21774] <= 8'h10 ;
			data[21775] <= 8'h10 ;
			data[21776] <= 8'h10 ;
			data[21777] <= 8'h10 ;
			data[21778] <= 8'h10 ;
			data[21779] <= 8'h10 ;
			data[21780] <= 8'h10 ;
			data[21781] <= 8'h10 ;
			data[21782] <= 8'h10 ;
			data[21783] <= 8'h10 ;
			data[21784] <= 8'h10 ;
			data[21785] <= 8'h10 ;
			data[21786] <= 8'h10 ;
			data[21787] <= 8'h10 ;
			data[21788] <= 8'h10 ;
			data[21789] <= 8'h10 ;
			data[21790] <= 8'h10 ;
			data[21791] <= 8'h10 ;
			data[21792] <= 8'h10 ;
			data[21793] <= 8'h10 ;
			data[21794] <= 8'h10 ;
			data[21795] <= 8'h10 ;
			data[21796] <= 8'h10 ;
			data[21797] <= 8'h10 ;
			data[21798] <= 8'h10 ;
			data[21799] <= 8'h10 ;
			data[21800] <= 8'h10 ;
			data[21801] <= 8'h10 ;
			data[21802] <= 8'h10 ;
			data[21803] <= 8'h10 ;
			data[21804] <= 8'h10 ;
			data[21805] <= 8'h10 ;
			data[21806] <= 8'h10 ;
			data[21807] <= 8'h10 ;
			data[21808] <= 8'h10 ;
			data[21809] <= 8'h10 ;
			data[21810] <= 8'h10 ;
			data[21811] <= 8'h10 ;
			data[21812] <= 8'h10 ;
			data[21813] <= 8'h10 ;
			data[21814] <= 8'h10 ;
			data[21815] <= 8'h10 ;
			data[21816] <= 8'h10 ;
			data[21817] <= 8'h10 ;
			data[21818] <= 8'h10 ;
			data[21819] <= 8'h10 ;
			data[21820] <= 8'h10 ;
			data[21821] <= 8'h10 ;
			data[21822] <= 8'h10 ;
			data[21823] <= 8'h10 ;
			data[21824] <= 8'h10 ;
			data[21825] <= 8'h10 ;
			data[21826] <= 8'h10 ;
			data[21827] <= 8'h10 ;
			data[21828] <= 8'h10 ;
			data[21829] <= 8'h10 ;
			data[21830] <= 8'h10 ;
			data[21831] <= 8'h10 ;
			data[21832] <= 8'h10 ;
			data[21833] <= 8'h10 ;
			data[21834] <= 8'h10 ;
			data[21835] <= 8'h10 ;
			data[21836] <= 8'h10 ;
			data[21837] <= 8'h10 ;
			data[21838] <= 8'h10 ;
			data[21839] <= 8'h10 ;
			data[21840] <= 8'h10 ;
			data[21841] <= 8'h10 ;
			data[21842] <= 8'h10 ;
			data[21843] <= 8'h10 ;
			data[21844] <= 8'h10 ;
			data[21845] <= 8'h10 ;
			data[21846] <= 8'h10 ;
			data[21847] <= 8'h10 ;
			data[21848] <= 8'h10 ;
			data[21849] <= 8'h10 ;
			data[21850] <= 8'h10 ;
			data[21851] <= 8'h10 ;
			data[21852] <= 8'h10 ;
			data[21853] <= 8'h10 ;
			data[21854] <= 8'h10 ;
			data[21855] <= 8'h10 ;
			data[21856] <= 8'h10 ;
			data[21857] <= 8'h10 ;
			data[21858] <= 8'h10 ;
			data[21859] <= 8'h10 ;
			data[21860] <= 8'h10 ;
			data[21861] <= 8'h10 ;
			data[21862] <= 8'h10 ;
			data[21863] <= 8'h10 ;
			data[21864] <= 8'h10 ;
			data[21865] <= 8'h10 ;
			data[21866] <= 8'h10 ;
			data[21867] <= 8'h10 ;
			data[21868] <= 8'h10 ;
			data[21869] <= 8'h10 ;
			data[21870] <= 8'h10 ;
			data[21871] <= 8'h10 ;
			data[21872] <= 8'h10 ;
			data[21873] <= 8'h10 ;
			data[21874] <= 8'h10 ;
			data[21875] <= 8'h10 ;
			data[21876] <= 8'h10 ;
			data[21877] <= 8'h10 ;
			data[21878] <= 8'h10 ;
			data[21879] <= 8'h10 ;
			data[21880] <= 8'h10 ;
			data[21881] <= 8'h10 ;
			data[21882] <= 8'h10 ;
			data[21883] <= 8'h10 ;
			data[21884] <= 8'h10 ;
			data[21885] <= 8'h10 ;
			data[21886] <= 8'h10 ;
			data[21887] <= 8'h10 ;
			data[21888] <= 8'h10 ;
			data[21889] <= 8'h10 ;
			data[21890] <= 8'h10 ;
			data[21891] <= 8'h10 ;
			data[21892] <= 8'h10 ;
			data[21893] <= 8'h10 ;
			data[21894] <= 8'h10 ;
			data[21895] <= 8'h10 ;
			data[21896] <= 8'h10 ;
			data[21897] <= 8'h10 ;
			data[21898] <= 8'h10 ;
			data[21899] <= 8'h10 ;
			data[21900] <= 8'h10 ;
			data[21901] <= 8'h10 ;
			data[21902] <= 8'h10 ;
			data[21903] <= 8'h10 ;
			data[21904] <= 8'h10 ;
			data[21905] <= 8'h10 ;
			data[21906] <= 8'h10 ;
			data[21907] <= 8'h10 ;
			data[21908] <= 8'h10 ;
			data[21909] <= 8'h10 ;
			data[21910] <= 8'h10 ;
			data[21911] <= 8'h10 ;
			data[21912] <= 8'h10 ;
			data[21913] <= 8'h10 ;
			data[21914] <= 8'h10 ;
			data[21915] <= 8'h10 ;
			data[21916] <= 8'h10 ;
			data[21917] <= 8'h10 ;
			data[21918] <= 8'h10 ;
			data[21919] <= 8'h10 ;
			data[21920] <= 8'h10 ;
			data[21921] <= 8'h10 ;
			data[21922] <= 8'h10 ;
			data[21923] <= 8'h10 ;
			data[21924] <= 8'h10 ;
			data[21925] <= 8'h10 ;
			data[21926] <= 8'h10 ;
			data[21927] <= 8'h10 ;
			data[21928] <= 8'h10 ;
			data[21929] <= 8'h10 ;
			data[21930] <= 8'h10 ;
			data[21931] <= 8'h10 ;
			data[21932] <= 8'h10 ;
			data[21933] <= 8'h10 ;
			data[21934] <= 8'h10 ;
			data[21935] <= 8'h10 ;
			data[21936] <= 8'h10 ;
			data[21937] <= 8'h10 ;
			data[21938] <= 8'h10 ;
			data[21939] <= 8'h10 ;
			data[21940] <= 8'h10 ;
			data[21941] <= 8'h10 ;
			data[21942] <= 8'h10 ;
			data[21943] <= 8'h10 ;
			data[21944] <= 8'h10 ;
			data[21945] <= 8'h10 ;
			data[21946] <= 8'h10 ;
			data[21947] <= 8'h10 ;
			data[21948] <= 8'h10 ;
			data[21949] <= 8'h10 ;
			data[21950] <= 8'h10 ;
			data[21951] <= 8'h10 ;
			data[21952] <= 8'h10 ;
			data[21953] <= 8'h10 ;
			data[21954] <= 8'h10 ;
			data[21955] <= 8'h10 ;
			data[21956] <= 8'h10 ;
			data[21957] <= 8'h10 ;
			data[21958] <= 8'h10 ;
			data[21959] <= 8'h10 ;
			data[21960] <= 8'h10 ;
			data[21961] <= 8'h10 ;
			data[21962] <= 8'h10 ;
			data[21963] <= 8'h10 ;
			data[21964] <= 8'h10 ;
			data[21965] <= 8'h10 ;
			data[21966] <= 8'h10 ;
			data[21967] <= 8'h10 ;
			data[21968] <= 8'h10 ;
			data[21969] <= 8'h10 ;
			data[21970] <= 8'h10 ;
			data[21971] <= 8'h10 ;
			data[21972] <= 8'h10 ;
			data[21973] <= 8'h10 ;
			data[21974] <= 8'h10 ;
			data[21975] <= 8'h10 ;
			data[21976] <= 8'h10 ;
			data[21977] <= 8'h10 ;
			data[21978] <= 8'h10 ;
			data[21979] <= 8'h10 ;
			data[21980] <= 8'h10 ;
			data[21981] <= 8'h10 ;
			data[21982] <= 8'h10 ;
			data[21983] <= 8'h10 ;
			data[21984] <= 8'h10 ;
			data[21985] <= 8'h10 ;
			data[21986] <= 8'h10 ;
			data[21987] <= 8'h10 ;
			data[21988] <= 8'h10 ;
			data[21989] <= 8'h10 ;
			data[21990] <= 8'h10 ;
			data[21991] <= 8'h10 ;
			data[21992] <= 8'h10 ;
			data[21993] <= 8'h10 ;
			data[21994] <= 8'h10 ;
			data[21995] <= 8'h10 ;
			data[21996] <= 8'h10 ;
			data[21997] <= 8'h10 ;
			data[21998] <= 8'h10 ;
			data[21999] <= 8'h10 ;
			data[22000] <= 8'h10 ;
			data[22001] <= 8'h10 ;
			data[22002] <= 8'h10 ;
			data[22003] <= 8'h10 ;
			data[22004] <= 8'h10 ;
			data[22005] <= 8'h10 ;
			data[22006] <= 8'h10 ;
			data[22007] <= 8'h10 ;
			data[22008] <= 8'h10 ;
			data[22009] <= 8'h10 ;
			data[22010] <= 8'h10 ;
			data[22011] <= 8'h10 ;
			data[22012] <= 8'h10 ;
			data[22013] <= 8'h10 ;
			data[22014] <= 8'h10 ;
			data[22015] <= 8'h10 ;
			data[22016] <= 8'h10 ;
			data[22017] <= 8'h10 ;
			data[22018] <= 8'h10 ;
			data[22019] <= 8'h10 ;
			data[22020] <= 8'h10 ;
			data[22021] <= 8'h10 ;
			data[22022] <= 8'h10 ;
			data[22023] <= 8'h10 ;
			data[22024] <= 8'h10 ;
			data[22025] <= 8'h10 ;
			data[22026] <= 8'h10 ;
			data[22027] <= 8'h10 ;
			data[22028] <= 8'h10 ;
			data[22029] <= 8'h10 ;
			data[22030] <= 8'h10 ;
			data[22031] <= 8'h10 ;
			data[22032] <= 8'h10 ;
			data[22033] <= 8'h10 ;
			data[22034] <= 8'h10 ;
			data[22035] <= 8'h10 ;
			data[22036] <= 8'h10 ;
			data[22037] <= 8'h10 ;
			data[22038] <= 8'h10 ;
			data[22039] <= 8'h10 ;
			data[22040] <= 8'h10 ;
			data[22041] <= 8'h10 ;
			data[22042] <= 8'h10 ;
			data[22043] <= 8'h10 ;
			data[22044] <= 8'h10 ;
			data[22045] <= 8'h10 ;
			data[22046] <= 8'h10 ;
			data[22047] <= 8'h10 ;
			data[22048] <= 8'h10 ;
			data[22049] <= 8'h10 ;
			data[22050] <= 8'h10 ;
			data[22051] <= 8'h10 ;
			data[22052] <= 8'h10 ;
			data[22053] <= 8'h10 ;
			data[22054] <= 8'h10 ;
			data[22055] <= 8'h10 ;
			data[22056] <= 8'h10 ;
			data[22057] <= 8'h10 ;
			data[22058] <= 8'h10 ;
			data[22059] <= 8'h10 ;
			data[22060] <= 8'h10 ;
			data[22061] <= 8'h10 ;
			data[22062] <= 8'h10 ;
			data[22063] <= 8'h10 ;
			data[22064] <= 8'h10 ;
			data[22065] <= 8'h10 ;
			data[22066] <= 8'h10 ;
			data[22067] <= 8'h10 ;
			data[22068] <= 8'h10 ;
			data[22069] <= 8'h10 ;
			data[22070] <= 8'h10 ;
			data[22071] <= 8'h10 ;
			data[22072] <= 8'h10 ;
			data[22073] <= 8'h10 ;
			data[22074] <= 8'h10 ;
			data[22075] <= 8'h10 ;
			data[22076] <= 8'h10 ;
			data[22077] <= 8'h10 ;
			data[22078] <= 8'h10 ;
			data[22079] <= 8'h10 ;
			data[22080] <= 8'h10 ;
			data[22081] <= 8'h10 ;
			data[22082] <= 8'h10 ;
			data[22083] <= 8'h10 ;
			data[22084] <= 8'h10 ;
			data[22085] <= 8'h10 ;
			data[22086] <= 8'h10 ;
			data[22087] <= 8'h10 ;
			data[22088] <= 8'h10 ;
			data[22089] <= 8'h10 ;
			data[22090] <= 8'h10 ;
			data[22091] <= 8'h10 ;
			data[22092] <= 8'h10 ;
			data[22093] <= 8'h10 ;
			data[22094] <= 8'h10 ;
			data[22095] <= 8'h10 ;
			data[22096] <= 8'h10 ;
			data[22097] <= 8'h10 ;
			data[22098] <= 8'h10 ;
			data[22099] <= 8'h10 ;
			data[22100] <= 8'h10 ;
			data[22101] <= 8'h10 ;
			data[22102] <= 8'h10 ;
			data[22103] <= 8'h10 ;
			data[22104] <= 8'h10 ;
			data[22105] <= 8'h10 ;
			data[22106] <= 8'h10 ;
			data[22107] <= 8'h10 ;
			data[22108] <= 8'h10 ;
			data[22109] <= 8'h10 ;
			data[22110] <= 8'h10 ;
			data[22111] <= 8'h10 ;
			data[22112] <= 8'h10 ;
			data[22113] <= 8'h10 ;
			data[22114] <= 8'h10 ;
			data[22115] <= 8'h10 ;
			data[22116] <= 8'h10 ;
			data[22117] <= 8'h10 ;
			data[22118] <= 8'h10 ;
			data[22119] <= 8'h10 ;
			data[22120] <= 8'h10 ;
			data[22121] <= 8'h10 ;
			data[22122] <= 8'h10 ;
			data[22123] <= 8'h10 ;
			data[22124] <= 8'h10 ;
			data[22125] <= 8'h10 ;
			data[22126] <= 8'h10 ;
			data[22127] <= 8'h10 ;
			data[22128] <= 8'h10 ;
			data[22129] <= 8'h10 ;
			data[22130] <= 8'h10 ;
			data[22131] <= 8'h10 ;
			data[22132] <= 8'h10 ;
			data[22133] <= 8'h10 ;
			data[22134] <= 8'h10 ;
			data[22135] <= 8'h10 ;
			data[22136] <= 8'h10 ;
			data[22137] <= 8'h10 ;
			data[22138] <= 8'h10 ;
			data[22139] <= 8'h10 ;
			data[22140] <= 8'h10 ;
			data[22141] <= 8'h10 ;
			data[22142] <= 8'h10 ;
			data[22143] <= 8'h10 ;
			data[22144] <= 8'h10 ;
			data[22145] <= 8'h10 ;
			data[22146] <= 8'h10 ;
			data[22147] <= 8'h10 ;
			data[22148] <= 8'h10 ;
			data[22149] <= 8'h10 ;
			data[22150] <= 8'h10 ;
			data[22151] <= 8'h10 ;
			data[22152] <= 8'h10 ;
			data[22153] <= 8'h10 ;
			data[22154] <= 8'h10 ;
			data[22155] <= 8'h10 ;
			data[22156] <= 8'h10 ;
			data[22157] <= 8'h10 ;
			data[22158] <= 8'h10 ;
			data[22159] <= 8'h10 ;
			data[22160] <= 8'h10 ;
			data[22161] <= 8'h10 ;
			data[22162] <= 8'h10 ;
			data[22163] <= 8'h10 ;
			data[22164] <= 8'h10 ;
			data[22165] <= 8'h10 ;
			data[22166] <= 8'h10 ;
			data[22167] <= 8'h10 ;
			data[22168] <= 8'h10 ;
			data[22169] <= 8'h10 ;
			data[22170] <= 8'h10 ;
			data[22171] <= 8'h10 ;
			data[22172] <= 8'h10 ;
			data[22173] <= 8'h10 ;
			data[22174] <= 8'h10 ;
			data[22175] <= 8'h10 ;
			data[22176] <= 8'h10 ;
			data[22177] <= 8'h10 ;
			data[22178] <= 8'h10 ;
			data[22179] <= 8'h10 ;
			data[22180] <= 8'h10 ;
			data[22181] <= 8'h10 ;
			data[22182] <= 8'h10 ;
			data[22183] <= 8'h10 ;
			data[22184] <= 8'h10 ;
			data[22185] <= 8'h10 ;
			data[22186] <= 8'h10 ;
			data[22187] <= 8'h10 ;
			data[22188] <= 8'h10 ;
			data[22189] <= 8'h10 ;
			data[22190] <= 8'h10 ;
			data[22191] <= 8'h10 ;
			data[22192] <= 8'h10 ;
			data[22193] <= 8'h10 ;
			data[22194] <= 8'h10 ;
			data[22195] <= 8'h10 ;
			data[22196] <= 8'h10 ;
			data[22197] <= 8'h10 ;
			data[22198] <= 8'h10 ;
			data[22199] <= 8'h10 ;
			data[22200] <= 8'h10 ;
			data[22201] <= 8'h10 ;
			data[22202] <= 8'h10 ;
			data[22203] <= 8'h10 ;
			data[22204] <= 8'h10 ;
			data[22205] <= 8'h10 ;
			data[22206] <= 8'h10 ;
			data[22207] <= 8'h10 ;
			data[22208] <= 8'h10 ;
			data[22209] <= 8'h10 ;
			data[22210] <= 8'h10 ;
			data[22211] <= 8'h10 ;
			data[22212] <= 8'h10 ;
			data[22213] <= 8'h10 ;
			data[22214] <= 8'h10 ;
			data[22215] <= 8'h10 ;
			data[22216] <= 8'h10 ;
			data[22217] <= 8'h10 ;
			data[22218] <= 8'h10 ;
			data[22219] <= 8'h10 ;
			data[22220] <= 8'h10 ;
			data[22221] <= 8'h10 ;
			data[22222] <= 8'h10 ;
			data[22223] <= 8'h10 ;
			data[22224] <= 8'h10 ;
			data[22225] <= 8'h10 ;
			data[22226] <= 8'h10 ;
			data[22227] <= 8'h10 ;
			data[22228] <= 8'h10 ;
			data[22229] <= 8'h10 ;
			data[22230] <= 8'h10 ;
			data[22231] <= 8'h10 ;
			data[22232] <= 8'h10 ;
			data[22233] <= 8'h10 ;
			data[22234] <= 8'h10 ;
			data[22235] <= 8'h10 ;
			data[22236] <= 8'h10 ;
			data[22237] <= 8'h10 ;
			data[22238] <= 8'h10 ;
			data[22239] <= 8'h10 ;
			data[22240] <= 8'h10 ;
			data[22241] <= 8'h10 ;
			data[22242] <= 8'h10 ;
			data[22243] <= 8'h10 ;
			data[22244] <= 8'h10 ;
			data[22245] <= 8'h10 ;
			data[22246] <= 8'h10 ;
			data[22247] <= 8'h10 ;
			data[22248] <= 8'h10 ;
			data[22249] <= 8'h10 ;
			data[22250] <= 8'h10 ;
			data[22251] <= 8'h10 ;
			data[22252] <= 8'h10 ;
			data[22253] <= 8'h10 ;
			data[22254] <= 8'h10 ;
			data[22255] <= 8'h10 ;
			data[22256] <= 8'h10 ;
			data[22257] <= 8'h10 ;
			data[22258] <= 8'h10 ;
			data[22259] <= 8'h10 ;
			data[22260] <= 8'h10 ;
			data[22261] <= 8'h10 ;
			data[22262] <= 8'h10 ;
			data[22263] <= 8'h10 ;
			data[22264] <= 8'h10 ;
			data[22265] <= 8'h10 ;
			data[22266] <= 8'h10 ;
			data[22267] <= 8'h10 ;
			data[22268] <= 8'h10 ;
			data[22269] <= 8'h10 ;
			data[22270] <= 8'h10 ;
			data[22271] <= 8'h10 ;
			data[22272] <= 8'h10 ;
			data[22273] <= 8'h10 ;
			data[22274] <= 8'h10 ;
			data[22275] <= 8'h10 ;
			data[22276] <= 8'h10 ;
			data[22277] <= 8'h10 ;
			data[22278] <= 8'h10 ;
			data[22279] <= 8'h10 ;
			data[22280] <= 8'h10 ;
			data[22281] <= 8'h10 ;
			data[22282] <= 8'h10 ;
			data[22283] <= 8'h10 ;
			data[22284] <= 8'h10 ;
			data[22285] <= 8'h10 ;
			data[22286] <= 8'h10 ;
			data[22287] <= 8'h10 ;
			data[22288] <= 8'h10 ;
			data[22289] <= 8'h10 ;
			data[22290] <= 8'h10 ;
			data[22291] <= 8'h10 ;
			data[22292] <= 8'h10 ;
			data[22293] <= 8'h10 ;
			data[22294] <= 8'h10 ;
			data[22295] <= 8'h10 ;
			data[22296] <= 8'h10 ;
			data[22297] <= 8'h10 ;
			data[22298] <= 8'h10 ;
			data[22299] <= 8'h10 ;
			data[22300] <= 8'h10 ;
			data[22301] <= 8'h10 ;
			data[22302] <= 8'h10 ;
			data[22303] <= 8'h10 ;
			data[22304] <= 8'h10 ;
			data[22305] <= 8'h10 ;
			data[22306] <= 8'h10 ;
			data[22307] <= 8'h10 ;
			data[22308] <= 8'h10 ;
			data[22309] <= 8'h10 ;
			data[22310] <= 8'h10 ;
			data[22311] <= 8'h10 ;
			data[22312] <= 8'h10 ;
			data[22313] <= 8'h10 ;
			data[22314] <= 8'h10 ;
			data[22315] <= 8'h10 ;
			data[22316] <= 8'h10 ;
			data[22317] <= 8'h10 ;
			data[22318] <= 8'h10 ;
			data[22319] <= 8'h10 ;
			data[22320] <= 8'h10 ;
			data[22321] <= 8'h10 ;
			data[22322] <= 8'h10 ;
			data[22323] <= 8'h10 ;
			data[22324] <= 8'h10 ;
			data[22325] <= 8'h10 ;
			data[22326] <= 8'h10 ;
			data[22327] <= 8'h10 ;
			data[22328] <= 8'h10 ;
			data[22329] <= 8'h10 ;
			data[22330] <= 8'h10 ;
			data[22331] <= 8'h10 ;
			data[22332] <= 8'h10 ;
			data[22333] <= 8'h10 ;
			data[22334] <= 8'h10 ;
			data[22335] <= 8'h10 ;
			data[22336] <= 8'h10 ;
			data[22337] <= 8'h10 ;
			data[22338] <= 8'h10 ;
			data[22339] <= 8'h10 ;
			data[22340] <= 8'h10 ;
			data[22341] <= 8'h10 ;
			data[22342] <= 8'h10 ;
			data[22343] <= 8'h10 ;
			data[22344] <= 8'h10 ;
			data[22345] <= 8'h10 ;
			data[22346] <= 8'h10 ;
			data[22347] <= 8'h10 ;
			data[22348] <= 8'h10 ;
			data[22349] <= 8'h10 ;
			data[22350] <= 8'h10 ;
			data[22351] <= 8'h10 ;
			data[22352] <= 8'h10 ;
			data[22353] <= 8'h10 ;
			data[22354] <= 8'h10 ;
			data[22355] <= 8'h10 ;
			data[22356] <= 8'h10 ;
			data[22357] <= 8'h10 ;
			data[22358] <= 8'h10 ;
			data[22359] <= 8'h10 ;
			data[22360] <= 8'h10 ;
			data[22361] <= 8'h10 ;
			data[22362] <= 8'h10 ;
			data[22363] <= 8'h10 ;
			data[22364] <= 8'h10 ;
			data[22365] <= 8'h10 ;
			data[22366] <= 8'h10 ;
			data[22367] <= 8'h10 ;
			data[22368] <= 8'h10 ;
			data[22369] <= 8'h10 ;
			data[22370] <= 8'h10 ;
			data[22371] <= 8'h10 ;
			data[22372] <= 8'h10 ;
			data[22373] <= 8'h10 ;
			data[22374] <= 8'h10 ;
			data[22375] <= 8'h10 ;
			data[22376] <= 8'h10 ;
			data[22377] <= 8'h10 ;
			data[22378] <= 8'h10 ;
			data[22379] <= 8'h10 ;
			data[22380] <= 8'h10 ;
			data[22381] <= 8'h10 ;
			data[22382] <= 8'h10 ;
			data[22383] <= 8'h10 ;
			data[22384] <= 8'h10 ;
			data[22385] <= 8'h10 ;
			data[22386] <= 8'h10 ;
			data[22387] <= 8'h10 ;
			data[22388] <= 8'h10 ;
			data[22389] <= 8'h10 ;
			data[22390] <= 8'h10 ;
			data[22391] <= 8'h10 ;
			data[22392] <= 8'h10 ;
			data[22393] <= 8'h10 ;
			data[22394] <= 8'h10 ;
			data[22395] <= 8'h10 ;
			data[22396] <= 8'h10 ;
			data[22397] <= 8'h10 ;
			data[22398] <= 8'h10 ;
			data[22399] <= 8'h10 ;
			data[22400] <= 8'h10 ;
			data[22401] <= 8'h10 ;
			data[22402] <= 8'h10 ;
			data[22403] <= 8'h10 ;
			data[22404] <= 8'h10 ;
			data[22405] <= 8'h10 ;
			data[22406] <= 8'h10 ;
			data[22407] <= 8'h10 ;
			data[22408] <= 8'h10 ;
			data[22409] <= 8'h10 ;
			data[22410] <= 8'h10 ;
			data[22411] <= 8'h10 ;
			data[22412] <= 8'h10 ;
			data[22413] <= 8'h10 ;
			data[22414] <= 8'h10 ;
			data[22415] <= 8'h10 ;
			data[22416] <= 8'h10 ;
			data[22417] <= 8'h10 ;
			data[22418] <= 8'h10 ;
			data[22419] <= 8'h10 ;
			data[22420] <= 8'h10 ;
			data[22421] <= 8'h10 ;
			data[22422] <= 8'h10 ;
			data[22423] <= 8'h10 ;
			data[22424] <= 8'h10 ;
			data[22425] <= 8'h10 ;
			data[22426] <= 8'h10 ;
			data[22427] <= 8'h10 ;
			data[22428] <= 8'h10 ;
			data[22429] <= 8'h10 ;
			data[22430] <= 8'h10 ;
			data[22431] <= 8'h10 ;
			data[22432] <= 8'h10 ;
			data[22433] <= 8'h10 ;
			data[22434] <= 8'h10 ;
			data[22435] <= 8'h10 ;
			data[22436] <= 8'h10 ;
			data[22437] <= 8'h10 ;
			data[22438] <= 8'h10 ;
			data[22439] <= 8'h10 ;
			data[22440] <= 8'h10 ;
			data[22441] <= 8'h10 ;
			data[22442] <= 8'h10 ;
			data[22443] <= 8'h10 ;
			data[22444] <= 8'h10 ;
			data[22445] <= 8'h10 ;
			data[22446] <= 8'h10 ;
			data[22447] <= 8'h10 ;
			data[22448] <= 8'h10 ;
			data[22449] <= 8'h10 ;
			data[22450] <= 8'h10 ;
			data[22451] <= 8'h10 ;
			data[22452] <= 8'h10 ;
			data[22453] <= 8'h10 ;
			data[22454] <= 8'h10 ;
			data[22455] <= 8'h10 ;
			data[22456] <= 8'h10 ;
			data[22457] <= 8'h10 ;
			data[22458] <= 8'h10 ;
			data[22459] <= 8'h10 ;
			data[22460] <= 8'h10 ;
			data[22461] <= 8'h10 ;
			data[22462] <= 8'h10 ;
			data[22463] <= 8'h10 ;
			data[22464] <= 8'h10 ;
			data[22465] <= 8'h10 ;
			data[22466] <= 8'h10 ;
			data[22467] <= 8'h10 ;
			data[22468] <= 8'h10 ;
			data[22469] <= 8'h10 ;
			data[22470] <= 8'h10 ;
			data[22471] <= 8'h10 ;
			data[22472] <= 8'h10 ;
			data[22473] <= 8'h10 ;
			data[22474] <= 8'h10 ;
			data[22475] <= 8'h10 ;
			data[22476] <= 8'h10 ;
			data[22477] <= 8'h10 ;
			data[22478] <= 8'h10 ;
			data[22479] <= 8'h10 ;
			data[22480] <= 8'h10 ;
			data[22481] <= 8'h10 ;
			data[22482] <= 8'h10 ;
			data[22483] <= 8'h10 ;
			data[22484] <= 8'h10 ;
			data[22485] <= 8'h10 ;
			data[22486] <= 8'h10 ;
			data[22487] <= 8'h10 ;
			data[22488] <= 8'h10 ;
			data[22489] <= 8'h10 ;
			data[22490] <= 8'h10 ;
			data[22491] <= 8'h10 ;
			data[22492] <= 8'h10 ;
			data[22493] <= 8'h10 ;
			data[22494] <= 8'h10 ;
			data[22495] <= 8'h10 ;
			data[22496] <= 8'h10 ;
			data[22497] <= 8'h10 ;
			data[22498] <= 8'h10 ;
			data[22499] <= 8'h10 ;
			data[22500] <= 8'h10 ;
			data[22501] <= 8'h10 ;
			data[22502] <= 8'h10 ;
			data[22503] <= 8'h10 ;
			data[22504] <= 8'h10 ;
			data[22505] <= 8'h10 ;
			data[22506] <= 8'h10 ;
			data[22507] <= 8'h10 ;
			data[22508] <= 8'h10 ;
			data[22509] <= 8'h10 ;
			data[22510] <= 8'h10 ;
			data[22511] <= 8'h10 ;
			data[22512] <= 8'h10 ;
			data[22513] <= 8'h10 ;
			data[22514] <= 8'h10 ;
			data[22515] <= 8'h10 ;
			data[22516] <= 8'h10 ;
			data[22517] <= 8'h10 ;
			data[22518] <= 8'h10 ;
			data[22519] <= 8'h10 ;
			data[22520] <= 8'h10 ;
			data[22521] <= 8'h10 ;
			data[22522] <= 8'h10 ;
			data[22523] <= 8'h10 ;
			data[22524] <= 8'h10 ;
			data[22525] <= 8'h10 ;
			data[22526] <= 8'h10 ;
			data[22527] <= 8'h10 ;
			data[22528] <= 8'h10 ;
			data[22529] <= 8'h10 ;
			data[22530] <= 8'h10 ;
			data[22531] <= 8'h10 ;
			data[22532] <= 8'h10 ;
			data[22533] <= 8'h10 ;
			data[22534] <= 8'h10 ;
			data[22535] <= 8'h10 ;
			data[22536] <= 8'h10 ;
			data[22537] <= 8'h10 ;
			data[22538] <= 8'h10 ;
			data[22539] <= 8'h10 ;
			data[22540] <= 8'h10 ;
			data[22541] <= 8'h10 ;
			data[22542] <= 8'h10 ;
			data[22543] <= 8'h10 ;
			data[22544] <= 8'h10 ;
			data[22545] <= 8'h10 ;
			data[22546] <= 8'h10 ;
			data[22547] <= 8'h10 ;
			data[22548] <= 8'h10 ;
			data[22549] <= 8'h10 ;
			data[22550] <= 8'h10 ;
			data[22551] <= 8'h10 ;
			data[22552] <= 8'h10 ;
			data[22553] <= 8'h10 ;
			data[22554] <= 8'h10 ;
			data[22555] <= 8'h10 ;
			data[22556] <= 8'h10 ;
			data[22557] <= 8'h10 ;
			data[22558] <= 8'h10 ;
			data[22559] <= 8'h10 ;
			data[22560] <= 8'h10 ;
			data[22561] <= 8'h10 ;
			data[22562] <= 8'h10 ;
			data[22563] <= 8'h10 ;
			data[22564] <= 8'h10 ;
			data[22565] <= 8'h10 ;
			data[22566] <= 8'h10 ;
			data[22567] <= 8'h10 ;
			data[22568] <= 8'h10 ;
			data[22569] <= 8'h10 ;
			data[22570] <= 8'h10 ;
			data[22571] <= 8'h10 ;
			data[22572] <= 8'h10 ;
			data[22573] <= 8'h10 ;
			data[22574] <= 8'h10 ;
			data[22575] <= 8'h10 ;
			data[22576] <= 8'h10 ;
			data[22577] <= 8'h10 ;
			data[22578] <= 8'h10 ;
			data[22579] <= 8'h10 ;
			data[22580] <= 8'h10 ;
			data[22581] <= 8'h10 ;
			data[22582] <= 8'h10 ;
			data[22583] <= 8'h10 ;
			data[22584] <= 8'h10 ;
			data[22585] <= 8'h10 ;
			data[22586] <= 8'h10 ;
			data[22587] <= 8'h10 ;
			data[22588] <= 8'h10 ;
			data[22589] <= 8'h10 ;
			data[22590] <= 8'h10 ;
			data[22591] <= 8'h10 ;
			data[22592] <= 8'h10 ;
			data[22593] <= 8'h10 ;
			data[22594] <= 8'h10 ;
			data[22595] <= 8'h10 ;
			data[22596] <= 8'h10 ;
			data[22597] <= 8'h10 ;
			data[22598] <= 8'h10 ;
			data[22599] <= 8'h10 ;
			data[22600] <= 8'h10 ;
			data[22601] <= 8'h10 ;
			data[22602] <= 8'h10 ;
			data[22603] <= 8'h10 ;
			data[22604] <= 8'h10 ;
			data[22605] <= 8'h10 ;
			data[22606] <= 8'h10 ;
			data[22607] <= 8'h10 ;
			data[22608] <= 8'h10 ;
			data[22609] <= 8'h10 ;
			data[22610] <= 8'h10 ;
			data[22611] <= 8'h10 ;
			data[22612] <= 8'h10 ;
			data[22613] <= 8'h10 ;
			data[22614] <= 8'h10 ;
			data[22615] <= 8'h10 ;
			data[22616] <= 8'h10 ;
			data[22617] <= 8'h10 ;
			data[22618] <= 8'h10 ;
			data[22619] <= 8'h10 ;
			data[22620] <= 8'h10 ;
			data[22621] <= 8'h10 ;
			data[22622] <= 8'h10 ;
			data[22623] <= 8'h10 ;
			data[22624] <= 8'h10 ;
			data[22625] <= 8'h10 ;
			data[22626] <= 8'h10 ;
			data[22627] <= 8'h10 ;
			data[22628] <= 8'h10 ;
			data[22629] <= 8'h10 ;
			data[22630] <= 8'h10 ;
			data[22631] <= 8'h10 ;
			data[22632] <= 8'h10 ;
			data[22633] <= 8'h10 ;
			data[22634] <= 8'h10 ;
			data[22635] <= 8'h10 ;
			data[22636] <= 8'h10 ;
			data[22637] <= 8'h10 ;
			data[22638] <= 8'h10 ;
			data[22639] <= 8'h10 ;
			data[22640] <= 8'h10 ;
			data[22641] <= 8'h10 ;
			data[22642] <= 8'h10 ;
			data[22643] <= 8'h10 ;
			data[22644] <= 8'h10 ;
			data[22645] <= 8'h10 ;
			data[22646] <= 8'h10 ;
			data[22647] <= 8'h10 ;
			data[22648] <= 8'h10 ;
			data[22649] <= 8'h10 ;
			data[22650] <= 8'h10 ;
			data[22651] <= 8'h10 ;
			data[22652] <= 8'h10 ;
			data[22653] <= 8'h10 ;
			data[22654] <= 8'h10 ;
			data[22655] <= 8'h10 ;
			data[22656] <= 8'h10 ;
			data[22657] <= 8'h10 ;
			data[22658] <= 8'h10 ;
			data[22659] <= 8'h10 ;
			data[22660] <= 8'h10 ;
			data[22661] <= 8'h10 ;
			data[22662] <= 8'h10 ;
			data[22663] <= 8'h10 ;
			data[22664] <= 8'h10 ;
			data[22665] <= 8'h10 ;
			data[22666] <= 8'h10 ;
			data[22667] <= 8'h10 ;
			data[22668] <= 8'h10 ;
			data[22669] <= 8'h10 ;
			data[22670] <= 8'h10 ;
			data[22671] <= 8'h10 ;
			data[22672] <= 8'h10 ;
			data[22673] <= 8'h10 ;
			data[22674] <= 8'h10 ;
			data[22675] <= 8'h10 ;
			data[22676] <= 8'h10 ;
			data[22677] <= 8'h10 ;
			data[22678] <= 8'h10 ;
			data[22679] <= 8'h10 ;
			data[22680] <= 8'h10 ;
			data[22681] <= 8'h10 ;
			data[22682] <= 8'h10 ;
			data[22683] <= 8'h10 ;
			data[22684] <= 8'h10 ;
			data[22685] <= 8'h10 ;
			data[22686] <= 8'h10 ;
			data[22687] <= 8'h10 ;
			data[22688] <= 8'h10 ;
			data[22689] <= 8'h10 ;
			data[22690] <= 8'h10 ;
			data[22691] <= 8'h10 ;
			data[22692] <= 8'h10 ;
			data[22693] <= 8'h10 ;
			data[22694] <= 8'h10 ;
			data[22695] <= 8'h10 ;
			data[22696] <= 8'h10 ;
			data[22697] <= 8'h10 ;
			data[22698] <= 8'h10 ;
			data[22699] <= 8'h10 ;
			data[22700] <= 8'h10 ;
			data[22701] <= 8'h10 ;
			data[22702] <= 8'h10 ;
			data[22703] <= 8'h10 ;
			data[22704] <= 8'h10 ;
			data[22705] <= 8'h10 ;
			data[22706] <= 8'h10 ;
			data[22707] <= 8'h10 ;
			data[22708] <= 8'h10 ;
			data[22709] <= 8'h10 ;
			data[22710] <= 8'h10 ;
			data[22711] <= 8'h10 ;
			data[22712] <= 8'h10 ;
			data[22713] <= 8'h10 ;
			data[22714] <= 8'h10 ;
			data[22715] <= 8'h10 ;
			data[22716] <= 8'h10 ;
			data[22717] <= 8'h10 ;
			data[22718] <= 8'h10 ;
			data[22719] <= 8'h10 ;
			data[22720] <= 8'h10 ;
			data[22721] <= 8'h10 ;
			data[22722] <= 8'h10 ;
			data[22723] <= 8'h10 ;
			data[22724] <= 8'h10 ;
			data[22725] <= 8'h10 ;
			data[22726] <= 8'h10 ;
			data[22727] <= 8'h10 ;
			data[22728] <= 8'h10 ;
			data[22729] <= 8'h10 ;
			data[22730] <= 8'h10 ;
			data[22731] <= 8'h10 ;
			data[22732] <= 8'h10 ;
			data[22733] <= 8'h10 ;
			data[22734] <= 8'h10 ;
			data[22735] <= 8'h10 ;
			data[22736] <= 8'h10 ;
			data[22737] <= 8'h10 ;
			data[22738] <= 8'h10 ;
			data[22739] <= 8'h10 ;
			data[22740] <= 8'h10 ;
			data[22741] <= 8'h10 ;
			data[22742] <= 8'h10 ;
			data[22743] <= 8'h10 ;
			data[22744] <= 8'h10 ;
			data[22745] <= 8'h10 ;
			data[22746] <= 8'h10 ;
			data[22747] <= 8'h10 ;
			data[22748] <= 8'h10 ;
			data[22749] <= 8'h10 ;
			data[22750] <= 8'h10 ;
			data[22751] <= 8'h10 ;
			data[22752] <= 8'h10 ;
			data[22753] <= 8'h10 ;
			data[22754] <= 8'h10 ;
			data[22755] <= 8'h10 ;
			data[22756] <= 8'h10 ;
			data[22757] <= 8'h10 ;
			data[22758] <= 8'h10 ;
			data[22759] <= 8'h10 ;
			data[22760] <= 8'h10 ;
			data[22761] <= 8'h10 ;
			data[22762] <= 8'h10 ;
			data[22763] <= 8'h10 ;
			data[22764] <= 8'h10 ;
			data[22765] <= 8'h10 ;
			data[22766] <= 8'h10 ;
			data[22767] <= 8'h10 ;
			data[22768] <= 8'h10 ;
			data[22769] <= 8'h10 ;
			data[22770] <= 8'h10 ;
			data[22771] <= 8'h10 ;
			data[22772] <= 8'h10 ;
			data[22773] <= 8'h10 ;
			data[22774] <= 8'h10 ;
			data[22775] <= 8'h10 ;
			data[22776] <= 8'h10 ;
			data[22777] <= 8'h10 ;
			data[22778] <= 8'h10 ;
			data[22779] <= 8'h10 ;
			data[22780] <= 8'h10 ;
			data[22781] <= 8'h10 ;
			data[22782] <= 8'h10 ;
			data[22783] <= 8'h10 ;
			data[22784] <= 8'h10 ;
			data[22785] <= 8'h10 ;
			data[22786] <= 8'h10 ;
			data[22787] <= 8'h10 ;
			data[22788] <= 8'h10 ;
			data[22789] <= 8'h10 ;
			data[22790] <= 8'h10 ;
			data[22791] <= 8'h10 ;
			data[22792] <= 8'h10 ;
			data[22793] <= 8'h10 ;
			data[22794] <= 8'h10 ;
			data[22795] <= 8'h10 ;
			data[22796] <= 8'h10 ;
			data[22797] <= 8'h10 ;
			data[22798] <= 8'h10 ;
			data[22799] <= 8'h10 ;
			data[22800] <= 8'h10 ;
			data[22801] <= 8'h10 ;
			data[22802] <= 8'h10 ;
			data[22803] <= 8'h10 ;
			data[22804] <= 8'h10 ;
			data[22805] <= 8'h10 ;
			data[22806] <= 8'h10 ;
			data[22807] <= 8'h10 ;
			data[22808] <= 8'h10 ;
			data[22809] <= 8'h10 ;
			data[22810] <= 8'h10 ;
			data[22811] <= 8'h10 ;
			data[22812] <= 8'h10 ;
			data[22813] <= 8'h10 ;
			data[22814] <= 8'h10 ;
			data[22815] <= 8'h10 ;
			data[22816] <= 8'h10 ;
			data[22817] <= 8'h10 ;
			data[22818] <= 8'h10 ;
			data[22819] <= 8'h10 ;
			data[22820] <= 8'h10 ;
			data[22821] <= 8'h10 ;
			data[22822] <= 8'h10 ;
			data[22823] <= 8'h10 ;
			data[22824] <= 8'h10 ;
			data[22825] <= 8'h10 ;
			data[22826] <= 8'h10 ;
			data[22827] <= 8'h10 ;
			data[22828] <= 8'h10 ;
			data[22829] <= 8'h10 ;
			data[22830] <= 8'h10 ;
			data[22831] <= 8'h10 ;
			data[22832] <= 8'h10 ;
			data[22833] <= 8'h10 ;
			data[22834] <= 8'h10 ;
			data[22835] <= 8'h10 ;
			data[22836] <= 8'h10 ;
			data[22837] <= 8'h10 ;
			data[22838] <= 8'h10 ;
			data[22839] <= 8'h10 ;
			data[22840] <= 8'h10 ;
			data[22841] <= 8'h10 ;
			data[22842] <= 8'h10 ;
			data[22843] <= 8'h10 ;
			data[22844] <= 8'h10 ;
			data[22845] <= 8'h10 ;
			data[22846] <= 8'h10 ;
			data[22847] <= 8'h10 ;
			data[22848] <= 8'h10 ;
			data[22849] <= 8'h10 ;
			data[22850] <= 8'h10 ;
			data[22851] <= 8'h10 ;
			data[22852] <= 8'h10 ;
			data[22853] <= 8'h10 ;
			data[22854] <= 8'h10 ;
			data[22855] <= 8'h10 ;
			data[22856] <= 8'h10 ;
			data[22857] <= 8'h10 ;
			data[22858] <= 8'h10 ;
			data[22859] <= 8'h10 ;
			data[22860] <= 8'h10 ;
			data[22861] <= 8'h10 ;
			data[22862] <= 8'h10 ;
			data[22863] <= 8'h10 ;
			data[22864] <= 8'h10 ;
			data[22865] <= 8'h10 ;
			data[22866] <= 8'h10 ;
			data[22867] <= 8'h10 ;
			data[22868] <= 8'h10 ;
			data[22869] <= 8'h10 ;
			data[22870] <= 8'h10 ;
			data[22871] <= 8'h10 ;
			data[22872] <= 8'h10 ;
			data[22873] <= 8'h10 ;
			data[22874] <= 8'h10 ;
			data[22875] <= 8'h10 ;
			data[22876] <= 8'h10 ;
			data[22877] <= 8'h10 ;
			data[22878] <= 8'h10 ;
			data[22879] <= 8'h10 ;
			data[22880] <= 8'h10 ;
			data[22881] <= 8'h10 ;
			data[22882] <= 8'h10 ;
			data[22883] <= 8'h10 ;
			data[22884] <= 8'h10 ;
			data[22885] <= 8'h10 ;
			data[22886] <= 8'h10 ;
			data[22887] <= 8'h10 ;
			data[22888] <= 8'h10 ;
			data[22889] <= 8'h10 ;
			data[22890] <= 8'h10 ;
			data[22891] <= 8'h10 ;
			data[22892] <= 8'h10 ;
			data[22893] <= 8'h10 ;
			data[22894] <= 8'h10 ;
			data[22895] <= 8'h10 ;
			data[22896] <= 8'h10 ;
			data[22897] <= 8'h10 ;
			data[22898] <= 8'h10 ;
			data[22899] <= 8'h10 ;
			data[22900] <= 8'h10 ;
			data[22901] <= 8'h10 ;
			data[22902] <= 8'h10 ;
			data[22903] <= 8'h10 ;
			data[22904] <= 8'h10 ;
			data[22905] <= 8'h10 ;
			data[22906] <= 8'h10 ;
			data[22907] <= 8'h10 ;
			data[22908] <= 8'h10 ;
			data[22909] <= 8'h10 ;
			data[22910] <= 8'h10 ;
			data[22911] <= 8'h10 ;
			data[22912] <= 8'h10 ;
			data[22913] <= 8'h10 ;
			data[22914] <= 8'h10 ;
			data[22915] <= 8'h10 ;
			data[22916] <= 8'h10 ;
			data[22917] <= 8'h10 ;
			data[22918] <= 8'h10 ;
			data[22919] <= 8'h10 ;
			data[22920] <= 8'h10 ;
			data[22921] <= 8'h10 ;
			data[22922] <= 8'h10 ;
			data[22923] <= 8'h10 ;
			data[22924] <= 8'h10 ;
			data[22925] <= 8'h10 ;
			data[22926] <= 8'h10 ;
			data[22927] <= 8'h10 ;
			data[22928] <= 8'h10 ;
			data[22929] <= 8'h10 ;
			data[22930] <= 8'h10 ;
			data[22931] <= 8'h10 ;
			data[22932] <= 8'h10 ;
			data[22933] <= 8'h10 ;
			data[22934] <= 8'h10 ;
			data[22935] <= 8'h10 ;
			data[22936] <= 8'h10 ;
			data[22937] <= 8'h10 ;
			data[22938] <= 8'h10 ;
			data[22939] <= 8'h10 ;
			data[22940] <= 8'h10 ;
			data[22941] <= 8'h10 ;
			data[22942] <= 8'h10 ;
			data[22943] <= 8'h10 ;
			data[22944] <= 8'h10 ;
			data[22945] <= 8'h10 ;
			data[22946] <= 8'h10 ;
			data[22947] <= 8'h10 ;
			data[22948] <= 8'h10 ;
			data[22949] <= 8'h10 ;
			data[22950] <= 8'h10 ;
			data[22951] <= 8'h10 ;
			data[22952] <= 8'h10 ;
			data[22953] <= 8'h10 ;
			data[22954] <= 8'h10 ;
			data[22955] <= 8'h10 ;
			data[22956] <= 8'h10 ;
			data[22957] <= 8'h10 ;
			data[22958] <= 8'h10 ;
			data[22959] <= 8'h10 ;
			data[22960] <= 8'h10 ;
			data[22961] <= 8'h10 ;
			data[22962] <= 8'h10 ;
			data[22963] <= 8'h10 ;
			data[22964] <= 8'h10 ;
			data[22965] <= 8'h10 ;
			data[22966] <= 8'h10 ;
			data[22967] <= 8'h10 ;
			data[22968] <= 8'h10 ;
			data[22969] <= 8'h10 ;
			data[22970] <= 8'h10 ;
			data[22971] <= 8'h10 ;
			data[22972] <= 8'h10 ;
			data[22973] <= 8'h10 ;
			data[22974] <= 8'h10 ;
			data[22975] <= 8'h10 ;
			data[22976] <= 8'h10 ;
			data[22977] <= 8'h10 ;
			data[22978] <= 8'h10 ;
			data[22979] <= 8'h10 ;
			data[22980] <= 8'h10 ;
			data[22981] <= 8'h10 ;
			data[22982] <= 8'h10 ;
			data[22983] <= 8'h10 ;
			data[22984] <= 8'h10 ;
			data[22985] <= 8'h10 ;
			data[22986] <= 8'h10 ;
			data[22987] <= 8'h10 ;
			data[22988] <= 8'h10 ;
			data[22989] <= 8'h10 ;
			data[22990] <= 8'h10 ;
			data[22991] <= 8'h10 ;
			data[22992] <= 8'h10 ;
			data[22993] <= 8'h10 ;
			data[22994] <= 8'h10 ;
			data[22995] <= 8'h10 ;
			data[22996] <= 8'h10 ;
			data[22997] <= 8'h10 ;
			data[22998] <= 8'h10 ;
			data[22999] <= 8'h10 ;
			data[23000] <= 8'h10 ;
			data[23001] <= 8'h10 ;
			data[23002] <= 8'h10 ;
			data[23003] <= 8'h10 ;
			data[23004] <= 8'h10 ;
			data[23005] <= 8'h10 ;
			data[23006] <= 8'h10 ;
			data[23007] <= 8'h10 ;
			data[23008] <= 8'h10 ;
			data[23009] <= 8'h10 ;
			data[23010] <= 8'h10 ;
			data[23011] <= 8'h10 ;
			data[23012] <= 8'h10 ;
			data[23013] <= 8'h10 ;
			data[23014] <= 8'h10 ;
			data[23015] <= 8'h10 ;
			data[23016] <= 8'h10 ;
			data[23017] <= 8'h10 ;
			data[23018] <= 8'h10 ;
			data[23019] <= 8'h10 ;
			data[23020] <= 8'h10 ;
			data[23021] <= 8'h10 ;
			data[23022] <= 8'h10 ;
			data[23023] <= 8'h10 ;
			data[23024] <= 8'h10 ;
			data[23025] <= 8'h10 ;
			data[23026] <= 8'h10 ;
			data[23027] <= 8'h10 ;
			data[23028] <= 8'h10 ;
			data[23029] <= 8'h10 ;
			data[23030] <= 8'h10 ;
			data[23031] <= 8'h10 ;
			data[23032] <= 8'h10 ;
			data[23033] <= 8'h10 ;
			data[23034] <= 8'h10 ;
			data[23035] <= 8'h10 ;
			data[23036] <= 8'h10 ;
			data[23037] <= 8'h10 ;
			data[23038] <= 8'h10 ;
			data[23039] <= 8'h10 ;
			data[23040] <= 8'h10 ;
			data[23041] <= 8'h10 ;
			data[23042] <= 8'h10 ;
			data[23043] <= 8'h10 ;
			data[23044] <= 8'h10 ;
			data[23045] <= 8'h10 ;
			data[23046] <= 8'h10 ;
			data[23047] <= 8'h10 ;
			data[23048] <= 8'h10 ;
			data[23049] <= 8'h10 ;
			data[23050] <= 8'h10 ;
			data[23051] <= 8'h10 ;
			data[23052] <= 8'h10 ;
			data[23053] <= 8'h10 ;
			data[23054] <= 8'h10 ;
			data[23055] <= 8'h10 ;
			data[23056] <= 8'h10 ;
			data[23057] <= 8'h10 ;
			data[23058] <= 8'h10 ;
			data[23059] <= 8'h10 ;
			data[23060] <= 8'h10 ;
			data[23061] <= 8'h10 ;
			data[23062] <= 8'h10 ;
			data[23063] <= 8'h10 ;
			data[23064] <= 8'h10 ;
			data[23065] <= 8'h10 ;
			data[23066] <= 8'h10 ;
			data[23067] <= 8'h10 ;
			data[23068] <= 8'h10 ;
			data[23069] <= 8'h10 ;
			data[23070] <= 8'h10 ;
			data[23071] <= 8'h10 ;
			data[23072] <= 8'h10 ;
			data[23073] <= 8'h10 ;
			data[23074] <= 8'h10 ;
			data[23075] <= 8'h10 ;
			data[23076] <= 8'h10 ;
			data[23077] <= 8'h10 ;
			data[23078] <= 8'h10 ;
			data[23079] <= 8'h10 ;
			data[23080] <= 8'h10 ;
			data[23081] <= 8'h10 ;
			data[23082] <= 8'h10 ;
			data[23083] <= 8'h10 ;
			data[23084] <= 8'h10 ;
			data[23085] <= 8'h10 ;
			data[23086] <= 8'h10 ;
			data[23087] <= 8'h10 ;
			data[23088] <= 8'h10 ;
			data[23089] <= 8'h10 ;
			data[23090] <= 8'h10 ;
			data[23091] <= 8'h10 ;
			data[23092] <= 8'h10 ;
			data[23093] <= 8'h10 ;
			data[23094] <= 8'h10 ;
			data[23095] <= 8'h10 ;
			data[23096] <= 8'h10 ;
			data[23097] <= 8'h10 ;
			data[23098] <= 8'h10 ;
			data[23099] <= 8'h10 ;
			data[23100] <= 8'h10 ;
			data[23101] <= 8'h10 ;
			data[23102] <= 8'h10 ;
			data[23103] <= 8'h10 ;
			data[23104] <= 8'h10 ;
			data[23105] <= 8'h10 ;
			data[23106] <= 8'h10 ;
			data[23107] <= 8'h10 ;
			data[23108] <= 8'h10 ;
			data[23109] <= 8'h10 ;
			data[23110] <= 8'h10 ;
			data[23111] <= 8'h10 ;
			data[23112] <= 8'h10 ;
			data[23113] <= 8'h10 ;
			data[23114] <= 8'h10 ;
			data[23115] <= 8'h10 ;
			data[23116] <= 8'h10 ;
			data[23117] <= 8'h10 ;
			data[23118] <= 8'h10 ;
			data[23119] <= 8'h10 ;
			data[23120] <= 8'h10 ;
			data[23121] <= 8'h10 ;
			data[23122] <= 8'h10 ;
			data[23123] <= 8'h10 ;
			data[23124] <= 8'h10 ;
			data[23125] <= 8'h10 ;
			data[23126] <= 8'h10 ;
			data[23127] <= 8'h10 ;
			data[23128] <= 8'h10 ;
			data[23129] <= 8'h10 ;
			data[23130] <= 8'h10 ;
			data[23131] <= 8'h10 ;
			data[23132] <= 8'h10 ;
			data[23133] <= 8'h10 ;
			data[23134] <= 8'h10 ;
			data[23135] <= 8'h10 ;
			data[23136] <= 8'h10 ;
			data[23137] <= 8'h10 ;
			data[23138] <= 8'h10 ;
			data[23139] <= 8'h10 ;
			data[23140] <= 8'h10 ;
			data[23141] <= 8'h10 ;
			data[23142] <= 8'h10 ;
			data[23143] <= 8'h10 ;
			data[23144] <= 8'h10 ;
			data[23145] <= 8'h10 ;
			data[23146] <= 8'h10 ;
			data[23147] <= 8'h10 ;
			data[23148] <= 8'h10 ;
			data[23149] <= 8'h10 ;
			data[23150] <= 8'h10 ;
			data[23151] <= 8'h10 ;
			data[23152] <= 8'h10 ;
			data[23153] <= 8'h10 ;
			data[23154] <= 8'h10 ;
			data[23155] <= 8'h10 ;
			data[23156] <= 8'h10 ;
			data[23157] <= 8'h10 ;
			data[23158] <= 8'h10 ;
			data[23159] <= 8'h10 ;
			data[23160] <= 8'h10 ;
			data[23161] <= 8'h10 ;
			data[23162] <= 8'h10 ;
			data[23163] <= 8'h10 ;
			data[23164] <= 8'h10 ;
			data[23165] <= 8'h10 ;
			data[23166] <= 8'h10 ;
			data[23167] <= 8'h10 ;
			data[23168] <= 8'h10 ;
			data[23169] <= 8'h10 ;
			data[23170] <= 8'h10 ;
			data[23171] <= 8'h10 ;
			data[23172] <= 8'h10 ;
			data[23173] <= 8'h10 ;
			data[23174] <= 8'h10 ;
			data[23175] <= 8'h10 ;
			data[23176] <= 8'h10 ;
			data[23177] <= 8'h10 ;
			data[23178] <= 8'h10 ;
			data[23179] <= 8'h10 ;
			data[23180] <= 8'h10 ;
			data[23181] <= 8'h10 ;
			data[23182] <= 8'h10 ;
			data[23183] <= 8'h10 ;
			data[23184] <= 8'h10 ;
			data[23185] <= 8'h10 ;
			data[23186] <= 8'h10 ;
			data[23187] <= 8'h10 ;
			data[23188] <= 8'h10 ;
			data[23189] <= 8'h10 ;
			data[23190] <= 8'h10 ;
			data[23191] <= 8'h10 ;
			data[23192] <= 8'h10 ;
			data[23193] <= 8'h10 ;
			data[23194] <= 8'h10 ;
			data[23195] <= 8'h10 ;
			data[23196] <= 8'h10 ;
			data[23197] <= 8'h10 ;
			data[23198] <= 8'h10 ;
			data[23199] <= 8'h10 ;
			data[23200] <= 8'h10 ;
			data[23201] <= 8'h10 ;
			data[23202] <= 8'h10 ;
			data[23203] <= 8'h10 ;
			data[23204] <= 8'h10 ;
			data[23205] <= 8'h10 ;
			data[23206] <= 8'h10 ;
			data[23207] <= 8'h10 ;
			data[23208] <= 8'h10 ;
			data[23209] <= 8'h10 ;
			data[23210] <= 8'h10 ;
			data[23211] <= 8'h10 ;
			data[23212] <= 8'h10 ;
			data[23213] <= 8'h10 ;
			data[23214] <= 8'h10 ;
			data[23215] <= 8'h10 ;
			data[23216] <= 8'h10 ;
			data[23217] <= 8'h10 ;
			data[23218] <= 8'h10 ;
			data[23219] <= 8'h10 ;
			data[23220] <= 8'h10 ;
			data[23221] <= 8'h10 ;
			data[23222] <= 8'h10 ;
			data[23223] <= 8'h10 ;
			data[23224] <= 8'h10 ;
			data[23225] <= 8'h10 ;
			data[23226] <= 8'h10 ;
			data[23227] <= 8'h10 ;
			data[23228] <= 8'h10 ;
			data[23229] <= 8'h10 ;
			data[23230] <= 8'h10 ;
			data[23231] <= 8'h10 ;
			data[23232] <= 8'h10 ;
			data[23233] <= 8'h10 ;
			data[23234] <= 8'h10 ;
			data[23235] <= 8'h10 ;
			data[23236] <= 8'h10 ;
			data[23237] <= 8'h10 ;
			data[23238] <= 8'h10 ;
			data[23239] <= 8'h10 ;
			data[23240] <= 8'h10 ;
			data[23241] <= 8'h10 ;
			data[23242] <= 8'h10 ;
			data[23243] <= 8'h10 ;
			data[23244] <= 8'h10 ;
			data[23245] <= 8'h10 ;
			data[23246] <= 8'h10 ;
			data[23247] <= 8'h10 ;
			data[23248] <= 8'h10 ;
			data[23249] <= 8'h10 ;
			data[23250] <= 8'h10 ;
			data[23251] <= 8'h10 ;
			data[23252] <= 8'h10 ;
			data[23253] <= 8'h10 ;
			data[23254] <= 8'h10 ;
			data[23255] <= 8'h10 ;
			data[23256] <= 8'h10 ;
			data[23257] <= 8'h10 ;
			data[23258] <= 8'h10 ;
			data[23259] <= 8'h10 ;
			data[23260] <= 8'h10 ;
			data[23261] <= 8'h10 ;
			data[23262] <= 8'h10 ;
			data[23263] <= 8'h10 ;
			data[23264] <= 8'h10 ;
			data[23265] <= 8'h10 ;
			data[23266] <= 8'h10 ;
			data[23267] <= 8'h10 ;
			data[23268] <= 8'h10 ;
			data[23269] <= 8'h10 ;
			data[23270] <= 8'h10 ;
			data[23271] <= 8'h10 ;
			data[23272] <= 8'h10 ;
			data[23273] <= 8'h10 ;
			data[23274] <= 8'h10 ;
			data[23275] <= 8'h10 ;
			data[23276] <= 8'h10 ;
			data[23277] <= 8'h10 ;
			data[23278] <= 8'h10 ;
			data[23279] <= 8'h10 ;
			data[23280] <= 8'h10 ;
			data[23281] <= 8'h10 ;
			data[23282] <= 8'h10 ;
			data[23283] <= 8'h10 ;
			data[23284] <= 8'h10 ;
			data[23285] <= 8'h10 ;
			data[23286] <= 8'h10 ;
			data[23287] <= 8'h10 ;
			data[23288] <= 8'h10 ;
			data[23289] <= 8'h10 ;
			data[23290] <= 8'h10 ;
			data[23291] <= 8'h10 ;
			data[23292] <= 8'h10 ;
			data[23293] <= 8'h10 ;
			data[23294] <= 8'h10 ;
			data[23295] <= 8'h10 ;
			data[23296] <= 8'h10 ;
			data[23297] <= 8'h10 ;
			data[23298] <= 8'h10 ;
			data[23299] <= 8'h10 ;
			data[23300] <= 8'h10 ;
			data[23301] <= 8'h10 ;
			data[23302] <= 8'h10 ;
			data[23303] <= 8'h10 ;
			data[23304] <= 8'h10 ;
			data[23305] <= 8'h10 ;
			data[23306] <= 8'h10 ;
			data[23307] <= 8'h10 ;
			data[23308] <= 8'h10 ;
			data[23309] <= 8'h10 ;
			data[23310] <= 8'h10 ;
			data[23311] <= 8'h10 ;
			data[23312] <= 8'h10 ;
			data[23313] <= 8'h10 ;
			data[23314] <= 8'h10 ;
			data[23315] <= 8'h10 ;
			data[23316] <= 8'h10 ;
			data[23317] <= 8'h10 ;
			data[23318] <= 8'h10 ;
			data[23319] <= 8'h10 ;
			data[23320] <= 8'h10 ;
			data[23321] <= 8'h10 ;
			data[23322] <= 8'h10 ;
			data[23323] <= 8'h10 ;
			data[23324] <= 8'h10 ;
			data[23325] <= 8'h10 ;
			data[23326] <= 8'h10 ;
			data[23327] <= 8'h10 ;
			data[23328] <= 8'h10 ;
			data[23329] <= 8'h10 ;
			data[23330] <= 8'h10 ;
			data[23331] <= 8'h10 ;
			data[23332] <= 8'h10 ;
			data[23333] <= 8'h10 ;
			data[23334] <= 8'h10 ;
			data[23335] <= 8'h10 ;
			data[23336] <= 8'h10 ;
			data[23337] <= 8'h10 ;
			data[23338] <= 8'h10 ;
			data[23339] <= 8'h10 ;
			data[23340] <= 8'h10 ;
			data[23341] <= 8'h10 ;
			data[23342] <= 8'h10 ;
			data[23343] <= 8'h10 ;
			data[23344] <= 8'h10 ;
			data[23345] <= 8'h10 ;
			data[23346] <= 8'h10 ;
			data[23347] <= 8'h10 ;
			data[23348] <= 8'h10 ;
			data[23349] <= 8'h10 ;
			data[23350] <= 8'h10 ;
			data[23351] <= 8'h10 ;
			data[23352] <= 8'h10 ;
			data[23353] <= 8'h10 ;
			data[23354] <= 8'h10 ;
			data[23355] <= 8'h10 ;
			data[23356] <= 8'h10 ;
			data[23357] <= 8'h10 ;
			data[23358] <= 8'h10 ;
			data[23359] <= 8'h10 ;
			data[23360] <= 8'h10 ;
			data[23361] <= 8'h10 ;
			data[23362] <= 8'h10 ;
			data[23363] <= 8'h10 ;
			data[23364] <= 8'h10 ;
			data[23365] <= 8'h10 ;
			data[23366] <= 8'h10 ;
			data[23367] <= 8'h10 ;
			data[23368] <= 8'h10 ;
			data[23369] <= 8'h10 ;
			data[23370] <= 8'h10 ;
			data[23371] <= 8'h10 ;
			data[23372] <= 8'h10 ;
			data[23373] <= 8'h10 ;
			data[23374] <= 8'h10 ;
			data[23375] <= 8'h10 ;
			data[23376] <= 8'h10 ;
			data[23377] <= 8'h10 ;
			data[23378] <= 8'h10 ;
			data[23379] <= 8'h10 ;
			data[23380] <= 8'h10 ;
			data[23381] <= 8'h10 ;
			data[23382] <= 8'h10 ;
			data[23383] <= 8'h10 ;
			data[23384] <= 8'h10 ;
			data[23385] <= 8'h10 ;
			data[23386] <= 8'h10 ;
			data[23387] <= 8'h10 ;
			data[23388] <= 8'h10 ;
			data[23389] <= 8'h10 ;
			data[23390] <= 8'h10 ;
			data[23391] <= 8'h10 ;
			data[23392] <= 8'h10 ;
			data[23393] <= 8'h10 ;
			data[23394] <= 8'h10 ;
			data[23395] <= 8'h10 ;
			data[23396] <= 8'h10 ;
			data[23397] <= 8'h10 ;
			data[23398] <= 8'h10 ;
			data[23399] <= 8'h10 ;
			data[23400] <= 8'h10 ;
			data[23401] <= 8'h10 ;
			data[23402] <= 8'h10 ;
			data[23403] <= 8'h10 ;
			data[23404] <= 8'h10 ;
			data[23405] <= 8'h10 ;
			data[23406] <= 8'h10 ;
			data[23407] <= 8'h10 ;
			data[23408] <= 8'h10 ;
			data[23409] <= 8'h10 ;
			data[23410] <= 8'h10 ;
			data[23411] <= 8'h10 ;
			data[23412] <= 8'h10 ;
			data[23413] <= 8'h10 ;
			data[23414] <= 8'h10 ;
			data[23415] <= 8'h10 ;
			data[23416] <= 8'h10 ;
			data[23417] <= 8'h10 ;
			data[23418] <= 8'h10 ;
			data[23419] <= 8'h10 ;
			data[23420] <= 8'h10 ;
			data[23421] <= 8'h10 ;
			data[23422] <= 8'h10 ;
			data[23423] <= 8'h10 ;
			data[23424] <= 8'h10 ;
			data[23425] <= 8'h10 ;
			data[23426] <= 8'h10 ;
			data[23427] <= 8'h10 ;
			data[23428] <= 8'h10 ;
			data[23429] <= 8'h10 ;
			data[23430] <= 8'h10 ;
			data[23431] <= 8'h10 ;
			data[23432] <= 8'h10 ;
			data[23433] <= 8'h10 ;
			data[23434] <= 8'h10 ;
			data[23435] <= 8'h10 ;
			data[23436] <= 8'h10 ;
			data[23437] <= 8'h10 ;
			data[23438] <= 8'h10 ;
			data[23439] <= 8'h10 ;
			data[23440] <= 8'h10 ;
			data[23441] <= 8'h10 ;
			data[23442] <= 8'h10 ;
			data[23443] <= 8'h10 ;
			data[23444] <= 8'h10 ;
			data[23445] <= 8'h10 ;
			data[23446] <= 8'h10 ;
			data[23447] <= 8'h10 ;
			data[23448] <= 8'h10 ;
			data[23449] <= 8'h10 ;
			data[23450] <= 8'h10 ;
			data[23451] <= 8'h10 ;
			data[23452] <= 8'h10 ;
			data[23453] <= 8'h10 ;
			data[23454] <= 8'h10 ;
			data[23455] <= 8'h10 ;
			data[23456] <= 8'h10 ;
			data[23457] <= 8'h10 ;
			data[23458] <= 8'h10 ;
			data[23459] <= 8'h10 ;
			data[23460] <= 8'h10 ;
			data[23461] <= 8'h10 ;
			data[23462] <= 8'h10 ;
			data[23463] <= 8'h10 ;
			data[23464] <= 8'h10 ;
			data[23465] <= 8'h10 ;
			data[23466] <= 8'h10 ;
			data[23467] <= 8'h10 ;
			data[23468] <= 8'h10 ;
			data[23469] <= 8'h10 ;
			data[23470] <= 8'h10 ;
			data[23471] <= 8'h10 ;
			data[23472] <= 8'h10 ;
			data[23473] <= 8'h10 ;
			data[23474] <= 8'h10 ;
			data[23475] <= 8'h10 ;
			data[23476] <= 8'h10 ;
			data[23477] <= 8'h10 ;
			data[23478] <= 8'h10 ;
			data[23479] <= 8'h10 ;
			data[23480] <= 8'h10 ;
			data[23481] <= 8'h10 ;
			data[23482] <= 8'h10 ;
			data[23483] <= 8'h10 ;
			data[23484] <= 8'h10 ;
			data[23485] <= 8'h10 ;
			data[23486] <= 8'h10 ;
			data[23487] <= 8'h10 ;
			data[23488] <= 8'h10 ;
			data[23489] <= 8'h10 ;
			data[23490] <= 8'h10 ;
			data[23491] <= 8'h10 ;
			data[23492] <= 8'h10 ;
			data[23493] <= 8'h10 ;
			data[23494] <= 8'h10 ;
			data[23495] <= 8'h10 ;
			data[23496] <= 8'h10 ;
			data[23497] <= 8'h10 ;
			data[23498] <= 8'h10 ;
			data[23499] <= 8'h10 ;
			data[23500] <= 8'h10 ;
			data[23501] <= 8'h10 ;
			data[23502] <= 8'h10 ;
			data[23503] <= 8'h10 ;
			data[23504] <= 8'h10 ;
			data[23505] <= 8'h10 ;
			data[23506] <= 8'h10 ;
			data[23507] <= 8'h10 ;
			data[23508] <= 8'h10 ;
			data[23509] <= 8'h10 ;
			data[23510] <= 8'h10 ;
			data[23511] <= 8'h10 ;
			data[23512] <= 8'h10 ;
			data[23513] <= 8'h10 ;
			data[23514] <= 8'h10 ;
			data[23515] <= 8'h10 ;
			data[23516] <= 8'h10 ;
			data[23517] <= 8'h10 ;
			data[23518] <= 8'h10 ;
			data[23519] <= 8'h10 ;
			data[23520] <= 8'h10 ;
			data[23521] <= 8'h10 ;
			data[23522] <= 8'h10 ;
			data[23523] <= 8'h10 ;
			data[23524] <= 8'h10 ;
			data[23525] <= 8'h10 ;
			data[23526] <= 8'h10 ;
			data[23527] <= 8'h10 ;
			data[23528] <= 8'h10 ;
			data[23529] <= 8'h10 ;
			data[23530] <= 8'h10 ;
			data[23531] <= 8'h10 ;
			data[23532] <= 8'h10 ;
			data[23533] <= 8'h10 ;
			data[23534] <= 8'h10 ;
			data[23535] <= 8'h10 ;
			data[23536] <= 8'h10 ;
			data[23537] <= 8'h10 ;
			data[23538] <= 8'h10 ;
			data[23539] <= 8'h10 ;
			data[23540] <= 8'h10 ;
			data[23541] <= 8'h10 ;
			data[23542] <= 8'h10 ;
			data[23543] <= 8'h10 ;
			data[23544] <= 8'h10 ;
			data[23545] <= 8'h10 ;
			data[23546] <= 8'h10 ;
			data[23547] <= 8'h10 ;
			data[23548] <= 8'h10 ;
			data[23549] <= 8'h10 ;
			data[23550] <= 8'h10 ;
			data[23551] <= 8'h10 ;
			data[23552] <= 8'h10 ;
			data[23553] <= 8'h10 ;
			data[23554] <= 8'h10 ;
			data[23555] <= 8'h10 ;
			data[23556] <= 8'h10 ;
			data[23557] <= 8'h10 ;
			data[23558] <= 8'h10 ;
			data[23559] <= 8'h10 ;
			data[23560] <= 8'h10 ;
			data[23561] <= 8'h10 ;
			data[23562] <= 8'h10 ;
			data[23563] <= 8'h10 ;
			data[23564] <= 8'h10 ;
			data[23565] <= 8'h10 ;
			data[23566] <= 8'h10 ;
			data[23567] <= 8'h10 ;
			data[23568] <= 8'h10 ;
			data[23569] <= 8'h10 ;
			data[23570] <= 8'h10 ;
			data[23571] <= 8'h10 ;
			data[23572] <= 8'h10 ;
			data[23573] <= 8'h10 ;
			data[23574] <= 8'h10 ;
			data[23575] <= 8'h10 ;
			data[23576] <= 8'h10 ;
			data[23577] <= 8'h10 ;
			data[23578] <= 8'h10 ;
			data[23579] <= 8'h10 ;
			data[23580] <= 8'h10 ;
			data[23581] <= 8'h10 ;
			data[23582] <= 8'h10 ;
			data[23583] <= 8'h10 ;
			data[23584] <= 8'h10 ;
			data[23585] <= 8'h10 ;
			data[23586] <= 8'h10 ;
			data[23587] <= 8'h10 ;
			data[23588] <= 8'h10 ;
			data[23589] <= 8'h10 ;
			data[23590] <= 8'h10 ;
			data[23591] <= 8'h10 ;
			data[23592] <= 8'h10 ;
			data[23593] <= 8'h10 ;
			data[23594] <= 8'h10 ;
			data[23595] <= 8'h10 ;
			data[23596] <= 8'h10 ;
			data[23597] <= 8'h10 ;
			data[23598] <= 8'h10 ;
			data[23599] <= 8'h10 ;
			data[23600] <= 8'h10 ;
			data[23601] <= 8'h10 ;
			data[23602] <= 8'h10 ;
			data[23603] <= 8'h10 ;
			data[23604] <= 8'h10 ;
			data[23605] <= 8'h10 ;
			data[23606] <= 8'h10 ;
			data[23607] <= 8'h10 ;
			data[23608] <= 8'h10 ;
			data[23609] <= 8'h10 ;
			data[23610] <= 8'h10 ;
			data[23611] <= 8'h10 ;
			data[23612] <= 8'h10 ;
			data[23613] <= 8'h10 ;
			data[23614] <= 8'h10 ;
			data[23615] <= 8'h10 ;
			data[23616] <= 8'h10 ;
			data[23617] <= 8'h10 ;
			data[23618] <= 8'h10 ;
			data[23619] <= 8'h10 ;
			data[23620] <= 8'h10 ;
			data[23621] <= 8'h10 ;
			data[23622] <= 8'h10 ;
			data[23623] <= 8'h10 ;
			data[23624] <= 8'h10 ;
			data[23625] <= 8'h10 ;
			data[23626] <= 8'h10 ;
			data[23627] <= 8'h10 ;
			data[23628] <= 8'h10 ;
			data[23629] <= 8'h10 ;
			data[23630] <= 8'h10 ;
			data[23631] <= 8'h10 ;
			data[23632] <= 8'h10 ;
			data[23633] <= 8'h10 ;
			data[23634] <= 8'h10 ;
			data[23635] <= 8'h10 ;
			data[23636] <= 8'h10 ;
			data[23637] <= 8'h10 ;
			data[23638] <= 8'h10 ;
			data[23639] <= 8'h10 ;
			data[23640] <= 8'h10 ;
			data[23641] <= 8'h10 ;
			data[23642] <= 8'h10 ;
			data[23643] <= 8'h10 ;
			data[23644] <= 8'h10 ;
			data[23645] <= 8'h10 ;
			data[23646] <= 8'h10 ;
			data[23647] <= 8'h10 ;
			data[23648] <= 8'h10 ;
			data[23649] <= 8'h10 ;
			data[23650] <= 8'h10 ;
			data[23651] <= 8'h10 ;
			data[23652] <= 8'h10 ;
			data[23653] <= 8'h10 ;
			data[23654] <= 8'h10 ;
			data[23655] <= 8'h10 ;
			data[23656] <= 8'h10 ;
			data[23657] <= 8'h10 ;
			data[23658] <= 8'h10 ;
			data[23659] <= 8'h10 ;
			data[23660] <= 8'h10 ;
			data[23661] <= 8'h10 ;
			data[23662] <= 8'h10 ;
			data[23663] <= 8'h10 ;
			data[23664] <= 8'h10 ;
			data[23665] <= 8'h10 ;
			data[23666] <= 8'h10 ;
			data[23667] <= 8'h10 ;
			data[23668] <= 8'h10 ;
			data[23669] <= 8'h10 ;
			data[23670] <= 8'h10 ;
			data[23671] <= 8'h10 ;
			data[23672] <= 8'h10 ;
			data[23673] <= 8'h10 ;
			data[23674] <= 8'h10 ;
			data[23675] <= 8'h10 ;
			data[23676] <= 8'h10 ;
			data[23677] <= 8'h10 ;
			data[23678] <= 8'h10 ;
			data[23679] <= 8'h10 ;
			data[23680] <= 8'h10 ;
			data[23681] <= 8'h10 ;
			data[23682] <= 8'h10 ;
			data[23683] <= 8'h10 ;
			data[23684] <= 8'h10 ;
			data[23685] <= 8'h10 ;
			data[23686] <= 8'h10 ;
			data[23687] <= 8'h10 ;
			data[23688] <= 8'h10 ;
			data[23689] <= 8'h10 ;
			data[23690] <= 8'h10 ;
			data[23691] <= 8'h10 ;
			data[23692] <= 8'h10 ;
			data[23693] <= 8'h10 ;
			data[23694] <= 8'h10 ;
			data[23695] <= 8'h10 ;
			data[23696] <= 8'h10 ;
			data[23697] <= 8'h10 ;
			data[23698] <= 8'h10 ;
			data[23699] <= 8'h10 ;
			data[23700] <= 8'h10 ;
			data[23701] <= 8'h10 ;
			data[23702] <= 8'h10 ;
			data[23703] <= 8'h10 ;
			data[23704] <= 8'h10 ;
			data[23705] <= 8'h10 ;
			data[23706] <= 8'h10 ;
			data[23707] <= 8'h10 ;
			data[23708] <= 8'h10 ;
			data[23709] <= 8'h10 ;
			data[23710] <= 8'h10 ;
			data[23711] <= 8'h10 ;
			data[23712] <= 8'h10 ;
			data[23713] <= 8'h10 ;
			data[23714] <= 8'h10 ;
			data[23715] <= 8'h10 ;
			data[23716] <= 8'h10 ;
			data[23717] <= 8'h10 ;
			data[23718] <= 8'h10 ;
			data[23719] <= 8'h10 ;
			data[23720] <= 8'h10 ;
			data[23721] <= 8'h10 ;
			data[23722] <= 8'h10 ;
			data[23723] <= 8'h10 ;
			data[23724] <= 8'h10 ;
			data[23725] <= 8'h10 ;
			data[23726] <= 8'h10 ;
			data[23727] <= 8'h10 ;
			data[23728] <= 8'h10 ;
			data[23729] <= 8'h10 ;
			data[23730] <= 8'h10 ;
			data[23731] <= 8'h10 ;
			data[23732] <= 8'h10 ;
			data[23733] <= 8'h10 ;
			data[23734] <= 8'h10 ;
			data[23735] <= 8'h10 ;
			data[23736] <= 8'h10 ;
			data[23737] <= 8'h10 ;
			data[23738] <= 8'h10 ;
			data[23739] <= 8'h10 ;
			data[23740] <= 8'h10 ;
			data[23741] <= 8'h10 ;
			data[23742] <= 8'h10 ;
			data[23743] <= 8'h10 ;
			data[23744] <= 8'h10 ;
			data[23745] <= 8'h10 ;
			data[23746] <= 8'h10 ;
			data[23747] <= 8'h10 ;
			data[23748] <= 8'h10 ;
			data[23749] <= 8'h10 ;
			data[23750] <= 8'h10 ;
			data[23751] <= 8'h10 ;
			data[23752] <= 8'h10 ;
			data[23753] <= 8'h10 ;
			data[23754] <= 8'h10 ;
			data[23755] <= 8'h10 ;
			data[23756] <= 8'h10 ;
			data[23757] <= 8'h10 ;
			data[23758] <= 8'h10 ;
			data[23759] <= 8'h10 ;
			data[23760] <= 8'h10 ;
			data[23761] <= 8'h10 ;
			data[23762] <= 8'h10 ;
			data[23763] <= 8'h10 ;
			data[23764] <= 8'h10 ;
			data[23765] <= 8'h10 ;
			data[23766] <= 8'h10 ;
			data[23767] <= 8'h10 ;
			data[23768] <= 8'h10 ;
			data[23769] <= 8'h10 ;
			data[23770] <= 8'h10 ;
			data[23771] <= 8'h10 ;
			data[23772] <= 8'h10 ;
			data[23773] <= 8'h10 ;
			data[23774] <= 8'h10 ;
			data[23775] <= 8'h10 ;
			data[23776] <= 8'h10 ;
			data[23777] <= 8'h10 ;
			data[23778] <= 8'h10 ;
			data[23779] <= 8'h10 ;
			data[23780] <= 8'h10 ;
			data[23781] <= 8'h10 ;
			data[23782] <= 8'h10 ;
			data[23783] <= 8'h10 ;
			data[23784] <= 8'h10 ;
			data[23785] <= 8'h10 ;
			data[23786] <= 8'h10 ;
			data[23787] <= 8'h10 ;
			data[23788] <= 8'h10 ;
			data[23789] <= 8'h10 ;
			data[23790] <= 8'h10 ;
			data[23791] <= 8'h10 ;
			data[23792] <= 8'h10 ;
			data[23793] <= 8'h10 ;
			data[23794] <= 8'h10 ;
			data[23795] <= 8'h10 ;
			data[23796] <= 8'h10 ;
			data[23797] <= 8'h10 ;
			data[23798] <= 8'h10 ;
			data[23799] <= 8'h10 ;
			data[23800] <= 8'h10 ;
			data[23801] <= 8'h10 ;
			data[23802] <= 8'h10 ;
			data[23803] <= 8'h10 ;
			data[23804] <= 8'h10 ;
			data[23805] <= 8'h10 ;
			data[23806] <= 8'h10 ;
			data[23807] <= 8'h10 ;
			data[23808] <= 8'h10 ;
			data[23809] <= 8'h10 ;
			data[23810] <= 8'h10 ;
			data[23811] <= 8'h10 ;
			data[23812] <= 8'h10 ;
			data[23813] <= 8'h10 ;
			data[23814] <= 8'h10 ;
			data[23815] <= 8'h10 ;
			data[23816] <= 8'h10 ;
			data[23817] <= 8'h10 ;
			data[23818] <= 8'h10 ;
			data[23819] <= 8'h10 ;
			data[23820] <= 8'h10 ;
			data[23821] <= 8'h10 ;
			data[23822] <= 8'h10 ;
			data[23823] <= 8'h10 ;
			data[23824] <= 8'h10 ;
			data[23825] <= 8'h10 ;
			data[23826] <= 8'h10 ;
			data[23827] <= 8'h10 ;
			data[23828] <= 8'h10 ;
			data[23829] <= 8'h10 ;
			data[23830] <= 8'h10 ;
			data[23831] <= 8'h10 ;
			data[23832] <= 8'h10 ;
			data[23833] <= 8'h10 ;
			data[23834] <= 8'h10 ;
			data[23835] <= 8'h10 ;
			data[23836] <= 8'h10 ;
			data[23837] <= 8'h10 ;
			data[23838] <= 8'h10 ;
			data[23839] <= 8'h10 ;
			data[23840] <= 8'h10 ;
			data[23841] <= 8'h10 ;
			data[23842] <= 8'h10 ;
			data[23843] <= 8'h10 ;
			data[23844] <= 8'h10 ;
			data[23845] <= 8'h10 ;
			data[23846] <= 8'h10 ;
			data[23847] <= 8'h10 ;
			data[23848] <= 8'h10 ;
			data[23849] <= 8'h10 ;
			data[23850] <= 8'h10 ;
			data[23851] <= 8'h10 ;
			data[23852] <= 8'h10 ;
			data[23853] <= 8'h10 ;
			data[23854] <= 8'h10 ;
			data[23855] <= 8'h10 ;
			data[23856] <= 8'h10 ;
			data[23857] <= 8'h10 ;
			data[23858] <= 8'h10 ;
			data[23859] <= 8'h10 ;
			data[23860] <= 8'h10 ;
			data[23861] <= 8'h10 ;
			data[23862] <= 8'h10 ;
			data[23863] <= 8'h10 ;
			data[23864] <= 8'h10 ;
			data[23865] <= 8'h10 ;
			data[23866] <= 8'h10 ;
			data[23867] <= 8'h10 ;
			data[23868] <= 8'h10 ;
			data[23869] <= 8'h10 ;
			data[23870] <= 8'h10 ;
			data[23871] <= 8'h10 ;
			data[23872] <= 8'h10 ;
			data[23873] <= 8'h10 ;
			data[23874] <= 8'h10 ;
			data[23875] <= 8'h10 ;
			data[23876] <= 8'h10 ;
			data[23877] <= 8'h10 ;
			data[23878] <= 8'h10 ;
			data[23879] <= 8'h10 ;
			data[23880] <= 8'h10 ;
			data[23881] <= 8'h10 ;
			data[23882] <= 8'h10 ;
			data[23883] <= 8'h10 ;
			data[23884] <= 8'h10 ;
			data[23885] <= 8'h10 ;
			data[23886] <= 8'h10 ;
			data[23887] <= 8'h10 ;
			data[23888] <= 8'h10 ;
			data[23889] <= 8'h10 ;
			data[23890] <= 8'h10 ;
			data[23891] <= 8'h10 ;
			data[23892] <= 8'h10 ;
			data[23893] <= 8'h10 ;
			data[23894] <= 8'h10 ;
			data[23895] <= 8'h10 ;
			data[23896] <= 8'h10 ;
			data[23897] <= 8'h10 ;
			data[23898] <= 8'h10 ;
			data[23899] <= 8'h10 ;
			data[23900] <= 8'h10 ;
			data[23901] <= 8'h10 ;
			data[23902] <= 8'h10 ;
			data[23903] <= 8'h10 ;
			data[23904] <= 8'h10 ;
			data[23905] <= 8'h10 ;
			data[23906] <= 8'h10 ;
			data[23907] <= 8'h10 ;
			data[23908] <= 8'h10 ;
			data[23909] <= 8'h10 ;
			data[23910] <= 8'h10 ;
			data[23911] <= 8'h10 ;
			data[23912] <= 8'h10 ;
			data[23913] <= 8'h10 ;
			data[23914] <= 8'h10 ;
			data[23915] <= 8'h10 ;
			data[23916] <= 8'h10 ;
			data[23917] <= 8'h10 ;
			data[23918] <= 8'h10 ;
			data[23919] <= 8'h10 ;
			data[23920] <= 8'h10 ;
			data[23921] <= 8'h10 ;
			data[23922] <= 8'h10 ;
			data[23923] <= 8'h10 ;
			data[23924] <= 8'h10 ;
			data[23925] <= 8'h10 ;
			data[23926] <= 8'h10 ;
			data[23927] <= 8'h10 ;
			data[23928] <= 8'h10 ;
			data[23929] <= 8'h10 ;
			data[23930] <= 8'h10 ;
			data[23931] <= 8'h10 ;
			data[23932] <= 8'h10 ;
			data[23933] <= 8'h10 ;
			data[23934] <= 8'h10 ;
			data[23935] <= 8'h10 ;
			data[23936] <= 8'h10 ;
			data[23937] <= 8'h10 ;
			data[23938] <= 8'h10 ;
			data[23939] <= 8'h10 ;
			data[23940] <= 8'h10 ;
			data[23941] <= 8'h10 ;
			data[23942] <= 8'h10 ;
			data[23943] <= 8'h10 ;
			data[23944] <= 8'h10 ;
			data[23945] <= 8'h10 ;
			data[23946] <= 8'h10 ;
			data[23947] <= 8'h10 ;
			data[23948] <= 8'h10 ;
			data[23949] <= 8'h10 ;
			data[23950] <= 8'h10 ;
			data[23951] <= 8'h10 ;
			data[23952] <= 8'h10 ;
			data[23953] <= 8'h10 ;
			data[23954] <= 8'h10 ;
			data[23955] <= 8'h10 ;
			data[23956] <= 8'h10 ;
			data[23957] <= 8'h10 ;
			data[23958] <= 8'h10 ;
			data[23959] <= 8'h10 ;
			data[23960] <= 8'h10 ;
			data[23961] <= 8'h10 ;
			data[23962] <= 8'h10 ;
			data[23963] <= 8'h10 ;
			data[23964] <= 8'h10 ;
			data[23965] <= 8'h10 ;
			data[23966] <= 8'h10 ;
			data[23967] <= 8'h10 ;
			data[23968] <= 8'h10 ;
			data[23969] <= 8'h10 ;
			data[23970] <= 8'h10 ;
			data[23971] <= 8'h10 ;
			data[23972] <= 8'h10 ;
			data[23973] <= 8'h10 ;
			data[23974] <= 8'h10 ;
			data[23975] <= 8'h10 ;
			data[23976] <= 8'h10 ;
			data[23977] <= 8'h10 ;
			data[23978] <= 8'h10 ;
			data[23979] <= 8'h10 ;
			data[23980] <= 8'h10 ;
			data[23981] <= 8'h10 ;
			data[23982] <= 8'h10 ;
			data[23983] <= 8'h10 ;
			data[23984] <= 8'h10 ;
			data[23985] <= 8'h10 ;
			data[23986] <= 8'h10 ;
			data[23987] <= 8'h10 ;
			data[23988] <= 8'h10 ;
			data[23989] <= 8'h10 ;
			data[23990] <= 8'h10 ;
			data[23991] <= 8'h10 ;
			data[23992] <= 8'h10 ;
			data[23993] <= 8'h10 ;
			data[23994] <= 8'h10 ;
			data[23995] <= 8'h10 ;
			data[23996] <= 8'h10 ;
			data[23997] <= 8'h10 ;
			data[23998] <= 8'h10 ;
			data[23999] <= 8'h10 ;
			data[24000] <= 8'h10 ;
			data[24001] <= 8'h10 ;
			data[24002] <= 8'h10 ;
			data[24003] <= 8'h10 ;
			data[24004] <= 8'h10 ;
			data[24005] <= 8'h10 ;
			data[24006] <= 8'h10 ;
			data[24007] <= 8'h10 ;
			data[24008] <= 8'h10 ;
			data[24009] <= 8'h10 ;
			data[24010] <= 8'h10 ;
			data[24011] <= 8'h10 ;
			data[24012] <= 8'h10 ;
			data[24013] <= 8'h10 ;
			data[24014] <= 8'h10 ;
			data[24015] <= 8'h10 ;
			data[24016] <= 8'h10 ;
			data[24017] <= 8'h10 ;
			data[24018] <= 8'h10 ;
			data[24019] <= 8'h10 ;
			data[24020] <= 8'h10 ;
			data[24021] <= 8'h10 ;
			data[24022] <= 8'h10 ;
			data[24023] <= 8'h10 ;
			data[24024] <= 8'h10 ;
			data[24025] <= 8'h10 ;
			data[24026] <= 8'h10 ;
			data[24027] <= 8'h10 ;
			data[24028] <= 8'h10 ;
			data[24029] <= 8'h10 ;
			data[24030] <= 8'h10 ;
			data[24031] <= 8'h10 ;
			data[24032] <= 8'h10 ;
			data[24033] <= 8'h10 ;
			data[24034] <= 8'h10 ;
			data[24035] <= 8'h10 ;
			data[24036] <= 8'h10 ;
			data[24037] <= 8'h10 ;
			data[24038] <= 8'h10 ;
			data[24039] <= 8'h10 ;
			data[24040] <= 8'h10 ;
			data[24041] <= 8'h10 ;
			data[24042] <= 8'h10 ;
			data[24043] <= 8'h10 ;
			data[24044] <= 8'h10 ;
			data[24045] <= 8'h10 ;
			data[24046] <= 8'h10 ;
			data[24047] <= 8'h10 ;
			data[24048] <= 8'h10 ;
			data[24049] <= 8'h10 ;
			data[24050] <= 8'h10 ;
			data[24051] <= 8'h10 ;
			data[24052] <= 8'h10 ;
			data[24053] <= 8'h10 ;
			data[24054] <= 8'h10 ;
			data[24055] <= 8'h10 ;
			data[24056] <= 8'h10 ;
			data[24057] <= 8'h10 ;
			data[24058] <= 8'h10 ;
			data[24059] <= 8'h10 ;
			data[24060] <= 8'h10 ;
			data[24061] <= 8'h10 ;
			data[24062] <= 8'h10 ;
			data[24063] <= 8'h10 ;
			data[24064] <= 8'h10 ;
			data[24065] <= 8'h10 ;
			data[24066] <= 8'h10 ;
			data[24067] <= 8'h10 ;
			data[24068] <= 8'h10 ;
			data[24069] <= 8'h10 ;
			data[24070] <= 8'h10 ;
			data[24071] <= 8'h10 ;
			data[24072] <= 8'h10 ;
			data[24073] <= 8'h10 ;
			data[24074] <= 8'h10 ;
			data[24075] <= 8'h10 ;
			data[24076] <= 8'h10 ;
			data[24077] <= 8'h10 ;
			data[24078] <= 8'h10 ;
			data[24079] <= 8'h10 ;
			data[24080] <= 8'h10 ;
			data[24081] <= 8'h10 ;
			data[24082] <= 8'h10 ;
			data[24083] <= 8'h10 ;
			data[24084] <= 8'h10 ;
			data[24085] <= 8'h10 ;
			data[24086] <= 8'h10 ;
			data[24087] <= 8'h10 ;
			data[24088] <= 8'h10 ;
			data[24089] <= 8'h10 ;
			data[24090] <= 8'h10 ;
			data[24091] <= 8'h10 ;
			data[24092] <= 8'h10 ;
			data[24093] <= 8'h10 ;
			data[24094] <= 8'h10 ;
			data[24095] <= 8'h10 ;
			data[24096] <= 8'h10 ;
			data[24097] <= 8'h10 ;
			data[24098] <= 8'h10 ;
			data[24099] <= 8'h10 ;
			data[24100] <= 8'h10 ;
			data[24101] <= 8'h10 ;
			data[24102] <= 8'h10 ;
			data[24103] <= 8'h10 ;
			data[24104] <= 8'h10 ;
			data[24105] <= 8'h10 ;
			data[24106] <= 8'h10 ;
			data[24107] <= 8'h10 ;
			data[24108] <= 8'h10 ;
			data[24109] <= 8'h10 ;
			data[24110] <= 8'h10 ;
			data[24111] <= 8'h10 ;
			data[24112] <= 8'h10 ;
			data[24113] <= 8'h10 ;
			data[24114] <= 8'h10 ;
			data[24115] <= 8'h10 ;
			data[24116] <= 8'h10 ;
			data[24117] <= 8'h10 ;
			data[24118] <= 8'h10 ;
			data[24119] <= 8'h10 ;
			data[24120] <= 8'h10 ;
			data[24121] <= 8'h10 ;
			data[24122] <= 8'h10 ;
			data[24123] <= 8'h10 ;
			data[24124] <= 8'h10 ;
			data[24125] <= 8'h10 ;
			data[24126] <= 8'h10 ;
			data[24127] <= 8'h10 ;
			data[24128] <= 8'h10 ;
			data[24129] <= 8'h10 ;
			data[24130] <= 8'h10 ;
			data[24131] <= 8'h10 ;
			data[24132] <= 8'h10 ;
			data[24133] <= 8'h10 ;
			data[24134] <= 8'h10 ;
			data[24135] <= 8'h10 ;
			data[24136] <= 8'h10 ;
			data[24137] <= 8'h10 ;
			data[24138] <= 8'h10 ;
			data[24139] <= 8'h10 ;
			data[24140] <= 8'h10 ;
			data[24141] <= 8'h10 ;
			data[24142] <= 8'h10 ;
			data[24143] <= 8'h10 ;
			data[24144] <= 8'h10 ;
			data[24145] <= 8'h10 ;
			data[24146] <= 8'h10 ;
			data[24147] <= 8'h10 ;
			data[24148] <= 8'h10 ;
			data[24149] <= 8'h10 ;
			data[24150] <= 8'h10 ;
			data[24151] <= 8'h10 ;
			data[24152] <= 8'h10 ;
			data[24153] <= 8'h10 ;
			data[24154] <= 8'h10 ;
			data[24155] <= 8'h10 ;
			data[24156] <= 8'h10 ;
			data[24157] <= 8'h10 ;
			data[24158] <= 8'h10 ;
			data[24159] <= 8'h10 ;
			data[24160] <= 8'h10 ;
			data[24161] <= 8'h10 ;
			data[24162] <= 8'h10 ;
			data[24163] <= 8'h10 ;
			data[24164] <= 8'h10 ;
			data[24165] <= 8'h10 ;
			data[24166] <= 8'h10 ;
			data[24167] <= 8'h10 ;
			data[24168] <= 8'h10 ;
			data[24169] <= 8'h10 ;
			data[24170] <= 8'h10 ;
			data[24171] <= 8'h10 ;
			data[24172] <= 8'h10 ;
			data[24173] <= 8'h10 ;
			data[24174] <= 8'h10 ;
			data[24175] <= 8'h10 ;
			data[24176] <= 8'h10 ;
			data[24177] <= 8'h10 ;
			data[24178] <= 8'h10 ;
			data[24179] <= 8'h10 ;
			data[24180] <= 8'h10 ;
			data[24181] <= 8'h10 ;
			data[24182] <= 8'h10 ;
			data[24183] <= 8'h10 ;
			data[24184] <= 8'h10 ;
			data[24185] <= 8'h10 ;
			data[24186] <= 8'h10 ;
			data[24187] <= 8'h10 ;
			data[24188] <= 8'h10 ;
			data[24189] <= 8'h10 ;
			data[24190] <= 8'h10 ;
			data[24191] <= 8'h10 ;
			data[24192] <= 8'h10 ;
			data[24193] <= 8'h10 ;
			data[24194] <= 8'h10 ;
			data[24195] <= 8'h10 ;
			data[24196] <= 8'h10 ;
			data[24197] <= 8'h10 ;
			data[24198] <= 8'h10 ;
			data[24199] <= 8'h10 ;
			data[24200] <= 8'h10 ;
			data[24201] <= 8'h10 ;
			data[24202] <= 8'h10 ;
			data[24203] <= 8'h10 ;
			data[24204] <= 8'h10 ;
			data[24205] <= 8'h10 ;
			data[24206] <= 8'h10 ;
			data[24207] <= 8'h10 ;
			data[24208] <= 8'h10 ;
			data[24209] <= 8'h10 ;
			data[24210] <= 8'h10 ;
			data[24211] <= 8'h10 ;
			data[24212] <= 8'h10 ;
			data[24213] <= 8'h10 ;
			data[24214] <= 8'h10 ;
			data[24215] <= 8'h10 ;
			data[24216] <= 8'h10 ;
			data[24217] <= 8'h10 ;
			data[24218] <= 8'h10 ;
			data[24219] <= 8'h10 ;
			data[24220] <= 8'h10 ;
			data[24221] <= 8'h10 ;
			data[24222] <= 8'h10 ;
			data[24223] <= 8'h10 ;
			data[24224] <= 8'h10 ;
			data[24225] <= 8'h10 ;
			data[24226] <= 8'h10 ;
			data[24227] <= 8'h10 ;
			data[24228] <= 8'h10 ;
			data[24229] <= 8'h10 ;
			data[24230] <= 8'h10 ;
			data[24231] <= 8'h10 ;
			data[24232] <= 8'h10 ;
			data[24233] <= 8'h10 ;
			data[24234] <= 8'h10 ;
			data[24235] <= 8'h10 ;
			data[24236] <= 8'h10 ;
			data[24237] <= 8'h10 ;
			data[24238] <= 8'h10 ;
			data[24239] <= 8'h10 ;
			data[24240] <= 8'h10 ;
			data[24241] <= 8'h10 ;
			data[24242] <= 8'h10 ;
			data[24243] <= 8'h10 ;
			data[24244] <= 8'h10 ;
			data[24245] <= 8'h10 ;
			data[24246] <= 8'h10 ;
			data[24247] <= 8'h10 ;
			data[24248] <= 8'h10 ;
			data[24249] <= 8'h10 ;
			data[24250] <= 8'h10 ;
			data[24251] <= 8'h10 ;
			data[24252] <= 8'h10 ;
			data[24253] <= 8'h10 ;
			data[24254] <= 8'h10 ;
			data[24255] <= 8'h10 ;
			data[24256] <= 8'h10 ;
			data[24257] <= 8'h10 ;
			data[24258] <= 8'h10 ;
			data[24259] <= 8'h10 ;
			data[24260] <= 8'h10 ;
			data[24261] <= 8'h10 ;
			data[24262] <= 8'h10 ;
			data[24263] <= 8'h10 ;
			data[24264] <= 8'h10 ;
			data[24265] <= 8'h10 ;
			data[24266] <= 8'h10 ;
			data[24267] <= 8'h10 ;
			data[24268] <= 8'h10 ;
			data[24269] <= 8'h10 ;
			data[24270] <= 8'h10 ;
			data[24271] <= 8'h10 ;
			data[24272] <= 8'h10 ;
			data[24273] <= 8'h10 ;
			data[24274] <= 8'h10 ;
			data[24275] <= 8'h10 ;
			data[24276] <= 8'h10 ;
			data[24277] <= 8'h10 ;
			data[24278] <= 8'h10 ;
			data[24279] <= 8'h10 ;
			data[24280] <= 8'h10 ;
			data[24281] <= 8'h10 ;
			data[24282] <= 8'h10 ;
			data[24283] <= 8'h10 ;
			data[24284] <= 8'h10 ;
			data[24285] <= 8'h10 ;
			data[24286] <= 8'h10 ;
			data[24287] <= 8'h10 ;
			data[24288] <= 8'h10 ;
			data[24289] <= 8'h10 ;
			data[24290] <= 8'h10 ;
			data[24291] <= 8'h10 ;
			data[24292] <= 8'h10 ;
			data[24293] <= 8'h10 ;
			data[24294] <= 8'h10 ;
			data[24295] <= 8'h10 ;
			data[24296] <= 8'h10 ;
			data[24297] <= 8'h10 ;
			data[24298] <= 8'h10 ;
			data[24299] <= 8'h10 ;
			data[24300] <= 8'h10 ;
			data[24301] <= 8'h10 ;
			data[24302] <= 8'h10 ;
			data[24303] <= 8'h10 ;
			data[24304] <= 8'h10 ;
			data[24305] <= 8'h10 ;
			data[24306] <= 8'h10 ;
			data[24307] <= 8'h10 ;
			data[24308] <= 8'h10 ;
			data[24309] <= 8'h10 ;
			data[24310] <= 8'h10 ;
			data[24311] <= 8'h10 ;
			data[24312] <= 8'h10 ;
			data[24313] <= 8'h10 ;
			data[24314] <= 8'h10 ;
			data[24315] <= 8'h10 ;
			data[24316] <= 8'h10 ;
			data[24317] <= 8'h10 ;
			data[24318] <= 8'h10 ;
			data[24319] <= 8'h10 ;
			data[24320] <= 8'h10 ;
			data[24321] <= 8'h10 ;
			data[24322] <= 8'h10 ;
			data[24323] <= 8'h10 ;
			data[24324] <= 8'h10 ;
			data[24325] <= 8'h10 ;
			data[24326] <= 8'h10 ;
			data[24327] <= 8'h10 ;
			data[24328] <= 8'h10 ;
			data[24329] <= 8'h10 ;
			data[24330] <= 8'h10 ;
			data[24331] <= 8'h10 ;
			data[24332] <= 8'h10 ;
			data[24333] <= 8'h10 ;
			data[24334] <= 8'h10 ;
			data[24335] <= 8'h10 ;
			data[24336] <= 8'h10 ;
			data[24337] <= 8'h10 ;
			data[24338] <= 8'h10 ;
			data[24339] <= 8'h10 ;
			data[24340] <= 8'h10 ;
			data[24341] <= 8'h10 ;
			data[24342] <= 8'h10 ;
			data[24343] <= 8'h10 ;
			data[24344] <= 8'h10 ;
			data[24345] <= 8'h10 ;
			data[24346] <= 8'h10 ;
			data[24347] <= 8'h10 ;
			data[24348] <= 8'h10 ;
			data[24349] <= 8'h10 ;
			data[24350] <= 8'h10 ;
			data[24351] <= 8'h10 ;
			data[24352] <= 8'h10 ;
			data[24353] <= 8'h10 ;
			data[24354] <= 8'h10 ;
			data[24355] <= 8'h10 ;
			data[24356] <= 8'h10 ;
			data[24357] <= 8'h10 ;
			data[24358] <= 8'h10 ;
			data[24359] <= 8'h10 ;
			data[24360] <= 8'h10 ;
			data[24361] <= 8'h10 ;
			data[24362] <= 8'h10 ;
			data[24363] <= 8'h10 ;
			data[24364] <= 8'h10 ;
			data[24365] <= 8'h10 ;
			data[24366] <= 8'h10 ;
			data[24367] <= 8'h10 ;
			data[24368] <= 8'h10 ;
			data[24369] <= 8'h10 ;
			data[24370] <= 8'h10 ;
			data[24371] <= 8'h10 ;
			data[24372] <= 8'h10 ;
			data[24373] <= 8'h10 ;
			data[24374] <= 8'h10 ;
			data[24375] <= 8'h10 ;
			data[24376] <= 8'h10 ;
			data[24377] <= 8'h10 ;
			data[24378] <= 8'h10 ;
			data[24379] <= 8'h10 ;
			data[24380] <= 8'h10 ;
			data[24381] <= 8'h10 ;
			data[24382] <= 8'h10 ;
			data[24383] <= 8'h10 ;
			data[24384] <= 8'h10 ;
			data[24385] <= 8'h10 ;
			data[24386] <= 8'h10 ;
			data[24387] <= 8'h10 ;
			data[24388] <= 8'h10 ;
			data[24389] <= 8'h10 ;
			data[24390] <= 8'h10 ;
			data[24391] <= 8'h10 ;
			data[24392] <= 8'h10 ;
			data[24393] <= 8'h10 ;
			data[24394] <= 8'h10 ;
			data[24395] <= 8'h10 ;
			data[24396] <= 8'h10 ;
			data[24397] <= 8'h10 ;
			data[24398] <= 8'h10 ;
			data[24399] <= 8'h10 ;
			data[24400] <= 8'h10 ;
			data[24401] <= 8'h10 ;
			data[24402] <= 8'h10 ;
			data[24403] <= 8'h10 ;
			data[24404] <= 8'h10 ;
			data[24405] <= 8'h10 ;
			data[24406] <= 8'h10 ;
			data[24407] <= 8'h10 ;
			data[24408] <= 8'h10 ;
			data[24409] <= 8'h10 ;
			data[24410] <= 8'h10 ;
			data[24411] <= 8'h10 ;
			data[24412] <= 8'h10 ;
			data[24413] <= 8'h10 ;
			data[24414] <= 8'h10 ;
			data[24415] <= 8'h10 ;
			data[24416] <= 8'h10 ;
			data[24417] <= 8'h10 ;
			data[24418] <= 8'h10 ;
			data[24419] <= 8'h10 ;
			data[24420] <= 8'h10 ;
			data[24421] <= 8'h10 ;
			data[24422] <= 8'h10 ;
			data[24423] <= 8'h10 ;
			data[24424] <= 8'h10 ;
			data[24425] <= 8'h10 ;
			data[24426] <= 8'h10 ;
			data[24427] <= 8'h10 ;
			data[24428] <= 8'h10 ;
			data[24429] <= 8'h10 ;
			data[24430] <= 8'h10 ;
			data[24431] <= 8'h10 ;
			data[24432] <= 8'h10 ;
			data[24433] <= 8'h10 ;
			data[24434] <= 8'h10 ;
			data[24435] <= 8'h10 ;
			data[24436] <= 8'h10 ;
			data[24437] <= 8'h10 ;
			data[24438] <= 8'h10 ;
			data[24439] <= 8'h10 ;
			data[24440] <= 8'h10 ;
			data[24441] <= 8'h10 ;
			data[24442] <= 8'h10 ;
			data[24443] <= 8'h10 ;
			data[24444] <= 8'h10 ;
			data[24445] <= 8'h10 ;
			data[24446] <= 8'h10 ;
			data[24447] <= 8'h10 ;
			data[24448] <= 8'h10 ;
			data[24449] <= 8'h10 ;
			data[24450] <= 8'h10 ;
			data[24451] <= 8'h10 ;
			data[24452] <= 8'h10 ;
			data[24453] <= 8'h10 ;
			data[24454] <= 8'h10 ;
			data[24455] <= 8'h10 ;
			data[24456] <= 8'h10 ;
			data[24457] <= 8'h10 ;
			data[24458] <= 8'h10 ;
			data[24459] <= 8'h10 ;
			data[24460] <= 8'h10 ;
			data[24461] <= 8'h10 ;
			data[24462] <= 8'h10 ;
			data[24463] <= 8'h10 ;
			data[24464] <= 8'h10 ;
			data[24465] <= 8'h10 ;
			data[24466] <= 8'h10 ;
			data[24467] <= 8'h10 ;
			data[24468] <= 8'h10 ;
			data[24469] <= 8'h10 ;
			data[24470] <= 8'h10 ;
			data[24471] <= 8'h10 ;
			data[24472] <= 8'h10 ;
			data[24473] <= 8'h10 ;
			data[24474] <= 8'h10 ;
			data[24475] <= 8'h10 ;
			data[24476] <= 8'h10 ;
			data[24477] <= 8'h10 ;
			data[24478] <= 8'h10 ;
			data[24479] <= 8'h10 ;
			data[24480] <= 8'h10 ;
			data[24481] <= 8'h10 ;
			data[24482] <= 8'h10 ;
			data[24483] <= 8'h10 ;
			data[24484] <= 8'h10 ;
			data[24485] <= 8'h10 ;
			data[24486] <= 8'h10 ;
			data[24487] <= 8'h10 ;
			data[24488] <= 8'h10 ;
			data[24489] <= 8'h10 ;
			data[24490] <= 8'h10 ;
			data[24491] <= 8'h10 ;
			data[24492] <= 8'h10 ;
			data[24493] <= 8'h10 ;
			data[24494] <= 8'h10 ;
			data[24495] <= 8'h10 ;
			data[24496] <= 8'h10 ;
			data[24497] <= 8'h10 ;
			data[24498] <= 8'h10 ;
			data[24499] <= 8'h10 ;
			data[24500] <= 8'h10 ;
			data[24501] <= 8'h10 ;
			data[24502] <= 8'h10 ;
			data[24503] <= 8'h10 ;
			data[24504] <= 8'h10 ;
			data[24505] <= 8'h10 ;
			data[24506] <= 8'h10 ;
			data[24507] <= 8'h10 ;
			data[24508] <= 8'h10 ;
			data[24509] <= 8'h10 ;
			data[24510] <= 8'h10 ;
			data[24511] <= 8'h10 ;
			data[24512] <= 8'h10 ;
			data[24513] <= 8'h10 ;
			data[24514] <= 8'h10 ;
			data[24515] <= 8'h10 ;
			data[24516] <= 8'h10 ;
			data[24517] <= 8'h10 ;
			data[24518] <= 8'h10 ;
			data[24519] <= 8'h10 ;
			data[24520] <= 8'h10 ;
			data[24521] <= 8'h10 ;
			data[24522] <= 8'h10 ;
			data[24523] <= 8'h10 ;
			data[24524] <= 8'h10 ;
			data[24525] <= 8'h10 ;
			data[24526] <= 8'h10 ;
			data[24527] <= 8'h10 ;
			data[24528] <= 8'h10 ;
			data[24529] <= 8'h10 ;
			data[24530] <= 8'h10 ;
			data[24531] <= 8'h10 ;
			data[24532] <= 8'h10 ;
			data[24533] <= 8'h10 ;
			data[24534] <= 8'h10 ;
			data[24535] <= 8'h10 ;
			data[24536] <= 8'h10 ;
			data[24537] <= 8'h10 ;
			data[24538] <= 8'h10 ;
			data[24539] <= 8'h10 ;
			data[24540] <= 8'h10 ;
			data[24541] <= 8'h10 ;
			data[24542] <= 8'h10 ;
			data[24543] <= 8'h10 ;
			data[24544] <= 8'h10 ;
			data[24545] <= 8'h10 ;
			data[24546] <= 8'h10 ;
			data[24547] <= 8'h10 ;
			data[24548] <= 8'h10 ;
			data[24549] <= 8'h10 ;
			data[24550] <= 8'h10 ;
			data[24551] <= 8'h10 ;
			data[24552] <= 8'h10 ;
			data[24553] <= 8'h10 ;
			data[24554] <= 8'h10 ;
			data[24555] <= 8'h10 ;
			data[24556] <= 8'h10 ;
			data[24557] <= 8'h10 ;
			data[24558] <= 8'h10 ;
			data[24559] <= 8'h10 ;
			data[24560] <= 8'h10 ;
			data[24561] <= 8'h10 ;
			data[24562] <= 8'h10 ;
			data[24563] <= 8'h10 ;
			data[24564] <= 8'h10 ;
			data[24565] <= 8'h10 ;
			data[24566] <= 8'h10 ;
			data[24567] <= 8'h10 ;
			data[24568] <= 8'h10 ;
			data[24569] <= 8'h10 ;
			data[24570] <= 8'h10 ;
			data[24571] <= 8'h10 ;
			data[24572] <= 8'h10 ;
			data[24573] <= 8'h10 ;
			data[24574] <= 8'h10 ;
			data[24575] <= 8'h10 ;
			data[24576] <= 8'h10 ;
			data[24577] <= 8'h10 ;
			data[24578] <= 8'h10 ;
			data[24579] <= 8'h10 ;
			data[24580] <= 8'h10 ;
			data[24581] <= 8'h10 ;
			data[24582] <= 8'h10 ;
			data[24583] <= 8'h10 ;
			data[24584] <= 8'h10 ;
			data[24585] <= 8'h10 ;
			data[24586] <= 8'h10 ;
			data[24587] <= 8'h10 ;
			data[24588] <= 8'h10 ;
			data[24589] <= 8'h10 ;
			data[24590] <= 8'h10 ;
			data[24591] <= 8'h10 ;
			data[24592] <= 8'h10 ;
			data[24593] <= 8'h10 ;
			data[24594] <= 8'h10 ;
			data[24595] <= 8'h10 ;
			data[24596] <= 8'h10 ;
			data[24597] <= 8'h10 ;
			data[24598] <= 8'h10 ;
			data[24599] <= 8'h10 ;
			data[24600] <= 8'h10 ;
			data[24601] <= 8'h10 ;
			data[24602] <= 8'h10 ;
			data[24603] <= 8'h10 ;
			data[24604] <= 8'h10 ;
			data[24605] <= 8'h10 ;
			data[24606] <= 8'h10 ;
			data[24607] <= 8'h10 ;
			data[24608] <= 8'h10 ;
			data[24609] <= 8'h10 ;
			data[24610] <= 8'h10 ;
			data[24611] <= 8'h10 ;
			data[24612] <= 8'h10 ;
			data[24613] <= 8'h10 ;
			data[24614] <= 8'h10 ;
			data[24615] <= 8'h10 ;
			data[24616] <= 8'h10 ;
			data[24617] <= 8'h10 ;
			data[24618] <= 8'h10 ;
			data[24619] <= 8'h10 ;
			data[24620] <= 8'h10 ;
			data[24621] <= 8'h10 ;
			data[24622] <= 8'h10 ;
			data[24623] <= 8'h10 ;
			data[24624] <= 8'h10 ;
			data[24625] <= 8'h10 ;
			data[24626] <= 8'h10 ;
			data[24627] <= 8'h10 ;
			data[24628] <= 8'h10 ;
			data[24629] <= 8'h10 ;
			data[24630] <= 8'h10 ;
			data[24631] <= 8'h10 ;
			data[24632] <= 8'h10 ;
			data[24633] <= 8'h10 ;
			data[24634] <= 8'h10 ;
			data[24635] <= 8'h10 ;
			data[24636] <= 8'h10 ;
			data[24637] <= 8'h10 ;
			data[24638] <= 8'h10 ;
			data[24639] <= 8'h10 ;
			data[24640] <= 8'h10 ;
			data[24641] <= 8'h10 ;
			data[24642] <= 8'h10 ;
			data[24643] <= 8'h10 ;
			data[24644] <= 8'h10 ;
			data[24645] <= 8'h10 ;
			data[24646] <= 8'h10 ;
			data[24647] <= 8'h10 ;
			data[24648] <= 8'h10 ;
			data[24649] <= 8'h10 ;
			data[24650] <= 8'h10 ;
			data[24651] <= 8'h10 ;
			data[24652] <= 8'h10 ;
			data[24653] <= 8'h10 ;
			data[24654] <= 8'h10 ;
			data[24655] <= 8'h10 ;
			data[24656] <= 8'h10 ;
			data[24657] <= 8'h10 ;
			data[24658] <= 8'h10 ;
			data[24659] <= 8'h10 ;
			data[24660] <= 8'h10 ;
			data[24661] <= 8'h10 ;
			data[24662] <= 8'h10 ;
			data[24663] <= 8'h10 ;
			data[24664] <= 8'h10 ;
			data[24665] <= 8'h10 ;
			data[24666] <= 8'h10 ;
			data[24667] <= 8'h10 ;
			data[24668] <= 8'h10 ;
			data[24669] <= 8'h10 ;
			data[24670] <= 8'h10 ;
			data[24671] <= 8'h10 ;
			data[24672] <= 8'h10 ;
			data[24673] <= 8'h10 ;
			data[24674] <= 8'h10 ;
			data[24675] <= 8'h10 ;
			data[24676] <= 8'h10 ;
			data[24677] <= 8'h10 ;
			data[24678] <= 8'h10 ;
			data[24679] <= 8'h10 ;
			data[24680] <= 8'h10 ;
			data[24681] <= 8'h10 ;
			data[24682] <= 8'h10 ;
			data[24683] <= 8'h10 ;
			data[24684] <= 8'h10 ;
			data[24685] <= 8'h10 ;
			data[24686] <= 8'h10 ;
			data[24687] <= 8'h10 ;
			data[24688] <= 8'h10 ;
			data[24689] <= 8'h10 ;
			data[24690] <= 8'h10 ;
			data[24691] <= 8'h10 ;
			data[24692] <= 8'h10 ;
			data[24693] <= 8'h10 ;
			data[24694] <= 8'h10 ;
			data[24695] <= 8'h10 ;
			data[24696] <= 8'h10 ;
			data[24697] <= 8'h10 ;
			data[24698] <= 8'h10 ;
			data[24699] <= 8'h10 ;
			data[24700] <= 8'h10 ;
			data[24701] <= 8'h10 ;
			data[24702] <= 8'h10 ;
			data[24703] <= 8'h10 ;
			data[24704] <= 8'h10 ;
			data[24705] <= 8'h10 ;
			data[24706] <= 8'h10 ;
			data[24707] <= 8'h10 ;
			data[24708] <= 8'h10 ;
			data[24709] <= 8'h10 ;
			data[24710] <= 8'h10 ;
			data[24711] <= 8'h10 ;
			data[24712] <= 8'h10 ;
			data[24713] <= 8'h10 ;
			data[24714] <= 8'h10 ;
			data[24715] <= 8'h10 ;
			data[24716] <= 8'h10 ;
			data[24717] <= 8'h10 ;
			data[24718] <= 8'h10 ;
			data[24719] <= 8'h10 ;
			data[24720] <= 8'h10 ;
			data[24721] <= 8'h10 ;
			data[24722] <= 8'h10 ;
			data[24723] <= 8'h10 ;
			data[24724] <= 8'h10 ;
			data[24725] <= 8'h10 ;
			data[24726] <= 8'h10 ;
			data[24727] <= 8'h10 ;
			data[24728] <= 8'h10 ;
			data[24729] <= 8'h10 ;
			data[24730] <= 8'h10 ;
			data[24731] <= 8'h10 ;
			data[24732] <= 8'h10 ;
			data[24733] <= 8'h10 ;
			data[24734] <= 8'h10 ;
			data[24735] <= 8'h10 ;
			data[24736] <= 8'h10 ;
			data[24737] <= 8'h10 ;
			data[24738] <= 8'h10 ;
			data[24739] <= 8'h10 ;
			data[24740] <= 8'h10 ;
			data[24741] <= 8'h10 ;
			data[24742] <= 8'h10 ;
			data[24743] <= 8'h10 ;
			data[24744] <= 8'h10 ;
			data[24745] <= 8'h10 ;
			data[24746] <= 8'h10 ;
			data[24747] <= 8'h10 ;
			data[24748] <= 8'h10 ;
			data[24749] <= 8'h10 ;
			data[24750] <= 8'h10 ;
			data[24751] <= 8'h10 ;
			data[24752] <= 8'h10 ;
			data[24753] <= 8'h10 ;
			data[24754] <= 8'h10 ;
			data[24755] <= 8'h10 ;
			data[24756] <= 8'h10 ;
			data[24757] <= 8'h10 ;
			data[24758] <= 8'h10 ;
			data[24759] <= 8'h10 ;
			data[24760] <= 8'h10 ;
			data[24761] <= 8'h10 ;
			data[24762] <= 8'h10 ;
			data[24763] <= 8'h10 ;
			data[24764] <= 8'h10 ;
			data[24765] <= 8'h10 ;
			data[24766] <= 8'h10 ;
			data[24767] <= 8'h10 ;
			data[24768] <= 8'h10 ;
			data[24769] <= 8'h10 ;
			data[24770] <= 8'h10 ;
			data[24771] <= 8'h10 ;
			data[24772] <= 8'h10 ;
			data[24773] <= 8'h10 ;
			data[24774] <= 8'h10 ;
			data[24775] <= 8'h10 ;
			data[24776] <= 8'h10 ;
			data[24777] <= 8'h10 ;
			data[24778] <= 8'h10 ;
			data[24779] <= 8'h10 ;
			data[24780] <= 8'h10 ;
			data[24781] <= 8'h10 ;
			data[24782] <= 8'h10 ;
			data[24783] <= 8'h10 ;
			data[24784] <= 8'h10 ;
			data[24785] <= 8'h10 ;
			data[24786] <= 8'h10 ;
			data[24787] <= 8'h10 ;
			data[24788] <= 8'h10 ;
			data[24789] <= 8'h10 ;
			data[24790] <= 8'h10 ;
			data[24791] <= 8'h10 ;
			data[24792] <= 8'h10 ;
			data[24793] <= 8'h10 ;
			data[24794] <= 8'h10 ;
			data[24795] <= 8'h10 ;
			data[24796] <= 8'h10 ;
			data[24797] <= 8'h10 ;
			data[24798] <= 8'h10 ;
			data[24799] <= 8'h10 ;
			data[24800] <= 8'h10 ;
			data[24801] <= 8'h10 ;
			data[24802] <= 8'h10 ;
			data[24803] <= 8'h10 ;
			data[24804] <= 8'h10 ;
			data[24805] <= 8'h10 ;
			data[24806] <= 8'h10 ;
			data[24807] <= 8'h10 ;
			data[24808] <= 8'h10 ;
			data[24809] <= 8'h10 ;
			data[24810] <= 8'h10 ;
			data[24811] <= 8'h10 ;
			data[24812] <= 8'h10 ;
			data[24813] <= 8'h10 ;
			data[24814] <= 8'h10 ;
			data[24815] <= 8'h10 ;
			data[24816] <= 8'h10 ;
			data[24817] <= 8'h10 ;
			data[24818] <= 8'h10 ;
			data[24819] <= 8'h10 ;
			data[24820] <= 8'h10 ;
			data[24821] <= 8'h10 ;
			data[24822] <= 8'h10 ;
			data[24823] <= 8'h10 ;
			data[24824] <= 8'h10 ;
			data[24825] <= 8'h10 ;
			data[24826] <= 8'h10 ;
			data[24827] <= 8'h10 ;
			data[24828] <= 8'h10 ;
			data[24829] <= 8'h10 ;
			data[24830] <= 8'h10 ;
			data[24831] <= 8'h10 ;
			data[24832] <= 8'h10 ;
			data[24833] <= 8'h10 ;
			data[24834] <= 8'h10 ;
			data[24835] <= 8'h10 ;
			data[24836] <= 8'h10 ;
			data[24837] <= 8'h10 ;
			data[24838] <= 8'h10 ;
			data[24839] <= 8'h10 ;
			data[24840] <= 8'h10 ;
			data[24841] <= 8'h10 ;
			data[24842] <= 8'h10 ;
			data[24843] <= 8'h10 ;
			data[24844] <= 8'h10 ;
			data[24845] <= 8'h10 ;
			data[24846] <= 8'h10 ;
			data[24847] <= 8'h10 ;
			data[24848] <= 8'h10 ;
			data[24849] <= 8'h10 ;
			data[24850] <= 8'h10 ;
			data[24851] <= 8'h10 ;
			data[24852] <= 8'h10 ;
			data[24853] <= 8'h10 ;
			data[24854] <= 8'h10 ;
			data[24855] <= 8'h10 ;
			data[24856] <= 8'h10 ;
			data[24857] <= 8'h10 ;
			data[24858] <= 8'h10 ;
			data[24859] <= 8'h10 ;
			data[24860] <= 8'h10 ;
			data[24861] <= 8'h10 ;
			data[24862] <= 8'h10 ;
			data[24863] <= 8'h10 ;
			data[24864] <= 8'h10 ;
			data[24865] <= 8'h10 ;
			data[24866] <= 8'h10 ;
			data[24867] <= 8'h10 ;
			data[24868] <= 8'h10 ;
			data[24869] <= 8'h10 ;
			data[24870] <= 8'h10 ;
			data[24871] <= 8'h10 ;
			data[24872] <= 8'h10 ;
			data[24873] <= 8'h10 ;
			data[24874] <= 8'h10 ;
			data[24875] <= 8'h10 ;
			data[24876] <= 8'h10 ;
			data[24877] <= 8'h10 ;
			data[24878] <= 8'h10 ;
			data[24879] <= 8'h10 ;
			data[24880] <= 8'h10 ;
			data[24881] <= 8'h10 ;
			data[24882] <= 8'h10 ;
			data[24883] <= 8'h10 ;
			data[24884] <= 8'h10 ;
			data[24885] <= 8'h10 ;
			data[24886] <= 8'h10 ;
			data[24887] <= 8'h10 ;
			data[24888] <= 8'h10 ;
			data[24889] <= 8'h10 ;
			data[24890] <= 8'h10 ;
			data[24891] <= 8'h10 ;
			data[24892] <= 8'h10 ;
			data[24893] <= 8'h10 ;
			data[24894] <= 8'h10 ;
			data[24895] <= 8'h10 ;
			data[24896] <= 8'h10 ;
			data[24897] <= 8'h10 ;
			data[24898] <= 8'h10 ;
			data[24899] <= 8'h10 ;
			data[24900] <= 8'h10 ;
			data[24901] <= 8'h10 ;
			data[24902] <= 8'h10 ;
			data[24903] <= 8'h10 ;
			data[24904] <= 8'h10 ;
			data[24905] <= 8'h10 ;
			data[24906] <= 8'h10 ;
			data[24907] <= 8'h10 ;
			data[24908] <= 8'h10 ;
			data[24909] <= 8'h10 ;
			data[24910] <= 8'h10 ;
			data[24911] <= 8'h10 ;
			data[24912] <= 8'h10 ;
			data[24913] <= 8'h10 ;
			data[24914] <= 8'h10 ;
			data[24915] <= 8'h10 ;
			data[24916] <= 8'h10 ;
			data[24917] <= 8'h10 ;
			data[24918] <= 8'h10 ;
			data[24919] <= 8'h10 ;
			data[24920] <= 8'h10 ;
			data[24921] <= 8'h10 ;
			data[24922] <= 8'h10 ;
			data[24923] <= 8'h10 ;
			data[24924] <= 8'h10 ;
			data[24925] <= 8'h10 ;
			data[24926] <= 8'h10 ;
			data[24927] <= 8'h10 ;
			data[24928] <= 8'h10 ;
			data[24929] <= 8'h10 ;
			data[24930] <= 8'h10 ;
			data[24931] <= 8'h10 ;
			data[24932] <= 8'h10 ;
			data[24933] <= 8'h10 ;
			data[24934] <= 8'h10 ;
			data[24935] <= 8'h10 ;
			data[24936] <= 8'h10 ;
			data[24937] <= 8'h10 ;
			data[24938] <= 8'h10 ;
			data[24939] <= 8'h10 ;
			data[24940] <= 8'h10 ;
			data[24941] <= 8'h10 ;
			data[24942] <= 8'h10 ;
			data[24943] <= 8'h10 ;
			data[24944] <= 8'h10 ;
			data[24945] <= 8'h10 ;
			data[24946] <= 8'h10 ;
			data[24947] <= 8'h10 ;
			data[24948] <= 8'h10 ;
			data[24949] <= 8'h10 ;
			data[24950] <= 8'h10 ;
			data[24951] <= 8'h10 ;
			data[24952] <= 8'h10 ;
			data[24953] <= 8'h10 ;
			data[24954] <= 8'h10 ;
			data[24955] <= 8'h10 ;
			data[24956] <= 8'h10 ;
			data[24957] <= 8'h10 ;
			data[24958] <= 8'h10 ;
			data[24959] <= 8'h10 ;
			data[24960] <= 8'h10 ;
			data[24961] <= 8'h10 ;
			data[24962] <= 8'h10 ;
			data[24963] <= 8'h10 ;
			data[24964] <= 8'h10 ;
			data[24965] <= 8'h10 ;
			data[24966] <= 8'h10 ;
			data[24967] <= 8'h10 ;
			data[24968] <= 8'h10 ;
			data[24969] <= 8'h10 ;
			data[24970] <= 8'h10 ;
			data[24971] <= 8'h10 ;
			data[24972] <= 8'h10 ;
			data[24973] <= 8'h10 ;
			data[24974] <= 8'h10 ;
			data[24975] <= 8'h10 ;
			data[24976] <= 8'h10 ;
			data[24977] <= 8'h10 ;
			data[24978] <= 8'h10 ;
			data[24979] <= 8'h10 ;
			data[24980] <= 8'h10 ;
			data[24981] <= 8'h10 ;
			data[24982] <= 8'h10 ;
			data[24983] <= 8'h10 ;
			data[24984] <= 8'h10 ;
			data[24985] <= 8'h10 ;
			data[24986] <= 8'h10 ;
			data[24987] <= 8'h10 ;
			data[24988] <= 8'h10 ;
			data[24989] <= 8'h10 ;
			data[24990] <= 8'h10 ;
			data[24991] <= 8'h10 ;
			data[24992] <= 8'h10 ;
			data[24993] <= 8'h10 ;
			data[24994] <= 8'h10 ;
			data[24995] <= 8'h10 ;
			data[24996] <= 8'h10 ;
			data[24997] <= 8'h10 ;
			data[24998] <= 8'h10 ;
			data[24999] <= 8'h10 ;
			data[25000] <= 8'h10 ;
			data[25001] <= 8'h10 ;
			data[25002] <= 8'h10 ;
			data[25003] <= 8'h10 ;
			data[25004] <= 8'h10 ;
			data[25005] <= 8'h10 ;
			data[25006] <= 8'h10 ;
			data[25007] <= 8'h10 ;
			data[25008] <= 8'h10 ;
			data[25009] <= 8'h10 ;
			data[25010] <= 8'h10 ;
			data[25011] <= 8'h10 ;
			data[25012] <= 8'h10 ;
			data[25013] <= 8'h10 ;
			data[25014] <= 8'h10 ;
			data[25015] <= 8'h10 ;
			data[25016] <= 8'h10 ;
			data[25017] <= 8'h10 ;
			data[25018] <= 8'h10 ;
			data[25019] <= 8'h10 ;
			data[25020] <= 8'h10 ;
			data[25021] <= 8'h10 ;
			data[25022] <= 8'h10 ;
			data[25023] <= 8'h10 ;
			data[25024] <= 8'h10 ;
			data[25025] <= 8'h10 ;
			data[25026] <= 8'h10 ;
			data[25027] <= 8'h10 ;
			data[25028] <= 8'h10 ;
			data[25029] <= 8'h10 ;
			data[25030] <= 8'h10 ;
			data[25031] <= 8'h10 ;
			data[25032] <= 8'h10 ;
			data[25033] <= 8'h10 ;
			data[25034] <= 8'h10 ;
			data[25035] <= 8'h10 ;
			data[25036] <= 8'h10 ;
			data[25037] <= 8'h10 ;
			data[25038] <= 8'h10 ;
			data[25039] <= 8'h10 ;
			data[25040] <= 8'h10 ;
			data[25041] <= 8'h10 ;
			data[25042] <= 8'h10 ;
			data[25043] <= 8'h10 ;
			data[25044] <= 8'h10 ;
			data[25045] <= 8'h10 ;
			data[25046] <= 8'h10 ;
			data[25047] <= 8'h10 ;
			data[25048] <= 8'h10 ;
			data[25049] <= 8'h10 ;
			data[25050] <= 8'h10 ;
			data[25051] <= 8'h10 ;
			data[25052] <= 8'h10 ;
			data[25053] <= 8'h10 ;
			data[25054] <= 8'h10 ;
			data[25055] <= 8'h10 ;
			data[25056] <= 8'h10 ;
			data[25057] <= 8'h10 ;
			data[25058] <= 8'h10 ;
			data[25059] <= 8'h10 ;
			data[25060] <= 8'h10 ;
			data[25061] <= 8'h10 ;
			data[25062] <= 8'h10 ;
			data[25063] <= 8'h10 ;
			data[25064] <= 8'h10 ;
			data[25065] <= 8'h10 ;
			data[25066] <= 8'h10 ;
			data[25067] <= 8'h10 ;
			data[25068] <= 8'h10 ;
			data[25069] <= 8'h10 ;
			data[25070] <= 8'h10 ;
			data[25071] <= 8'h10 ;
			data[25072] <= 8'h10 ;
			data[25073] <= 8'h10 ;
			data[25074] <= 8'h10 ;
			data[25075] <= 8'h10 ;
			data[25076] <= 8'h10 ;
			data[25077] <= 8'h10 ;
			data[25078] <= 8'h10 ;
			data[25079] <= 8'h10 ;
			data[25080] <= 8'h10 ;
			data[25081] <= 8'h10 ;
			data[25082] <= 8'h10 ;
			data[25083] <= 8'h10 ;
			data[25084] <= 8'h10 ;
			data[25085] <= 8'h10 ;
			data[25086] <= 8'h10 ;
			data[25087] <= 8'h10 ;
			data[25088] <= 8'h10 ;
			data[25089] <= 8'h10 ;
			data[25090] <= 8'h10 ;
			data[25091] <= 8'h10 ;
			data[25092] <= 8'h10 ;
			data[25093] <= 8'h10 ;
			data[25094] <= 8'h10 ;
			data[25095] <= 8'h10 ;
			data[25096] <= 8'h10 ;
			data[25097] <= 8'h10 ;
			data[25098] <= 8'h10 ;
			data[25099] <= 8'h10 ;
			data[25100] <= 8'h10 ;
			data[25101] <= 8'h10 ;
			data[25102] <= 8'h10 ;
			data[25103] <= 8'h10 ;
			data[25104] <= 8'h10 ;
			data[25105] <= 8'h10 ;
			data[25106] <= 8'h10 ;
			data[25107] <= 8'h10 ;
			data[25108] <= 8'h10 ;
			data[25109] <= 8'h10 ;
			data[25110] <= 8'h10 ;
			data[25111] <= 8'h10 ;
			data[25112] <= 8'h10 ;
			data[25113] <= 8'h10 ;
			data[25114] <= 8'h10 ;
			data[25115] <= 8'h10 ;
			data[25116] <= 8'h10 ;
			data[25117] <= 8'h10 ;
			data[25118] <= 8'h10 ;
			data[25119] <= 8'h10 ;
			data[25120] <= 8'h10 ;
			data[25121] <= 8'h10 ;
			data[25122] <= 8'h10 ;
			data[25123] <= 8'h10 ;
			data[25124] <= 8'h10 ;
			data[25125] <= 8'h10 ;
			data[25126] <= 8'h10 ;
			data[25127] <= 8'h10 ;
			data[25128] <= 8'h10 ;
			data[25129] <= 8'h10 ;
			data[25130] <= 8'h10 ;
			data[25131] <= 8'h10 ;
			data[25132] <= 8'h10 ;
			data[25133] <= 8'h10 ;
			data[25134] <= 8'h10 ;
			data[25135] <= 8'h10 ;
			data[25136] <= 8'h10 ;
			data[25137] <= 8'h10 ;
			data[25138] <= 8'h10 ;
			data[25139] <= 8'h10 ;
			data[25140] <= 8'h10 ;
			data[25141] <= 8'h10 ;
			data[25142] <= 8'h10 ;
			data[25143] <= 8'h10 ;
			data[25144] <= 8'h10 ;
			data[25145] <= 8'h10 ;
			data[25146] <= 8'h10 ;
			data[25147] <= 8'h10 ;
			data[25148] <= 8'h10 ;
			data[25149] <= 8'h10 ;
			data[25150] <= 8'h10 ;
			data[25151] <= 8'h10 ;
			data[25152] <= 8'h10 ;
			data[25153] <= 8'h10 ;
			data[25154] <= 8'h10 ;
			data[25155] <= 8'h10 ;
			data[25156] <= 8'h10 ;
			data[25157] <= 8'h10 ;
			data[25158] <= 8'h10 ;
			data[25159] <= 8'h10 ;
			data[25160] <= 8'h10 ;
			data[25161] <= 8'h10 ;
			data[25162] <= 8'h10 ;
			data[25163] <= 8'h10 ;
			data[25164] <= 8'h10 ;
			data[25165] <= 8'h10 ;
			data[25166] <= 8'h10 ;
			data[25167] <= 8'h10 ;
			data[25168] <= 8'h10 ;
			data[25169] <= 8'h10 ;
			data[25170] <= 8'h10 ;
			data[25171] <= 8'h10 ;
			data[25172] <= 8'h10 ;
			data[25173] <= 8'h10 ;
			data[25174] <= 8'h10 ;
			data[25175] <= 8'h10 ;
			data[25176] <= 8'h10 ;
			data[25177] <= 8'h10 ;
			data[25178] <= 8'h10 ;
			data[25179] <= 8'h10 ;
			data[25180] <= 8'h10 ;
			data[25181] <= 8'h10 ;
			data[25182] <= 8'h10 ;
			data[25183] <= 8'h10 ;
			data[25184] <= 8'h10 ;
			data[25185] <= 8'h10 ;
			data[25186] <= 8'h10 ;
			data[25187] <= 8'h10 ;
			data[25188] <= 8'h10 ;
			data[25189] <= 8'h10 ;
			data[25190] <= 8'h10 ;
			data[25191] <= 8'h10 ;
			data[25192] <= 8'h10 ;
			data[25193] <= 8'h10 ;
			data[25194] <= 8'h10 ;
			data[25195] <= 8'h10 ;
			data[25196] <= 8'h10 ;
			data[25197] <= 8'h10 ;
			data[25198] <= 8'h10 ;
			data[25199] <= 8'h10 ;
			data[25200] <= 8'h10 ;
			data[25201] <= 8'h10 ;
			data[25202] <= 8'h10 ;
			data[25203] <= 8'h10 ;
			data[25204] <= 8'h10 ;
			data[25205] <= 8'h10 ;
			data[25206] <= 8'h10 ;
			data[25207] <= 8'h10 ;
			data[25208] <= 8'h10 ;
			data[25209] <= 8'h10 ;
			data[25210] <= 8'h10 ;
			data[25211] <= 8'h10 ;
			data[25212] <= 8'h10 ;
			data[25213] <= 8'h10 ;
			data[25214] <= 8'h10 ;
			data[25215] <= 8'h10 ;
			data[25216] <= 8'h10 ;
			data[25217] <= 8'h10 ;
			data[25218] <= 8'h10 ;
			data[25219] <= 8'h10 ;
			data[25220] <= 8'h10 ;
			data[25221] <= 8'h10 ;
			data[25222] <= 8'h10 ;
			data[25223] <= 8'h10 ;
			data[25224] <= 8'h10 ;
			data[25225] <= 8'h10 ;
			data[25226] <= 8'h10 ;
			data[25227] <= 8'h10 ;
			data[25228] <= 8'h10 ;
			data[25229] <= 8'h10 ;
			data[25230] <= 8'h10 ;
			data[25231] <= 8'h10 ;
			data[25232] <= 8'h10 ;
			data[25233] <= 8'h10 ;
			data[25234] <= 8'h10 ;
			data[25235] <= 8'h10 ;
			data[25236] <= 8'h10 ;
			data[25237] <= 8'h10 ;
			data[25238] <= 8'h10 ;
			data[25239] <= 8'h10 ;
			data[25240] <= 8'h10 ;
			data[25241] <= 8'h10 ;
			data[25242] <= 8'h10 ;
			data[25243] <= 8'h10 ;
			data[25244] <= 8'h10 ;
			data[25245] <= 8'h10 ;
			data[25246] <= 8'h10 ;
			data[25247] <= 8'h10 ;
			data[25248] <= 8'h10 ;
			data[25249] <= 8'h10 ;
			data[25250] <= 8'h10 ;
			data[25251] <= 8'h10 ;
			data[25252] <= 8'h10 ;
			data[25253] <= 8'h10 ;
			data[25254] <= 8'h10 ;
			data[25255] <= 8'h10 ;
			data[25256] <= 8'h10 ;
			data[25257] <= 8'h10 ;
			data[25258] <= 8'h10 ;
			data[25259] <= 8'h10 ;
			data[25260] <= 8'h10 ;
			data[25261] <= 8'h10 ;
			data[25262] <= 8'h10 ;
			data[25263] <= 8'h10 ;
			data[25264] <= 8'h10 ;
			data[25265] <= 8'h10 ;
			data[25266] <= 8'h10 ;
			data[25267] <= 8'h10 ;
			data[25268] <= 8'h10 ;
			data[25269] <= 8'h10 ;
			data[25270] <= 8'h10 ;
			data[25271] <= 8'h10 ;
			data[25272] <= 8'h10 ;
			data[25273] <= 8'h10 ;
			data[25274] <= 8'h10 ;
			data[25275] <= 8'h10 ;
			data[25276] <= 8'h10 ;
			data[25277] <= 8'h10 ;
			data[25278] <= 8'h10 ;
			data[25279] <= 8'h10 ;
			data[25280] <= 8'h10 ;
			data[25281] <= 8'h10 ;
			data[25282] <= 8'h10 ;
			data[25283] <= 8'h10 ;
			data[25284] <= 8'h10 ;
			data[25285] <= 8'h10 ;
			data[25286] <= 8'h10 ;
			data[25287] <= 8'h10 ;
			data[25288] <= 8'h10 ;
			data[25289] <= 8'h10 ;
			data[25290] <= 8'h10 ;
			data[25291] <= 8'h10 ;
			data[25292] <= 8'h10 ;
			data[25293] <= 8'h10 ;
			data[25294] <= 8'h10 ;
			data[25295] <= 8'h10 ;
			data[25296] <= 8'h10 ;
			data[25297] <= 8'h10 ;
			data[25298] <= 8'h10 ;
			data[25299] <= 8'h10 ;
			data[25300] <= 8'h10 ;
			data[25301] <= 8'h10 ;
			data[25302] <= 8'h10 ;
			data[25303] <= 8'h10 ;
			data[25304] <= 8'h10 ;
			data[25305] <= 8'h10 ;
			data[25306] <= 8'h10 ;
			data[25307] <= 8'h10 ;
			data[25308] <= 8'h10 ;
			data[25309] <= 8'h10 ;
			data[25310] <= 8'h10 ;
			data[25311] <= 8'h10 ;
			data[25312] <= 8'h10 ;
			data[25313] <= 8'h10 ;
			data[25314] <= 8'h10 ;
			data[25315] <= 8'h10 ;
			data[25316] <= 8'h10 ;
			data[25317] <= 8'h10 ;
			data[25318] <= 8'h10 ;
			data[25319] <= 8'h10 ;
			data[25320] <= 8'h10 ;
			data[25321] <= 8'h10 ;
			data[25322] <= 8'h10 ;
			data[25323] <= 8'h10 ;
			data[25324] <= 8'h10 ;
			data[25325] <= 8'h10 ;
			data[25326] <= 8'h10 ;
			data[25327] <= 8'h10 ;
			data[25328] <= 8'h10 ;
			data[25329] <= 8'h10 ;
			data[25330] <= 8'h10 ;
			data[25331] <= 8'h10 ;
			data[25332] <= 8'h10 ;
			data[25333] <= 8'h10 ;
			data[25334] <= 8'h10 ;
			data[25335] <= 8'h10 ;
			data[25336] <= 8'h10 ;
			data[25337] <= 8'h10 ;
			data[25338] <= 8'h10 ;
			data[25339] <= 8'h10 ;
			data[25340] <= 8'h10 ;
			data[25341] <= 8'h10 ;
			data[25342] <= 8'h10 ;
			data[25343] <= 8'h10 ;
			data[25344] <= 8'h10 ;
			data[25345] <= 8'h10 ;
			data[25346] <= 8'h10 ;
			data[25347] <= 8'h10 ;
			data[25348] <= 8'h10 ;
			data[25349] <= 8'h10 ;
			data[25350] <= 8'h10 ;
			data[25351] <= 8'h10 ;
			data[25352] <= 8'h10 ;
			data[25353] <= 8'h10 ;
			data[25354] <= 8'h10 ;
			data[25355] <= 8'h10 ;
			data[25356] <= 8'h10 ;
			data[25357] <= 8'h10 ;
			data[25358] <= 8'h10 ;
			data[25359] <= 8'h10 ;
			data[25360] <= 8'h10 ;
			data[25361] <= 8'h10 ;
			data[25362] <= 8'h10 ;
			data[25363] <= 8'h10 ;
			data[25364] <= 8'h10 ;
			data[25365] <= 8'h10 ;
			data[25366] <= 8'h10 ;
			data[25367] <= 8'h10 ;
			data[25368] <= 8'h10 ;
			data[25369] <= 8'h10 ;
			data[25370] <= 8'h10 ;
			data[25371] <= 8'h10 ;
			data[25372] <= 8'h10 ;
			data[25373] <= 8'h10 ;
			data[25374] <= 8'h10 ;
			data[25375] <= 8'h10 ;
			data[25376] <= 8'h10 ;
			data[25377] <= 8'h10 ;
			data[25378] <= 8'h10 ;
			data[25379] <= 8'h10 ;
			data[25380] <= 8'h10 ;
			data[25381] <= 8'h10 ;
			data[25382] <= 8'h10 ;
			data[25383] <= 8'h10 ;
			data[25384] <= 8'h10 ;
			data[25385] <= 8'h10 ;
			data[25386] <= 8'h10 ;
			data[25387] <= 8'h10 ;
			data[25388] <= 8'h10 ;
			data[25389] <= 8'h10 ;
			data[25390] <= 8'h10 ;
			data[25391] <= 8'h10 ;
			data[25392] <= 8'h10 ;
			data[25393] <= 8'h10 ;
			data[25394] <= 8'h10 ;
			data[25395] <= 8'h10 ;
			data[25396] <= 8'h10 ;
			data[25397] <= 8'h10 ;
			data[25398] <= 8'h10 ;
			data[25399] <= 8'h10 ;
			data[25400] <= 8'h10 ;
			data[25401] <= 8'h10 ;
			data[25402] <= 8'h10 ;
			data[25403] <= 8'h10 ;
			data[25404] <= 8'h10 ;
			data[25405] <= 8'h10 ;
			data[25406] <= 8'h10 ;
			data[25407] <= 8'h10 ;
			data[25408] <= 8'h10 ;
			data[25409] <= 8'h10 ;
			data[25410] <= 8'h10 ;
			data[25411] <= 8'h10 ;
			data[25412] <= 8'h10 ;
			data[25413] <= 8'h10 ;
			data[25414] <= 8'h10 ;
			data[25415] <= 8'h10 ;
			data[25416] <= 8'h10 ;
			data[25417] <= 8'h10 ;
			data[25418] <= 8'h10 ;
			data[25419] <= 8'h10 ;
			data[25420] <= 8'h10 ;
			data[25421] <= 8'h10 ;
			data[25422] <= 8'h10 ;
			data[25423] <= 8'h10 ;
			data[25424] <= 8'h10 ;
			data[25425] <= 8'h10 ;
			data[25426] <= 8'h10 ;
			data[25427] <= 8'h10 ;
			data[25428] <= 8'h10 ;
			data[25429] <= 8'h10 ;
			data[25430] <= 8'h10 ;
			data[25431] <= 8'h10 ;
			data[25432] <= 8'h10 ;
			data[25433] <= 8'h10 ;
			data[25434] <= 8'h10 ;
			data[25435] <= 8'h10 ;
			data[25436] <= 8'h10 ;
			data[25437] <= 8'h10 ;
			data[25438] <= 8'h10 ;
			data[25439] <= 8'h10 ;
			data[25440] <= 8'h10 ;
			data[25441] <= 8'h10 ;
			data[25442] <= 8'h10 ;
			data[25443] <= 8'h10 ;
			data[25444] <= 8'h10 ;
			data[25445] <= 8'h10 ;
			data[25446] <= 8'h10 ;
			data[25447] <= 8'h10 ;
			data[25448] <= 8'h10 ;
			data[25449] <= 8'h10 ;
			data[25450] <= 8'h10 ;
			data[25451] <= 8'h10 ;
			data[25452] <= 8'h10 ;
			data[25453] <= 8'h10 ;
			data[25454] <= 8'h10 ;
			data[25455] <= 8'h10 ;
			data[25456] <= 8'h10 ;
			data[25457] <= 8'h10 ;
			data[25458] <= 8'h10 ;
			data[25459] <= 8'h10 ;
			data[25460] <= 8'h10 ;
			data[25461] <= 8'h10 ;
			data[25462] <= 8'h10 ;
			data[25463] <= 8'h10 ;
			data[25464] <= 8'h10 ;
			data[25465] <= 8'h10 ;
			data[25466] <= 8'h10 ;
			data[25467] <= 8'h10 ;
			data[25468] <= 8'h10 ;
			data[25469] <= 8'h10 ;
			data[25470] <= 8'h10 ;
			data[25471] <= 8'h10 ;
			data[25472] <= 8'h10 ;
			data[25473] <= 8'h10 ;
			data[25474] <= 8'h10 ;
			data[25475] <= 8'h10 ;
			data[25476] <= 8'h10 ;
			data[25477] <= 8'h10 ;
			data[25478] <= 8'h10 ;
			data[25479] <= 8'h10 ;
			data[25480] <= 8'h10 ;
			data[25481] <= 8'h10 ;
			data[25482] <= 8'h10 ;
			data[25483] <= 8'h10 ;
			data[25484] <= 8'h10 ;
			data[25485] <= 8'h10 ;
			data[25486] <= 8'h10 ;
			data[25487] <= 8'h10 ;
			data[25488] <= 8'h10 ;
			data[25489] <= 8'h10 ;
			data[25490] <= 8'h10 ;
			data[25491] <= 8'h10 ;
			data[25492] <= 8'h10 ;
			data[25493] <= 8'h10 ;
			data[25494] <= 8'h10 ;
			data[25495] <= 8'h10 ;
			data[25496] <= 8'h10 ;
			data[25497] <= 8'h10 ;
			data[25498] <= 8'h10 ;
			data[25499] <= 8'h10 ;
			data[25500] <= 8'h10 ;
			data[25501] <= 8'h10 ;
			data[25502] <= 8'h10 ;
			data[25503] <= 8'h10 ;
			data[25504] <= 8'h10 ;
			data[25505] <= 8'h10 ;
			data[25506] <= 8'h10 ;
			data[25507] <= 8'h10 ;
			data[25508] <= 8'h10 ;
			data[25509] <= 8'h10 ;
			data[25510] <= 8'h10 ;
			data[25511] <= 8'h10 ;
			data[25512] <= 8'h10 ;
			data[25513] <= 8'h10 ;
			data[25514] <= 8'h10 ;
			data[25515] <= 8'h10 ;
			data[25516] <= 8'h10 ;
			data[25517] <= 8'h10 ;
			data[25518] <= 8'h10 ;
			data[25519] <= 8'h10 ;
			data[25520] <= 8'h10 ;
			data[25521] <= 8'h10 ;
			data[25522] <= 8'h10 ;
			data[25523] <= 8'h10 ;
			data[25524] <= 8'h10 ;
			data[25525] <= 8'h10 ;
			data[25526] <= 8'h10 ;
			data[25527] <= 8'h10 ;
			data[25528] <= 8'h10 ;
			data[25529] <= 8'h10 ;
			data[25530] <= 8'h10 ;
			data[25531] <= 8'h10 ;
			data[25532] <= 8'h10 ;
			data[25533] <= 8'h10 ;
			data[25534] <= 8'h10 ;
			data[25535] <= 8'h10 ;
			data[25536] <= 8'h10 ;
			data[25537] <= 8'h10 ;
			data[25538] <= 8'h10 ;
			data[25539] <= 8'h10 ;
			data[25540] <= 8'h10 ;
			data[25541] <= 8'h10 ;
			data[25542] <= 8'h10 ;
			data[25543] <= 8'h10 ;
			data[25544] <= 8'h10 ;
			data[25545] <= 8'h10 ;
			data[25546] <= 8'h10 ;
			data[25547] <= 8'h10 ;
			data[25548] <= 8'h10 ;
			data[25549] <= 8'h10 ;
			data[25550] <= 8'h10 ;
			data[25551] <= 8'h10 ;
			data[25552] <= 8'h10 ;
			data[25553] <= 8'h10 ;
			data[25554] <= 8'h10 ;
			data[25555] <= 8'h10 ;
			data[25556] <= 8'h10 ;
			data[25557] <= 8'h10 ;
			data[25558] <= 8'h10 ;
			data[25559] <= 8'h10 ;
			data[25560] <= 8'h10 ;
			data[25561] <= 8'h10 ;
			data[25562] <= 8'h10 ;
			data[25563] <= 8'h10 ;
			data[25564] <= 8'h10 ;
			data[25565] <= 8'h10 ;
			data[25566] <= 8'h10 ;
			data[25567] <= 8'h10 ;
			data[25568] <= 8'h10 ;
			data[25569] <= 8'h10 ;
			data[25570] <= 8'h10 ;
			data[25571] <= 8'h10 ;
			data[25572] <= 8'h10 ;
			data[25573] <= 8'h10 ;
			data[25574] <= 8'h10 ;
			data[25575] <= 8'h10 ;
			data[25576] <= 8'h10 ;
			data[25577] <= 8'h10 ;
			data[25578] <= 8'h10 ;
			data[25579] <= 8'h10 ;
			data[25580] <= 8'h10 ;
			data[25581] <= 8'h10 ;
			data[25582] <= 8'h10 ;
			data[25583] <= 8'h10 ;
			data[25584] <= 8'h10 ;
			data[25585] <= 8'h10 ;
			data[25586] <= 8'h10 ;
			data[25587] <= 8'h10 ;
			data[25588] <= 8'h10 ;
			data[25589] <= 8'h10 ;
			data[25590] <= 8'h10 ;
			data[25591] <= 8'h10 ;
			data[25592] <= 8'h10 ;
			data[25593] <= 8'h10 ;
			data[25594] <= 8'h10 ;
			data[25595] <= 8'h10 ;
			data[25596] <= 8'h10 ;
			data[25597] <= 8'h10 ;
			data[25598] <= 8'h10 ;
			data[25599] <= 8'h10 ;
			data[25600] <= 8'h10 ;
			data[25601] <= 8'h10 ;
			data[25602] <= 8'h10 ;
			data[25603] <= 8'h10 ;
			data[25604] <= 8'h10 ;
			data[25605] <= 8'h10 ;
			data[25606] <= 8'h10 ;
			data[25607] <= 8'h10 ;
			data[25608] <= 8'h10 ;
			data[25609] <= 8'h10 ;
			data[25610] <= 8'h10 ;
			data[25611] <= 8'h10 ;
			data[25612] <= 8'h10 ;
			data[25613] <= 8'h10 ;
			data[25614] <= 8'h10 ;
			data[25615] <= 8'h10 ;
			data[25616] <= 8'h10 ;
			data[25617] <= 8'h10 ;
			data[25618] <= 8'h10 ;
			data[25619] <= 8'h10 ;
			data[25620] <= 8'h10 ;
			data[25621] <= 8'h10 ;
			data[25622] <= 8'h10 ;
			data[25623] <= 8'h10 ;
			data[25624] <= 8'h10 ;
			data[25625] <= 8'h10 ;
			data[25626] <= 8'h10 ;
			data[25627] <= 8'h10 ;
			data[25628] <= 8'h10 ;
			data[25629] <= 8'h10 ;
			data[25630] <= 8'h10 ;
			data[25631] <= 8'h10 ;
			data[25632] <= 8'h10 ;
			data[25633] <= 8'h10 ;
			data[25634] <= 8'h10 ;
			data[25635] <= 8'h10 ;
			data[25636] <= 8'h10 ;
			data[25637] <= 8'h10 ;
			data[25638] <= 8'h10 ;
			data[25639] <= 8'h10 ;
			data[25640] <= 8'h10 ;
			data[25641] <= 8'h10 ;
			data[25642] <= 8'h10 ;
			data[25643] <= 8'h10 ;
			data[25644] <= 8'h10 ;
			data[25645] <= 8'h10 ;
			data[25646] <= 8'h10 ;
			data[25647] <= 8'h10 ;
			data[25648] <= 8'h10 ;
			data[25649] <= 8'h10 ;
			data[25650] <= 8'h10 ;
			data[25651] <= 8'h10 ;
			data[25652] <= 8'h10 ;
			data[25653] <= 8'h10 ;
			data[25654] <= 8'h10 ;
			data[25655] <= 8'h10 ;
			data[25656] <= 8'h10 ;
			data[25657] <= 8'h10 ;
			data[25658] <= 8'h10 ;
			data[25659] <= 8'h10 ;
			data[25660] <= 8'h10 ;
			data[25661] <= 8'h10 ;
			data[25662] <= 8'h10 ;
			data[25663] <= 8'h10 ;
			data[25664] <= 8'h10 ;
			data[25665] <= 8'h10 ;
			data[25666] <= 8'h10 ;
			data[25667] <= 8'h10 ;
			data[25668] <= 8'h10 ;
			data[25669] <= 8'h10 ;
			data[25670] <= 8'h10 ;
			data[25671] <= 8'h10 ;
			data[25672] <= 8'h10 ;
			data[25673] <= 8'h10 ;
			data[25674] <= 8'h10 ;
			data[25675] <= 8'h10 ;
			data[25676] <= 8'h10 ;
			data[25677] <= 8'h10 ;
			data[25678] <= 8'h10 ;
			data[25679] <= 8'h10 ;
			data[25680] <= 8'h10 ;
			data[25681] <= 8'h10 ;
			data[25682] <= 8'h10 ;
			data[25683] <= 8'h10 ;
			data[25684] <= 8'h10 ;
			data[25685] <= 8'h10 ;
			data[25686] <= 8'h10 ;
			data[25687] <= 8'h10 ;
			data[25688] <= 8'h10 ;
			data[25689] <= 8'h10 ;
			data[25690] <= 8'h10 ;
			data[25691] <= 8'h10 ;
			data[25692] <= 8'h10 ;
			data[25693] <= 8'h10 ;
			data[25694] <= 8'h10 ;
			data[25695] <= 8'h10 ;
			data[25696] <= 8'h10 ;
			data[25697] <= 8'h10 ;
			data[25698] <= 8'h10 ;
			data[25699] <= 8'h10 ;
			data[25700] <= 8'h10 ;
			data[25701] <= 8'h10 ;
			data[25702] <= 8'h10 ;
			data[25703] <= 8'h10 ;
			data[25704] <= 8'h10 ;
			data[25705] <= 8'h10 ;
			data[25706] <= 8'h10 ;
			data[25707] <= 8'h10 ;
			data[25708] <= 8'h10 ;
			data[25709] <= 8'h10 ;
			data[25710] <= 8'h10 ;
			data[25711] <= 8'h10 ;
			data[25712] <= 8'h10 ;
			data[25713] <= 8'h10 ;
			data[25714] <= 8'h10 ;
			data[25715] <= 8'h10 ;
			data[25716] <= 8'h10 ;
			data[25717] <= 8'h10 ;
			data[25718] <= 8'h10 ;
			data[25719] <= 8'h10 ;
			data[25720] <= 8'h10 ;
			data[25721] <= 8'h10 ;
			data[25722] <= 8'h10 ;
			data[25723] <= 8'h10 ;
			data[25724] <= 8'h10 ;
			data[25725] <= 8'h10 ;
			data[25726] <= 8'h10 ;
			data[25727] <= 8'h10 ;
			data[25728] <= 8'h10 ;
			data[25729] <= 8'h10 ;
			data[25730] <= 8'h10 ;
			data[25731] <= 8'h10 ;
			data[25732] <= 8'h10 ;
			data[25733] <= 8'h10 ;
			data[25734] <= 8'h10 ;
			data[25735] <= 8'h10 ;
			data[25736] <= 8'h10 ;
			data[25737] <= 8'h10 ;
			data[25738] <= 8'h10 ;
			data[25739] <= 8'h10 ;
			data[25740] <= 8'h10 ;
			data[25741] <= 8'h10 ;
			data[25742] <= 8'h10 ;
			data[25743] <= 8'h10 ;
			data[25744] <= 8'h10 ;
			data[25745] <= 8'h10 ;
			data[25746] <= 8'h10 ;
			data[25747] <= 8'h10 ;
			data[25748] <= 8'h10 ;
			data[25749] <= 8'h10 ;
			data[25750] <= 8'h10 ;
			data[25751] <= 8'h10 ;
			data[25752] <= 8'h10 ;
			data[25753] <= 8'h10 ;
			data[25754] <= 8'h10 ;
			data[25755] <= 8'h10 ;
			data[25756] <= 8'h10 ;
			data[25757] <= 8'h10 ;
			data[25758] <= 8'h10 ;
			data[25759] <= 8'h10 ;
			data[25760] <= 8'h10 ;
			data[25761] <= 8'h10 ;
			data[25762] <= 8'h10 ;
			data[25763] <= 8'h10 ;
			data[25764] <= 8'h10 ;
			data[25765] <= 8'h10 ;
			data[25766] <= 8'h10 ;
			data[25767] <= 8'h10 ;
			data[25768] <= 8'h10 ;
			data[25769] <= 8'h10 ;
			data[25770] <= 8'h10 ;
			data[25771] <= 8'h10 ;
			data[25772] <= 8'h10 ;
			data[25773] <= 8'h10 ;
			data[25774] <= 8'h10 ;
			data[25775] <= 8'h10 ;
			data[25776] <= 8'h10 ;
			data[25777] <= 8'h10 ;
			data[25778] <= 8'h10 ;
			data[25779] <= 8'h10 ;
			data[25780] <= 8'h10 ;
			data[25781] <= 8'h10 ;
			data[25782] <= 8'h10 ;
			data[25783] <= 8'h10 ;
			data[25784] <= 8'h10 ;
			data[25785] <= 8'h10 ;
			data[25786] <= 8'h10 ;
			data[25787] <= 8'h10 ;
			data[25788] <= 8'h10 ;
			data[25789] <= 8'h10 ;
			data[25790] <= 8'h10 ;
			data[25791] <= 8'h10 ;
			data[25792] <= 8'h10 ;
			data[25793] <= 8'h10 ;
			data[25794] <= 8'h10 ;
			data[25795] <= 8'h10 ;
			data[25796] <= 8'h10 ;
			data[25797] <= 8'h10 ;
			data[25798] <= 8'h10 ;
			data[25799] <= 8'h10 ;
			data[25800] <= 8'h10 ;
			data[25801] <= 8'h10 ;
			data[25802] <= 8'h10 ;
			data[25803] <= 8'h10 ;
			data[25804] <= 8'h10 ;
			data[25805] <= 8'h10 ;
			data[25806] <= 8'h10 ;
			data[25807] <= 8'h10 ;
			data[25808] <= 8'h10 ;
			data[25809] <= 8'h10 ;
			data[25810] <= 8'h10 ;
			data[25811] <= 8'h10 ;
			data[25812] <= 8'h10 ;
			data[25813] <= 8'h10 ;
			data[25814] <= 8'h10 ;
			data[25815] <= 8'h10 ;
			data[25816] <= 8'h10 ;
			data[25817] <= 8'h10 ;
			data[25818] <= 8'h10 ;
			data[25819] <= 8'h10 ;
			data[25820] <= 8'h10 ;
			data[25821] <= 8'h10 ;
			data[25822] <= 8'h10 ;
			data[25823] <= 8'h10 ;
			data[25824] <= 8'h10 ;
			data[25825] <= 8'h10 ;
			data[25826] <= 8'h10 ;
			data[25827] <= 8'h10 ;
			data[25828] <= 8'h10 ;
			data[25829] <= 8'h10 ;
			data[25830] <= 8'h10 ;
			data[25831] <= 8'h10 ;
			data[25832] <= 8'h10 ;
			data[25833] <= 8'h10 ;
			data[25834] <= 8'h10 ;
			data[25835] <= 8'h10 ;
			data[25836] <= 8'h10 ;
			data[25837] <= 8'h10 ;
			data[25838] <= 8'h10 ;
			data[25839] <= 8'h10 ;
			data[25840] <= 8'h10 ;
			data[25841] <= 8'h10 ;
			data[25842] <= 8'h10 ;
			data[25843] <= 8'h10 ;
			data[25844] <= 8'h10 ;
			data[25845] <= 8'h10 ;
			data[25846] <= 8'h10 ;
			data[25847] <= 8'h10 ;
			data[25848] <= 8'h10 ;
			data[25849] <= 8'h10 ;
			data[25850] <= 8'h10 ;
			data[25851] <= 8'h10 ;
			data[25852] <= 8'h10 ;
			data[25853] <= 8'h10 ;
			data[25854] <= 8'h10 ;
			data[25855] <= 8'h10 ;
			data[25856] <= 8'h10 ;
			data[25857] <= 8'h10 ;
			data[25858] <= 8'h10 ;
			data[25859] <= 8'h10 ;
			data[25860] <= 8'h10 ;
			data[25861] <= 8'h10 ;
			data[25862] <= 8'h10 ;
			data[25863] <= 8'h10 ;
			data[25864] <= 8'h10 ;
			data[25865] <= 8'h10 ;
			data[25866] <= 8'h10 ;
			data[25867] <= 8'h10 ;
			data[25868] <= 8'h10 ;
			data[25869] <= 8'h10 ;
			data[25870] <= 8'h10 ;
			data[25871] <= 8'h10 ;
			data[25872] <= 8'h10 ;
			data[25873] <= 8'h10 ;
			data[25874] <= 8'h10 ;
			data[25875] <= 8'h10 ;
			data[25876] <= 8'h10 ;
			data[25877] <= 8'h10 ;
			data[25878] <= 8'h10 ;
			data[25879] <= 8'h10 ;
			data[25880] <= 8'h10 ;
			data[25881] <= 8'h10 ;
			data[25882] <= 8'h10 ;
			data[25883] <= 8'h10 ;
			data[25884] <= 8'h10 ;
			data[25885] <= 8'h10 ;
			data[25886] <= 8'h10 ;
			data[25887] <= 8'h10 ;
			data[25888] <= 8'h10 ;
			data[25889] <= 8'h10 ;
			data[25890] <= 8'h10 ;
			data[25891] <= 8'h10 ;
			data[25892] <= 8'h10 ;
			data[25893] <= 8'h10 ;
			data[25894] <= 8'h10 ;
			data[25895] <= 8'h10 ;
			data[25896] <= 8'h10 ;
			data[25897] <= 8'h10 ;
			data[25898] <= 8'h10 ;
			data[25899] <= 8'h10 ;
			data[25900] <= 8'h10 ;
			data[25901] <= 8'h10 ;
			data[25902] <= 8'h10 ;
			data[25903] <= 8'h10 ;
			data[25904] <= 8'h10 ;
			data[25905] <= 8'h10 ;
			data[25906] <= 8'h10 ;
			data[25907] <= 8'h10 ;
			data[25908] <= 8'h10 ;
			data[25909] <= 8'h10 ;
			data[25910] <= 8'h10 ;
			data[25911] <= 8'h10 ;
			data[25912] <= 8'h10 ;
			data[25913] <= 8'h10 ;
			data[25914] <= 8'h10 ;
			data[25915] <= 8'h10 ;
			data[25916] <= 8'h10 ;
			data[25917] <= 8'h10 ;
			data[25918] <= 8'h10 ;
			data[25919] <= 8'h10 ;
			data[25920] <= 8'h10 ;
			data[25921] <= 8'h10 ;
			data[25922] <= 8'h10 ;
			data[25923] <= 8'h10 ;
			data[25924] <= 8'h10 ;
			data[25925] <= 8'h10 ;
			data[25926] <= 8'h10 ;
			data[25927] <= 8'h10 ;
			data[25928] <= 8'h10 ;
			data[25929] <= 8'h10 ;
			data[25930] <= 8'h10 ;
			data[25931] <= 8'h10 ;
			data[25932] <= 8'h10 ;
			data[25933] <= 8'h10 ;
			data[25934] <= 8'h10 ;
			data[25935] <= 8'h10 ;
			data[25936] <= 8'h10 ;
			data[25937] <= 8'h10 ;
			data[25938] <= 8'h10 ;
			data[25939] <= 8'h10 ;
			data[25940] <= 8'h10 ;
			data[25941] <= 8'h10 ;
			data[25942] <= 8'h10 ;
			data[25943] <= 8'h10 ;
			data[25944] <= 8'h10 ;
			data[25945] <= 8'h10 ;
			data[25946] <= 8'h10 ;
			data[25947] <= 8'h10 ;
			data[25948] <= 8'h10 ;
			data[25949] <= 8'h10 ;
			data[25950] <= 8'h10 ;
			data[25951] <= 8'h10 ;
			data[25952] <= 8'h10 ;
			data[25953] <= 8'h10 ;
			data[25954] <= 8'h10 ;
			data[25955] <= 8'h10 ;
			data[25956] <= 8'h10 ;
			data[25957] <= 8'h10 ;
			data[25958] <= 8'h10 ;
			data[25959] <= 8'h10 ;
			data[25960] <= 8'h10 ;
			data[25961] <= 8'h10 ;
			data[25962] <= 8'h10 ;
			data[25963] <= 8'h10 ;
			data[25964] <= 8'h10 ;
			data[25965] <= 8'h10 ;
			data[25966] <= 8'h10 ;
			data[25967] <= 8'h10 ;
			data[25968] <= 8'h10 ;
			data[25969] <= 8'h10 ;
			data[25970] <= 8'h10 ;
			data[25971] <= 8'h10 ;
			data[25972] <= 8'h10 ;
			data[25973] <= 8'h10 ;
			data[25974] <= 8'h10 ;
			data[25975] <= 8'h10 ;
			data[25976] <= 8'h10 ;
			data[25977] <= 8'h10 ;
			data[25978] <= 8'h10 ;
			data[25979] <= 8'h10 ;
			data[25980] <= 8'h10 ;
			data[25981] <= 8'h10 ;
			data[25982] <= 8'h10 ;
			data[25983] <= 8'h10 ;
			data[25984] <= 8'h10 ;
			data[25985] <= 8'h10 ;
			data[25986] <= 8'h10 ;
			data[25987] <= 8'h10 ;
			data[25988] <= 8'h10 ;
			data[25989] <= 8'h10 ;
			data[25990] <= 8'h10 ;
			data[25991] <= 8'h10 ;
			data[25992] <= 8'h10 ;
			data[25993] <= 8'h10 ;
			data[25994] <= 8'h10 ;
			data[25995] <= 8'h10 ;
			data[25996] <= 8'h10 ;
			data[25997] <= 8'h10 ;
			data[25998] <= 8'h10 ;
			data[25999] <= 8'h10 ;
			data[26000] <= 8'h10 ;
			data[26001] <= 8'h10 ;
			data[26002] <= 8'h10 ;
			data[26003] <= 8'h10 ;
			data[26004] <= 8'h10 ;
			data[26005] <= 8'h10 ;
			data[26006] <= 8'h10 ;
			data[26007] <= 8'h10 ;
			data[26008] <= 8'h10 ;
			data[26009] <= 8'h10 ;
			data[26010] <= 8'h10 ;
			data[26011] <= 8'h10 ;
			data[26012] <= 8'h10 ;
			data[26013] <= 8'h10 ;
			data[26014] <= 8'h10 ;
			data[26015] <= 8'h10 ;
			data[26016] <= 8'h10 ;
			data[26017] <= 8'h10 ;
			data[26018] <= 8'h10 ;
			data[26019] <= 8'h10 ;
			data[26020] <= 8'h10 ;
			data[26021] <= 8'h10 ;
			data[26022] <= 8'h10 ;
			data[26023] <= 8'h10 ;
			data[26024] <= 8'h10 ;
			data[26025] <= 8'h10 ;
			data[26026] <= 8'h10 ;
			data[26027] <= 8'h10 ;
			data[26028] <= 8'h10 ;
			data[26029] <= 8'h10 ;
			data[26030] <= 8'h10 ;
			data[26031] <= 8'h10 ;
			data[26032] <= 8'h10 ;
			data[26033] <= 8'h10 ;
			data[26034] <= 8'h10 ;
			data[26035] <= 8'h10 ;
			data[26036] <= 8'h10 ;
			data[26037] <= 8'h10 ;
			data[26038] <= 8'h10 ;
			data[26039] <= 8'h10 ;
			data[26040] <= 8'h10 ;
			data[26041] <= 8'h10 ;
			data[26042] <= 8'h10 ;
			data[26043] <= 8'h10 ;
			data[26044] <= 8'h10 ;
			data[26045] <= 8'h10 ;
			data[26046] <= 8'h10 ;
			data[26047] <= 8'h10 ;
			data[26048] <= 8'h10 ;
			data[26049] <= 8'h10 ;
			data[26050] <= 8'h10 ;
			data[26051] <= 8'h10 ;
			data[26052] <= 8'h10 ;
			data[26053] <= 8'h10 ;
			data[26054] <= 8'h10 ;
			data[26055] <= 8'h10 ;
			data[26056] <= 8'h10 ;
			data[26057] <= 8'h10 ;
			data[26058] <= 8'h10 ;
			data[26059] <= 8'h10 ;
			data[26060] <= 8'h10 ;
			data[26061] <= 8'h10 ;
			data[26062] <= 8'h10 ;
			data[26063] <= 8'h10 ;
			data[26064] <= 8'h10 ;
			data[26065] <= 8'h10 ;
			data[26066] <= 8'h10 ;
			data[26067] <= 8'h10 ;
			data[26068] <= 8'h10 ;
			data[26069] <= 8'h10 ;
			data[26070] <= 8'h10 ;
			data[26071] <= 8'h10 ;
			data[26072] <= 8'h10 ;
			data[26073] <= 8'h10 ;
			data[26074] <= 8'h10 ;
			data[26075] <= 8'h10 ;
			data[26076] <= 8'h10 ;
			data[26077] <= 8'h10 ;
			data[26078] <= 8'h10 ;
			data[26079] <= 8'h10 ;
			data[26080] <= 8'h10 ;
			data[26081] <= 8'h10 ;
			data[26082] <= 8'h10 ;
			data[26083] <= 8'h10 ;
			data[26084] <= 8'h10 ;
			data[26085] <= 8'h10 ;
			data[26086] <= 8'h10 ;
			data[26087] <= 8'h10 ;
			data[26088] <= 8'h10 ;
			data[26089] <= 8'h10 ;
			data[26090] <= 8'h10 ;
			data[26091] <= 8'h10 ;
			data[26092] <= 8'h10 ;
			data[26093] <= 8'h10 ;
			data[26094] <= 8'h10 ;
			data[26095] <= 8'h10 ;
			data[26096] <= 8'h10 ;
			data[26097] <= 8'h10 ;
			data[26098] <= 8'h10 ;
			data[26099] <= 8'h10 ;
			data[26100] <= 8'h10 ;
			data[26101] <= 8'h10 ;
			data[26102] <= 8'h10 ;
			data[26103] <= 8'h10 ;
			data[26104] <= 8'h10 ;
			data[26105] <= 8'h10 ;
			data[26106] <= 8'h10 ;
			data[26107] <= 8'h10 ;
			data[26108] <= 8'h10 ;
			data[26109] <= 8'h10 ;
			data[26110] <= 8'h10 ;
			data[26111] <= 8'h10 ;
			data[26112] <= 8'h10 ;
			data[26113] <= 8'h10 ;
			data[26114] <= 8'h10 ;
			data[26115] <= 8'h10 ;
			data[26116] <= 8'h10 ;
			data[26117] <= 8'h10 ;
			data[26118] <= 8'h10 ;
			data[26119] <= 8'h10 ;
			data[26120] <= 8'h10 ;
			data[26121] <= 8'h10 ;
			data[26122] <= 8'h10 ;
			data[26123] <= 8'h10 ;
			data[26124] <= 8'h10 ;
			data[26125] <= 8'h10 ;
			data[26126] <= 8'h10 ;
			data[26127] <= 8'h10 ;
			data[26128] <= 8'h10 ;
			data[26129] <= 8'h10 ;
			data[26130] <= 8'h10 ;
			data[26131] <= 8'h10 ;
			data[26132] <= 8'h10 ;
			data[26133] <= 8'h10 ;
			data[26134] <= 8'h10 ;
			data[26135] <= 8'h10 ;
			data[26136] <= 8'h10 ;
			data[26137] <= 8'h10 ;
			data[26138] <= 8'h10 ;
			data[26139] <= 8'h10 ;
			data[26140] <= 8'h10 ;
			data[26141] <= 8'h10 ;
			data[26142] <= 8'h10 ;
			data[26143] <= 8'h10 ;
			data[26144] <= 8'h10 ;
			data[26145] <= 8'h10 ;
			data[26146] <= 8'h10 ;
			data[26147] <= 8'h10 ;
			data[26148] <= 8'h10 ;
			data[26149] <= 8'h10 ;
			data[26150] <= 8'h10 ;
			data[26151] <= 8'h10 ;
			data[26152] <= 8'h10 ;
			data[26153] <= 8'h10 ;
			data[26154] <= 8'h10 ;
			data[26155] <= 8'h10 ;
			data[26156] <= 8'h10 ;
			data[26157] <= 8'h10 ;
			data[26158] <= 8'h10 ;
			data[26159] <= 8'h10 ;
			data[26160] <= 8'h10 ;
			data[26161] <= 8'h10 ;
			data[26162] <= 8'h10 ;
			data[26163] <= 8'h10 ;
			data[26164] <= 8'h10 ;
			data[26165] <= 8'h10 ;
			data[26166] <= 8'h10 ;
			data[26167] <= 8'h10 ;
			data[26168] <= 8'h10 ;
			data[26169] <= 8'h10 ;
			data[26170] <= 8'h10 ;
			data[26171] <= 8'h10 ;
			data[26172] <= 8'h10 ;
			data[26173] <= 8'h10 ;
			data[26174] <= 8'h10 ;
			data[26175] <= 8'h10 ;
			data[26176] <= 8'h10 ;
			data[26177] <= 8'h10 ;
			data[26178] <= 8'h10 ;
			data[26179] <= 8'h10 ;
			data[26180] <= 8'h10 ;
			data[26181] <= 8'h10 ;
			data[26182] <= 8'h10 ;
			data[26183] <= 8'h10 ;
			data[26184] <= 8'h10 ;
			data[26185] <= 8'h10 ;
			data[26186] <= 8'h10 ;
			data[26187] <= 8'h10 ;
			data[26188] <= 8'h10 ;
			data[26189] <= 8'h10 ;
			data[26190] <= 8'h10 ;
			data[26191] <= 8'h10 ;
			data[26192] <= 8'h10 ;
			data[26193] <= 8'h10 ;
			data[26194] <= 8'h10 ;
			data[26195] <= 8'h10 ;
			data[26196] <= 8'h10 ;
			data[26197] <= 8'h10 ;
			data[26198] <= 8'h10 ;
			data[26199] <= 8'h10 ;
			data[26200] <= 8'h10 ;
			data[26201] <= 8'h10 ;
			data[26202] <= 8'h10 ;
			data[26203] <= 8'h10 ;
			data[26204] <= 8'h10 ;
			data[26205] <= 8'h10 ;
			data[26206] <= 8'h10 ;
			data[26207] <= 8'h10 ;
			data[26208] <= 8'h10 ;
			data[26209] <= 8'h10 ;
			data[26210] <= 8'h10 ;
			data[26211] <= 8'h10 ;
			data[26212] <= 8'h10 ;
			data[26213] <= 8'h10 ;
			data[26214] <= 8'h10 ;
			data[26215] <= 8'h10 ;
			data[26216] <= 8'h10 ;
			data[26217] <= 8'h10 ;
			data[26218] <= 8'h10 ;
			data[26219] <= 8'h10 ;
			data[26220] <= 8'h10 ;
			data[26221] <= 8'h10 ;
			data[26222] <= 8'h10 ;
			data[26223] <= 8'h10 ;
			data[26224] <= 8'h10 ;
			data[26225] <= 8'h10 ;
			data[26226] <= 8'h10 ;
			data[26227] <= 8'h10 ;
			data[26228] <= 8'h10 ;
			data[26229] <= 8'h10 ;
			data[26230] <= 8'h10 ;
			data[26231] <= 8'h10 ;
			data[26232] <= 8'h10 ;
			data[26233] <= 8'h10 ;
			data[26234] <= 8'h10 ;
			data[26235] <= 8'h10 ;
			data[26236] <= 8'h10 ;
			data[26237] <= 8'h10 ;
			data[26238] <= 8'h10 ;
			data[26239] <= 8'h10 ;
			data[26240] <= 8'h10 ;
			data[26241] <= 8'h10 ;
			data[26242] <= 8'h10 ;
			data[26243] <= 8'h10 ;
			data[26244] <= 8'h10 ;
			data[26245] <= 8'h10 ;
			data[26246] <= 8'h10 ;
			data[26247] <= 8'h10 ;
			data[26248] <= 8'h10 ;
			data[26249] <= 8'h10 ;
			data[26250] <= 8'h10 ;
			data[26251] <= 8'h10 ;
			data[26252] <= 8'h10 ;
			data[26253] <= 8'h10 ;
			data[26254] <= 8'h10 ;
			data[26255] <= 8'h10 ;
			data[26256] <= 8'h10 ;
			data[26257] <= 8'h10 ;
			data[26258] <= 8'h10 ;
			data[26259] <= 8'h10 ;
			data[26260] <= 8'h10 ;
			data[26261] <= 8'h10 ;
			data[26262] <= 8'h10 ;
			data[26263] <= 8'h10 ;
			data[26264] <= 8'h10 ;
			data[26265] <= 8'h10 ;
			data[26266] <= 8'h10 ;
			data[26267] <= 8'h10 ;
			data[26268] <= 8'h10 ;
			data[26269] <= 8'h10 ;
			data[26270] <= 8'h10 ;
			data[26271] <= 8'h10 ;
			data[26272] <= 8'h10 ;
			data[26273] <= 8'h10 ;
			data[26274] <= 8'h10 ;
			data[26275] <= 8'h10 ;
			data[26276] <= 8'h10 ;
			data[26277] <= 8'h10 ;
			data[26278] <= 8'h10 ;
			data[26279] <= 8'h10 ;
			data[26280] <= 8'h10 ;
			data[26281] <= 8'h10 ;
			data[26282] <= 8'h10 ;
			data[26283] <= 8'h10 ;
			data[26284] <= 8'h10 ;
			data[26285] <= 8'h10 ;
			data[26286] <= 8'h10 ;
			data[26287] <= 8'h10 ;
			data[26288] <= 8'h10 ;
			data[26289] <= 8'h10 ;
			data[26290] <= 8'h10 ;
			data[26291] <= 8'h10 ;
			data[26292] <= 8'h10 ;
			data[26293] <= 8'h10 ;
			data[26294] <= 8'h10 ;
			data[26295] <= 8'h10 ;
			data[26296] <= 8'h10 ;
			data[26297] <= 8'h10 ;
			data[26298] <= 8'h10 ;
			data[26299] <= 8'h10 ;
			data[26300] <= 8'h10 ;
			data[26301] <= 8'h10 ;
			data[26302] <= 8'h10 ;
			data[26303] <= 8'h10 ;
			data[26304] <= 8'h10 ;
			data[26305] <= 8'h10 ;
			data[26306] <= 8'h10 ;
			data[26307] <= 8'h10 ;
			data[26308] <= 8'h10 ;
			data[26309] <= 8'h10 ;
			data[26310] <= 8'h10 ;
			data[26311] <= 8'h10 ;
			data[26312] <= 8'h10 ;
			data[26313] <= 8'h10 ;
			data[26314] <= 8'h10 ;
			data[26315] <= 8'h10 ;
			data[26316] <= 8'h10 ;
			data[26317] <= 8'h10 ;
			data[26318] <= 8'h10 ;
			data[26319] <= 8'h10 ;
			data[26320] <= 8'h10 ;
			data[26321] <= 8'h10 ;
			data[26322] <= 8'h10 ;
			data[26323] <= 8'h10 ;
			data[26324] <= 8'h10 ;
			data[26325] <= 8'h10 ;
			data[26326] <= 8'h10 ;
			data[26327] <= 8'h10 ;
			data[26328] <= 8'h10 ;
			data[26329] <= 8'h10 ;
			data[26330] <= 8'h10 ;
			data[26331] <= 8'h10 ;
			data[26332] <= 8'h10 ;
			data[26333] <= 8'h10 ;
			data[26334] <= 8'h10 ;
			data[26335] <= 8'h10 ;
			data[26336] <= 8'h10 ;
			data[26337] <= 8'h10 ;
			data[26338] <= 8'h10 ;
			data[26339] <= 8'h10 ;
			data[26340] <= 8'h10 ;
			data[26341] <= 8'h10 ;
			data[26342] <= 8'h10 ;
			data[26343] <= 8'h10 ;
			data[26344] <= 8'h10 ;
			data[26345] <= 8'h10 ;
			data[26346] <= 8'h10 ;
			data[26347] <= 8'h10 ;
			data[26348] <= 8'h10 ;
			data[26349] <= 8'h10 ;
			data[26350] <= 8'h10 ;
			data[26351] <= 8'h10 ;
			data[26352] <= 8'h10 ;
			data[26353] <= 8'h10 ;
			data[26354] <= 8'h10 ;
			data[26355] <= 8'h10 ;
			data[26356] <= 8'h10 ;
			data[26357] <= 8'h10 ;
			data[26358] <= 8'h10 ;
			data[26359] <= 8'h10 ;
			data[26360] <= 8'h10 ;
			data[26361] <= 8'h10 ;
			data[26362] <= 8'h10 ;
			data[26363] <= 8'h10 ;
			data[26364] <= 8'h10 ;
			data[26365] <= 8'h10 ;
			data[26366] <= 8'h10 ;
			data[26367] <= 8'h10 ;
			data[26368] <= 8'h10 ;
			data[26369] <= 8'h10 ;
			data[26370] <= 8'h10 ;
			data[26371] <= 8'h10 ;
			data[26372] <= 8'h10 ;
			data[26373] <= 8'h10 ;
			data[26374] <= 8'h10 ;
			data[26375] <= 8'h10 ;
			data[26376] <= 8'h10 ;
			data[26377] <= 8'h10 ;
			data[26378] <= 8'h10 ;
			data[26379] <= 8'h10 ;
			data[26380] <= 8'h10 ;
			data[26381] <= 8'h10 ;
			data[26382] <= 8'h10 ;
			data[26383] <= 8'h10 ;
			data[26384] <= 8'h10 ;
			data[26385] <= 8'h10 ;
			data[26386] <= 8'h10 ;
			data[26387] <= 8'h10 ;
			data[26388] <= 8'h10 ;
			data[26389] <= 8'h10 ;
			data[26390] <= 8'h10 ;
			data[26391] <= 8'h10 ;
			data[26392] <= 8'h10 ;
			data[26393] <= 8'h10 ;
			data[26394] <= 8'h10 ;
			data[26395] <= 8'h10 ;
			data[26396] <= 8'h10 ;
			data[26397] <= 8'h10 ;
			data[26398] <= 8'h10 ;
			data[26399] <= 8'h10 ;
			data[26400] <= 8'h10 ;
			data[26401] <= 8'h10 ;
			data[26402] <= 8'h10 ;
			data[26403] <= 8'h10 ;
			data[26404] <= 8'h10 ;
			data[26405] <= 8'h10 ;
			data[26406] <= 8'h10 ;
			data[26407] <= 8'h10 ;
			data[26408] <= 8'h10 ;
			data[26409] <= 8'h10 ;
			data[26410] <= 8'h10 ;
			data[26411] <= 8'h10 ;
			data[26412] <= 8'h10 ;
			data[26413] <= 8'h10 ;
			data[26414] <= 8'h10 ;
			data[26415] <= 8'h10 ;
			data[26416] <= 8'h10 ;
			data[26417] <= 8'h10 ;
			data[26418] <= 8'h10 ;
			data[26419] <= 8'h10 ;
			data[26420] <= 8'h10 ;
			data[26421] <= 8'h10 ;
			data[26422] <= 8'h10 ;
			data[26423] <= 8'h10 ;
			data[26424] <= 8'h10 ;
			data[26425] <= 8'h10 ;
			data[26426] <= 8'h10 ;
			data[26427] <= 8'h10 ;
			data[26428] <= 8'h10 ;
			data[26429] <= 8'h10 ;
			data[26430] <= 8'h10 ;
			data[26431] <= 8'h10 ;
			data[26432] <= 8'h10 ;
			data[26433] <= 8'h10 ;
			data[26434] <= 8'h10 ;
			data[26435] <= 8'h10 ;
			data[26436] <= 8'h10 ;
			data[26437] <= 8'h10 ;
			data[26438] <= 8'h10 ;
			data[26439] <= 8'h10 ;
			data[26440] <= 8'h10 ;
			data[26441] <= 8'h10 ;
			data[26442] <= 8'h10 ;
			data[26443] <= 8'h10 ;
			data[26444] <= 8'h10 ;
			data[26445] <= 8'h10 ;
			data[26446] <= 8'h10 ;
			data[26447] <= 8'h10 ;
			data[26448] <= 8'h10 ;
			data[26449] <= 8'h10 ;
			data[26450] <= 8'h10 ;
			data[26451] <= 8'h10 ;
			data[26452] <= 8'h10 ;
			data[26453] <= 8'h10 ;
			data[26454] <= 8'h10 ;
			data[26455] <= 8'h10 ;
			data[26456] <= 8'h10 ;
			data[26457] <= 8'h10 ;
			data[26458] <= 8'h10 ;
			data[26459] <= 8'h10 ;
			data[26460] <= 8'h10 ;
			data[26461] <= 8'h10 ;
			data[26462] <= 8'h10 ;
			data[26463] <= 8'h10 ;
			data[26464] <= 8'h10 ;
			data[26465] <= 8'h10 ;
			data[26466] <= 8'h10 ;
			data[26467] <= 8'h10 ;
			data[26468] <= 8'h10 ;
			data[26469] <= 8'h10 ;
			data[26470] <= 8'h10 ;
			data[26471] <= 8'h10 ;
			data[26472] <= 8'h10 ;
			data[26473] <= 8'h10 ;
			data[26474] <= 8'h10 ;
			data[26475] <= 8'h10 ;
			data[26476] <= 8'h10 ;
			data[26477] <= 8'h10 ;
			data[26478] <= 8'h10 ;
			data[26479] <= 8'h10 ;
			data[26480] <= 8'h10 ;
			data[26481] <= 8'h10 ;
			data[26482] <= 8'h10 ;
			data[26483] <= 8'h10 ;
			data[26484] <= 8'h10 ;
			data[26485] <= 8'h10 ;
			data[26486] <= 8'h10 ;
			data[26487] <= 8'h10 ;
			data[26488] <= 8'h10 ;
			data[26489] <= 8'h10 ;
			data[26490] <= 8'h10 ;
			data[26491] <= 8'h10 ;
			data[26492] <= 8'h10 ;
			data[26493] <= 8'h10 ;
			data[26494] <= 8'h10 ;
			data[26495] <= 8'h10 ;
			data[26496] <= 8'h10 ;
			data[26497] <= 8'h10 ;
			data[26498] <= 8'h10 ;
			data[26499] <= 8'h10 ;
			data[26500] <= 8'h10 ;
			data[26501] <= 8'h10 ;
			data[26502] <= 8'h10 ;
			data[26503] <= 8'h10 ;
			data[26504] <= 8'h10 ;
			data[26505] <= 8'h10 ;
			data[26506] <= 8'h10 ;
			data[26507] <= 8'h10 ;
			data[26508] <= 8'h10 ;
			data[26509] <= 8'h10 ;
			data[26510] <= 8'h10 ;
			data[26511] <= 8'h10 ;
			data[26512] <= 8'h10 ;
			data[26513] <= 8'h10 ;
			data[26514] <= 8'h10 ;
			data[26515] <= 8'h10 ;
			data[26516] <= 8'h10 ;
			data[26517] <= 8'h10 ;
			data[26518] <= 8'h10 ;
			data[26519] <= 8'h10 ;
			data[26520] <= 8'h10 ;
			data[26521] <= 8'h10 ;
			data[26522] <= 8'h10 ;
			data[26523] <= 8'h10 ;
			data[26524] <= 8'h10 ;
			data[26525] <= 8'h10 ;
			data[26526] <= 8'h10 ;
			data[26527] <= 8'h10 ;
			data[26528] <= 8'h10 ;
			data[26529] <= 8'h10 ;
			data[26530] <= 8'h10 ;
			data[26531] <= 8'h10 ;
			data[26532] <= 8'h10 ;
			data[26533] <= 8'h10 ;
			data[26534] <= 8'h10 ;
			data[26535] <= 8'h10 ;
			data[26536] <= 8'h10 ;
			data[26537] <= 8'h10 ;
			data[26538] <= 8'h10 ;
			data[26539] <= 8'h10 ;
			data[26540] <= 8'h10 ;
			data[26541] <= 8'h10 ;
			data[26542] <= 8'h10 ;
			data[26543] <= 8'h10 ;
			data[26544] <= 8'h10 ;
			data[26545] <= 8'h10 ;
			data[26546] <= 8'h10 ;
			data[26547] <= 8'h10 ;
			data[26548] <= 8'h10 ;
			data[26549] <= 8'h10 ;
			data[26550] <= 8'h10 ;
			data[26551] <= 8'h10 ;
			data[26552] <= 8'h10 ;
			data[26553] <= 8'h10 ;
			data[26554] <= 8'h10 ;
			data[26555] <= 8'h10 ;
			data[26556] <= 8'h10 ;
			data[26557] <= 8'h10 ;
			data[26558] <= 8'h10 ;
			data[26559] <= 8'h10 ;
			data[26560] <= 8'h10 ;
			data[26561] <= 8'h10 ;
			data[26562] <= 8'h10 ;
			data[26563] <= 8'h10 ;
			data[26564] <= 8'h10 ;
			data[26565] <= 8'h10 ;
			data[26566] <= 8'h10 ;
			data[26567] <= 8'h10 ;
			data[26568] <= 8'h10 ;
			data[26569] <= 8'h10 ;
			data[26570] <= 8'h10 ;
			data[26571] <= 8'h10 ;
			data[26572] <= 8'h10 ;
			data[26573] <= 8'h10 ;
			data[26574] <= 8'h10 ;
			data[26575] <= 8'h10 ;
			data[26576] <= 8'h10 ;
			data[26577] <= 8'h10 ;
			data[26578] <= 8'h10 ;
			data[26579] <= 8'h10 ;
			data[26580] <= 8'h10 ;
			data[26581] <= 8'h10 ;
			data[26582] <= 8'h10 ;
			data[26583] <= 8'h10 ;
			data[26584] <= 8'h10 ;
			data[26585] <= 8'h10 ;
			data[26586] <= 8'h10 ;
			data[26587] <= 8'h10 ;
			data[26588] <= 8'h10 ;
			data[26589] <= 8'h10 ;
			data[26590] <= 8'h10 ;
			data[26591] <= 8'h10 ;
			data[26592] <= 8'h10 ;
			data[26593] <= 8'h10 ;
			data[26594] <= 8'h10 ;
			data[26595] <= 8'h10 ;
			data[26596] <= 8'h10 ;
			data[26597] <= 8'h10 ;
			data[26598] <= 8'h10 ;
			data[26599] <= 8'h10 ;
			data[26600] <= 8'h10 ;
			data[26601] <= 8'h10 ;
			data[26602] <= 8'h10 ;
			data[26603] <= 8'h10 ;
			data[26604] <= 8'h10 ;
			data[26605] <= 8'h10 ;
			data[26606] <= 8'h10 ;
			data[26607] <= 8'h10 ;
			data[26608] <= 8'h10 ;
			data[26609] <= 8'h10 ;
			data[26610] <= 8'h10 ;
			data[26611] <= 8'h10 ;
			data[26612] <= 8'h10 ;
			data[26613] <= 8'h10 ;
			data[26614] <= 8'h10 ;
			data[26615] <= 8'h10 ;
			data[26616] <= 8'h10 ;
			data[26617] <= 8'h10 ;
			data[26618] <= 8'h10 ;
			data[26619] <= 8'h10 ;
			data[26620] <= 8'h10 ;
			data[26621] <= 8'h10 ;
			data[26622] <= 8'h10 ;
			data[26623] <= 8'h10 ;
			data[26624] <= 8'h10 ;
			data[26625] <= 8'h10 ;
			data[26626] <= 8'h10 ;
			data[26627] <= 8'h10 ;
			data[26628] <= 8'h10 ;
			data[26629] <= 8'h10 ;
			data[26630] <= 8'h10 ;
			data[26631] <= 8'h10 ;
			data[26632] <= 8'h10 ;
			data[26633] <= 8'h10 ;
			data[26634] <= 8'h10 ;
			data[26635] <= 8'h10 ;
			data[26636] <= 8'h10 ;
			data[26637] <= 8'h10 ;
			data[26638] <= 8'h10 ;
			data[26639] <= 8'h10 ;
			data[26640] <= 8'h10 ;
			data[26641] <= 8'h10 ;
			data[26642] <= 8'h10 ;
			data[26643] <= 8'h10 ;
			data[26644] <= 8'h10 ;
			data[26645] <= 8'h10 ;
			data[26646] <= 8'h10 ;
			data[26647] <= 8'h10 ;
			data[26648] <= 8'h10 ;
			data[26649] <= 8'h10 ;
			data[26650] <= 8'h10 ;
			data[26651] <= 8'h10 ;
			data[26652] <= 8'h10 ;
			data[26653] <= 8'h10 ;
			data[26654] <= 8'h10 ;
			data[26655] <= 8'h10 ;
			data[26656] <= 8'h10 ;
			data[26657] <= 8'h10 ;
			data[26658] <= 8'h10 ;
			data[26659] <= 8'h10 ;
			data[26660] <= 8'h10 ;
			data[26661] <= 8'h10 ;
			data[26662] <= 8'h10 ;
			data[26663] <= 8'h10 ;
			data[26664] <= 8'h10 ;
			data[26665] <= 8'h10 ;
			data[26666] <= 8'h10 ;
			data[26667] <= 8'h10 ;
			data[26668] <= 8'h10 ;
			data[26669] <= 8'h10 ;
			data[26670] <= 8'h10 ;
			data[26671] <= 8'h10 ;
			data[26672] <= 8'h10 ;
			data[26673] <= 8'h10 ;
			data[26674] <= 8'h10 ;
			data[26675] <= 8'h10 ;
			data[26676] <= 8'h10 ;
			data[26677] <= 8'h10 ;
			data[26678] <= 8'h10 ;
			data[26679] <= 8'h10 ;
			data[26680] <= 8'h10 ;
			data[26681] <= 8'h10 ;
			data[26682] <= 8'h10 ;
			data[26683] <= 8'h10 ;
			data[26684] <= 8'h10 ;
			data[26685] <= 8'h10 ;
			data[26686] <= 8'h10 ;
			data[26687] <= 8'h10 ;
			data[26688] <= 8'h10 ;
			data[26689] <= 8'h10 ;
			data[26690] <= 8'h10 ;
			data[26691] <= 8'h10 ;
			data[26692] <= 8'h10 ;
			data[26693] <= 8'h10 ;
			data[26694] <= 8'h10 ;
			data[26695] <= 8'h10 ;
			data[26696] <= 8'h10 ;
			data[26697] <= 8'h10 ;
			data[26698] <= 8'h10 ;
			data[26699] <= 8'h10 ;
			data[26700] <= 8'h10 ;
			data[26701] <= 8'h10 ;
			data[26702] <= 8'h10 ;
			data[26703] <= 8'h10 ;
			data[26704] <= 8'h10 ;
			data[26705] <= 8'h10 ;
			data[26706] <= 8'h10 ;
			data[26707] <= 8'h10 ;
			data[26708] <= 8'h10 ;
			data[26709] <= 8'h10 ;
			data[26710] <= 8'h10 ;
			data[26711] <= 8'h10 ;
			data[26712] <= 8'h10 ;
			data[26713] <= 8'h10 ;
			data[26714] <= 8'h10 ;
			data[26715] <= 8'h10 ;
			data[26716] <= 8'h10 ;
			data[26717] <= 8'h10 ;
			data[26718] <= 8'h10 ;
			data[26719] <= 8'h10 ;
			data[26720] <= 8'h10 ;
			data[26721] <= 8'h10 ;
			data[26722] <= 8'h10 ;
			data[26723] <= 8'h10 ;
			data[26724] <= 8'h10 ;
			data[26725] <= 8'h10 ;
			data[26726] <= 8'h10 ;
			data[26727] <= 8'h10 ;
			data[26728] <= 8'h10 ;
			data[26729] <= 8'h10 ;
			data[26730] <= 8'h10 ;
			data[26731] <= 8'h10 ;
			data[26732] <= 8'h10 ;
			data[26733] <= 8'h10 ;
			data[26734] <= 8'h10 ;
			data[26735] <= 8'h10 ;
			data[26736] <= 8'h10 ;
			data[26737] <= 8'h10 ;
			data[26738] <= 8'h10 ;
			data[26739] <= 8'h10 ;
			data[26740] <= 8'h10 ;
			data[26741] <= 8'h10 ;
			data[26742] <= 8'h10 ;
			data[26743] <= 8'h10 ;
			data[26744] <= 8'h10 ;
			data[26745] <= 8'h10 ;
			data[26746] <= 8'h10 ;
			data[26747] <= 8'h10 ;
			data[26748] <= 8'h10 ;
			data[26749] <= 8'h10 ;
			data[26750] <= 8'h10 ;
			data[26751] <= 8'h10 ;
			data[26752] <= 8'h10 ;
			data[26753] <= 8'h10 ;
			data[26754] <= 8'h10 ;
			data[26755] <= 8'h10 ;
			data[26756] <= 8'h10 ;
			data[26757] <= 8'h10 ;
			data[26758] <= 8'h10 ;
			data[26759] <= 8'h10 ;
			data[26760] <= 8'h10 ;
			data[26761] <= 8'h10 ;
			data[26762] <= 8'h10 ;
			data[26763] <= 8'h10 ;
			data[26764] <= 8'h10 ;
			data[26765] <= 8'h10 ;
			data[26766] <= 8'h10 ;
			data[26767] <= 8'h10 ;
			data[26768] <= 8'h10 ;
			data[26769] <= 8'h10 ;
			data[26770] <= 8'h10 ;
			data[26771] <= 8'h10 ;
			data[26772] <= 8'h10 ;
			data[26773] <= 8'h10 ;
			data[26774] <= 8'h10 ;
			data[26775] <= 8'h10 ;
			data[26776] <= 8'h10 ;
			data[26777] <= 8'h10 ;
			data[26778] <= 8'h10 ;
			data[26779] <= 8'h10 ;
			data[26780] <= 8'h10 ;
			data[26781] <= 8'h10 ;
			data[26782] <= 8'h10 ;
			data[26783] <= 8'h10 ;
			data[26784] <= 8'h10 ;
			data[26785] <= 8'h10 ;
			data[26786] <= 8'h10 ;
			data[26787] <= 8'h10 ;
			data[26788] <= 8'h10 ;
			data[26789] <= 8'h10 ;
			data[26790] <= 8'h10 ;
			data[26791] <= 8'h10 ;
			data[26792] <= 8'h10 ;
			data[26793] <= 8'h10 ;
			data[26794] <= 8'h10 ;
			data[26795] <= 8'h10 ;
			data[26796] <= 8'h10 ;
			data[26797] <= 8'h10 ;
			data[26798] <= 8'h10 ;
			data[26799] <= 8'h10 ;
			data[26800] <= 8'h10 ;
			data[26801] <= 8'h10 ;
			data[26802] <= 8'h10 ;
			data[26803] <= 8'h10 ;
			data[26804] <= 8'h10 ;
			data[26805] <= 8'h10 ;
			data[26806] <= 8'h10 ;
			data[26807] <= 8'h10 ;
			data[26808] <= 8'h10 ;
			data[26809] <= 8'h10 ;
			data[26810] <= 8'h10 ;
			data[26811] <= 8'h10 ;
			data[26812] <= 8'h10 ;
			data[26813] <= 8'h10 ;
			data[26814] <= 8'h10 ;
			data[26815] <= 8'h10 ;
			data[26816] <= 8'h10 ;
			data[26817] <= 8'h10 ;
			data[26818] <= 8'h10 ;
			data[26819] <= 8'h10 ;
			data[26820] <= 8'h10 ;
			data[26821] <= 8'h10 ;
			data[26822] <= 8'h10 ;
			data[26823] <= 8'h10 ;
			data[26824] <= 8'h10 ;
			data[26825] <= 8'h10 ;
			data[26826] <= 8'h10 ;
			data[26827] <= 8'h10 ;
			data[26828] <= 8'h10 ;
			data[26829] <= 8'h10 ;
			data[26830] <= 8'h10 ;
			data[26831] <= 8'h10 ;
			data[26832] <= 8'h10 ;
			data[26833] <= 8'h10 ;
			data[26834] <= 8'h10 ;
			data[26835] <= 8'h10 ;
			data[26836] <= 8'h10 ;
			data[26837] <= 8'h10 ;
			data[26838] <= 8'h10 ;
			data[26839] <= 8'h10 ;
			data[26840] <= 8'h10 ;
			data[26841] <= 8'h10 ;
			data[26842] <= 8'h10 ;
			data[26843] <= 8'h10 ;
			data[26844] <= 8'h10 ;
			data[26845] <= 8'h10 ;
			data[26846] <= 8'h10 ;
			data[26847] <= 8'h10 ;
			data[26848] <= 8'h10 ;
			data[26849] <= 8'h10 ;
			data[26850] <= 8'h10 ;
			data[26851] <= 8'h10 ;
			data[26852] <= 8'h10 ;
			data[26853] <= 8'h10 ;
			data[26854] <= 8'h10 ;
			data[26855] <= 8'h10 ;
			data[26856] <= 8'h10 ;
			data[26857] <= 8'h10 ;
			data[26858] <= 8'h10 ;
			data[26859] <= 8'h10 ;
			data[26860] <= 8'h10 ;
			data[26861] <= 8'h10 ;
			data[26862] <= 8'h10 ;
			data[26863] <= 8'h10 ;
			data[26864] <= 8'h10 ;
			data[26865] <= 8'h10 ;
			data[26866] <= 8'h10 ;
			data[26867] <= 8'h10 ;
			data[26868] <= 8'h10 ;
			data[26869] <= 8'h10 ;
			data[26870] <= 8'h10 ;
			data[26871] <= 8'h10 ;
			data[26872] <= 8'h10 ;
			data[26873] <= 8'h10 ;
			data[26874] <= 8'h10 ;
			data[26875] <= 8'h10 ;
			data[26876] <= 8'h10 ;
			data[26877] <= 8'h10 ;
			data[26878] <= 8'h10 ;
			data[26879] <= 8'h10 ;
			data[26880] <= 8'h10 ;
			data[26881] <= 8'h10 ;
			data[26882] <= 8'h10 ;
			data[26883] <= 8'h10 ;
			data[26884] <= 8'h10 ;
			data[26885] <= 8'h10 ;
			data[26886] <= 8'h10 ;
			data[26887] <= 8'h10 ;
			data[26888] <= 8'h10 ;
			data[26889] <= 8'h10 ;
			data[26890] <= 8'h10 ;
			data[26891] <= 8'h10 ;
			data[26892] <= 8'h10 ;
			data[26893] <= 8'h10 ;
			data[26894] <= 8'h10 ;
			data[26895] <= 8'h10 ;
			data[26896] <= 8'h10 ;
			data[26897] <= 8'h10 ;
			data[26898] <= 8'h10 ;
			data[26899] <= 8'h10 ;
			data[26900] <= 8'h10 ;
			data[26901] <= 8'h10 ;
			data[26902] <= 8'h10 ;
			data[26903] <= 8'h10 ;
			data[26904] <= 8'h10 ;
			data[26905] <= 8'h10 ;
			data[26906] <= 8'h10 ;
			data[26907] <= 8'h10 ;
			data[26908] <= 8'h10 ;
			data[26909] <= 8'h10 ;
			data[26910] <= 8'h10 ;
			data[26911] <= 8'h10 ;
			data[26912] <= 8'h10 ;
			data[26913] <= 8'h10 ;
			data[26914] <= 8'h10 ;
			data[26915] <= 8'h10 ;
			data[26916] <= 8'h10 ;
			data[26917] <= 8'h10 ;
			data[26918] <= 8'h10 ;
			data[26919] <= 8'h10 ;
			data[26920] <= 8'h10 ;
			data[26921] <= 8'h10 ;
			data[26922] <= 8'h10 ;
			data[26923] <= 8'h10 ;
			data[26924] <= 8'h10 ;
			data[26925] <= 8'h10 ;
			data[26926] <= 8'h10 ;
			data[26927] <= 8'h10 ;
			data[26928] <= 8'h10 ;
			data[26929] <= 8'h10 ;
			data[26930] <= 8'h10 ;
			data[26931] <= 8'h10 ;
			data[26932] <= 8'h10 ;
			data[26933] <= 8'h10 ;
			data[26934] <= 8'h10 ;
			data[26935] <= 8'h10 ;
			data[26936] <= 8'h10 ;
			data[26937] <= 8'h10 ;
			data[26938] <= 8'h10 ;
			data[26939] <= 8'h10 ;
			data[26940] <= 8'h10 ;
			data[26941] <= 8'h10 ;
			data[26942] <= 8'h10 ;
			data[26943] <= 8'h10 ;
			data[26944] <= 8'h10 ;
			data[26945] <= 8'h10 ;
			data[26946] <= 8'h10 ;
			data[26947] <= 8'h10 ;
			data[26948] <= 8'h10 ;
			data[26949] <= 8'h10 ;
			data[26950] <= 8'h10 ;
			data[26951] <= 8'h10 ;
			data[26952] <= 8'h10 ;
			data[26953] <= 8'h10 ;
			data[26954] <= 8'h10 ;
			data[26955] <= 8'h10 ;
			data[26956] <= 8'h10 ;
			data[26957] <= 8'h10 ;
			data[26958] <= 8'h10 ;
			data[26959] <= 8'h10 ;
			data[26960] <= 8'h10 ;
			data[26961] <= 8'h10 ;
			data[26962] <= 8'h10 ;
			data[26963] <= 8'h10 ;
			data[26964] <= 8'h10 ;
			data[26965] <= 8'h10 ;
			data[26966] <= 8'h10 ;
			data[26967] <= 8'h10 ;
			data[26968] <= 8'h10 ;
			data[26969] <= 8'h10 ;
			data[26970] <= 8'h10 ;
			data[26971] <= 8'h10 ;
			data[26972] <= 8'h10 ;
			data[26973] <= 8'h10 ;
			data[26974] <= 8'h10 ;
			data[26975] <= 8'h10 ;
			data[26976] <= 8'h10 ;
			data[26977] <= 8'h10 ;
			data[26978] <= 8'h10 ;
			data[26979] <= 8'h10 ;
			data[26980] <= 8'h10 ;
			data[26981] <= 8'h10 ;
			data[26982] <= 8'h10 ;
			data[26983] <= 8'h10 ;
			data[26984] <= 8'h10 ;
			data[26985] <= 8'h10 ;
			data[26986] <= 8'h10 ;
			data[26987] <= 8'h10 ;
			data[26988] <= 8'h10 ;
			data[26989] <= 8'h10 ;
			data[26990] <= 8'h10 ;
			data[26991] <= 8'h10 ;
			data[26992] <= 8'h10 ;
			data[26993] <= 8'h10 ;
			data[26994] <= 8'h10 ;
			data[26995] <= 8'h10 ;
			data[26996] <= 8'h10 ;
			data[26997] <= 8'h10 ;
			data[26998] <= 8'h10 ;
			data[26999] <= 8'h10 ;
			data[27000] <= 8'h10 ;
			data[27001] <= 8'h10 ;
			data[27002] <= 8'h10 ;
			data[27003] <= 8'h10 ;
			data[27004] <= 8'h10 ;
			data[27005] <= 8'h10 ;
			data[27006] <= 8'h10 ;
			data[27007] <= 8'h10 ;
			data[27008] <= 8'h10 ;
			data[27009] <= 8'h10 ;
			data[27010] <= 8'h10 ;
			data[27011] <= 8'h10 ;
			data[27012] <= 8'h10 ;
			data[27013] <= 8'h10 ;
			data[27014] <= 8'h10 ;
			data[27015] <= 8'h10 ;
			data[27016] <= 8'h10 ;
			data[27017] <= 8'h10 ;
			data[27018] <= 8'h10 ;
			data[27019] <= 8'h10 ;
			data[27020] <= 8'h10 ;
			data[27021] <= 8'h10 ;
			data[27022] <= 8'h10 ;
			data[27023] <= 8'h10 ;
			data[27024] <= 8'h10 ;
			data[27025] <= 8'h10 ;
			data[27026] <= 8'h10 ;
			data[27027] <= 8'h10 ;
			data[27028] <= 8'h10 ;
			data[27029] <= 8'h10 ;
			data[27030] <= 8'h10 ;
			data[27031] <= 8'h10 ;
			data[27032] <= 8'h10 ;
			data[27033] <= 8'h10 ;
			data[27034] <= 8'h10 ;
			data[27035] <= 8'h10 ;
			data[27036] <= 8'h10 ;
			data[27037] <= 8'h10 ;
			data[27038] <= 8'h10 ;
			data[27039] <= 8'h10 ;
			data[27040] <= 8'h10 ;
			data[27041] <= 8'h10 ;
			data[27042] <= 8'h10 ;
			data[27043] <= 8'h10 ;
			data[27044] <= 8'h10 ;
			data[27045] <= 8'h10 ;
			data[27046] <= 8'h10 ;
			data[27047] <= 8'h10 ;
			data[27048] <= 8'h10 ;
			data[27049] <= 8'h10 ;
			data[27050] <= 8'h10 ;
			data[27051] <= 8'h10 ;
			data[27052] <= 8'h10 ;
			data[27053] <= 8'h10 ;
			data[27054] <= 8'h10 ;
			data[27055] <= 8'h10 ;
			data[27056] <= 8'h10 ;
			data[27057] <= 8'h10 ;
			data[27058] <= 8'h10 ;
			data[27059] <= 8'h10 ;
			data[27060] <= 8'h10 ;
			data[27061] <= 8'h10 ;
			data[27062] <= 8'h10 ;
			data[27063] <= 8'h10 ;
			data[27064] <= 8'h10 ;
			data[27065] <= 8'h10 ;
			data[27066] <= 8'h10 ;
			data[27067] <= 8'h10 ;
			data[27068] <= 8'h10 ;
			data[27069] <= 8'h10 ;
			data[27070] <= 8'h10 ;
			data[27071] <= 8'h10 ;
			data[27072] <= 8'h10 ;
			data[27073] <= 8'h10 ;
			data[27074] <= 8'h10 ;
			data[27075] <= 8'h10 ;
			data[27076] <= 8'h10 ;
			data[27077] <= 8'h10 ;
			data[27078] <= 8'h10 ;
			data[27079] <= 8'h10 ;
			data[27080] <= 8'h10 ;
			data[27081] <= 8'h10 ;
			data[27082] <= 8'h10 ;
			data[27083] <= 8'h10 ;
			data[27084] <= 8'h10 ;
			data[27085] <= 8'h10 ;
			data[27086] <= 8'h10 ;
			data[27087] <= 8'h10 ;
			data[27088] <= 8'h10 ;
			data[27089] <= 8'h10 ;
			data[27090] <= 8'h10 ;
			data[27091] <= 8'h10 ;
			data[27092] <= 8'h10 ;
			data[27093] <= 8'h10 ;
			data[27094] <= 8'h10 ;
			data[27095] <= 8'h10 ;
			data[27096] <= 8'h10 ;
			data[27097] <= 8'h10 ;
			data[27098] <= 8'h10 ;
			data[27099] <= 8'h10 ;
			data[27100] <= 8'h10 ;
			data[27101] <= 8'h10 ;
			data[27102] <= 8'h10 ;
			data[27103] <= 8'h10 ;
			data[27104] <= 8'h10 ;
			data[27105] <= 8'h10 ;
			data[27106] <= 8'h10 ;
			data[27107] <= 8'h10 ;
			data[27108] <= 8'h10 ;
			data[27109] <= 8'h10 ;
			data[27110] <= 8'h10 ;
			data[27111] <= 8'h10 ;
			data[27112] <= 8'h10 ;
			data[27113] <= 8'h10 ;
			data[27114] <= 8'h10 ;
			data[27115] <= 8'h10 ;
			data[27116] <= 8'h10 ;
			data[27117] <= 8'h10 ;
			data[27118] <= 8'h10 ;
			data[27119] <= 8'h10 ;
			data[27120] <= 8'h10 ;
			data[27121] <= 8'h10 ;
			data[27122] <= 8'h10 ;
			data[27123] <= 8'h10 ;
			data[27124] <= 8'h10 ;
			data[27125] <= 8'h10 ;
			data[27126] <= 8'h10 ;
			data[27127] <= 8'h10 ;
			data[27128] <= 8'h10 ;
			data[27129] <= 8'h10 ;
			data[27130] <= 8'h10 ;
			data[27131] <= 8'h10 ;
			data[27132] <= 8'h10 ;
			data[27133] <= 8'h10 ;
			data[27134] <= 8'h10 ;
			data[27135] <= 8'h10 ;
			data[27136] <= 8'h10 ;
			data[27137] <= 8'h10 ;
			data[27138] <= 8'h10 ;
			data[27139] <= 8'h10 ;
			data[27140] <= 8'h10 ;
			data[27141] <= 8'h10 ;
			data[27142] <= 8'h10 ;
			data[27143] <= 8'h10 ;
			data[27144] <= 8'h10 ;
			data[27145] <= 8'h10 ;
			data[27146] <= 8'h10 ;
			data[27147] <= 8'h10 ;
			data[27148] <= 8'h10 ;
			data[27149] <= 8'h10 ;
			data[27150] <= 8'h10 ;
			data[27151] <= 8'h10 ;
			data[27152] <= 8'h10 ;
			data[27153] <= 8'h10 ;
			data[27154] <= 8'h10 ;
			data[27155] <= 8'h10 ;
			data[27156] <= 8'h10 ;
			data[27157] <= 8'h10 ;
			data[27158] <= 8'h10 ;
			data[27159] <= 8'h10 ;
			data[27160] <= 8'h10 ;
			data[27161] <= 8'h10 ;
			data[27162] <= 8'h10 ;
			data[27163] <= 8'h10 ;
			data[27164] <= 8'h10 ;
			data[27165] <= 8'h10 ;
			data[27166] <= 8'h10 ;
			data[27167] <= 8'h10 ;
			data[27168] <= 8'h10 ;
			data[27169] <= 8'h10 ;
			data[27170] <= 8'h10 ;
			data[27171] <= 8'h10 ;
			data[27172] <= 8'h10 ;
			data[27173] <= 8'h10 ;
			data[27174] <= 8'h10 ;
			data[27175] <= 8'h10 ;
			data[27176] <= 8'h10 ;
			data[27177] <= 8'h10 ;
			data[27178] <= 8'h10 ;
			data[27179] <= 8'h10 ;
			data[27180] <= 8'h10 ;
			data[27181] <= 8'h10 ;
			data[27182] <= 8'h10 ;
			data[27183] <= 8'h10 ;
			data[27184] <= 8'h10 ;
			data[27185] <= 8'h10 ;
			data[27186] <= 8'h10 ;
			data[27187] <= 8'h10 ;
			data[27188] <= 8'h10 ;
			data[27189] <= 8'h10 ;
			data[27190] <= 8'h10 ;
			data[27191] <= 8'h10 ;
			data[27192] <= 8'h10 ;
			data[27193] <= 8'h10 ;
			data[27194] <= 8'h10 ;
			data[27195] <= 8'h10 ;
			data[27196] <= 8'h10 ;
			data[27197] <= 8'h10 ;
			data[27198] <= 8'h10 ;
			data[27199] <= 8'h10 ;
			data[27200] <= 8'h10 ;
			data[27201] <= 8'h10 ;
			data[27202] <= 8'h10 ;
			data[27203] <= 8'h10 ;
			data[27204] <= 8'h10 ;
			data[27205] <= 8'h10 ;
			data[27206] <= 8'h10 ;
			data[27207] <= 8'h10 ;
			data[27208] <= 8'h10 ;
			data[27209] <= 8'h10 ;
			data[27210] <= 8'h10 ;
			data[27211] <= 8'h10 ;
			data[27212] <= 8'h10 ;
			data[27213] <= 8'h10 ;
			data[27214] <= 8'h10 ;
			data[27215] <= 8'h10 ;
			data[27216] <= 8'h10 ;
			data[27217] <= 8'h10 ;
			data[27218] <= 8'h10 ;
			data[27219] <= 8'h10 ;
			data[27220] <= 8'h10 ;
			data[27221] <= 8'h10 ;
			data[27222] <= 8'h10 ;
			data[27223] <= 8'h10 ;
			data[27224] <= 8'h10 ;
			data[27225] <= 8'h10 ;
			data[27226] <= 8'h10 ;
			data[27227] <= 8'h10 ;
			data[27228] <= 8'h10 ;
			data[27229] <= 8'h10 ;
			data[27230] <= 8'h10 ;
			data[27231] <= 8'h10 ;
			data[27232] <= 8'h10 ;
			data[27233] <= 8'h10 ;
			data[27234] <= 8'h10 ;
			data[27235] <= 8'h10 ;
			data[27236] <= 8'h10 ;
			data[27237] <= 8'h10 ;
			data[27238] <= 8'h10 ;
			data[27239] <= 8'h10 ;
			data[27240] <= 8'h10 ;
			data[27241] <= 8'h10 ;
			data[27242] <= 8'h10 ;
			data[27243] <= 8'h10 ;
			data[27244] <= 8'h10 ;
			data[27245] <= 8'h10 ;
			data[27246] <= 8'h10 ;
			data[27247] <= 8'h10 ;
			data[27248] <= 8'h10 ;
			data[27249] <= 8'h10 ;
			data[27250] <= 8'h10 ;
			data[27251] <= 8'h10 ;
			data[27252] <= 8'h10 ;
			data[27253] <= 8'h10 ;
			data[27254] <= 8'h10 ;
			data[27255] <= 8'h10 ;
			data[27256] <= 8'h10 ;
			data[27257] <= 8'h10 ;
			data[27258] <= 8'h10 ;
			data[27259] <= 8'h10 ;
			data[27260] <= 8'h10 ;
			data[27261] <= 8'h10 ;
			data[27262] <= 8'h10 ;
			data[27263] <= 8'h10 ;
			data[27264] <= 8'h10 ;
			data[27265] <= 8'h10 ;
			data[27266] <= 8'h10 ;
			data[27267] <= 8'h10 ;
			data[27268] <= 8'h10 ;
			data[27269] <= 8'h10 ;
			data[27270] <= 8'h10 ;
			data[27271] <= 8'h10 ;
			data[27272] <= 8'h10 ;
			data[27273] <= 8'h10 ;
			data[27274] <= 8'h10 ;
			data[27275] <= 8'h10 ;
			data[27276] <= 8'h10 ;
			data[27277] <= 8'h10 ;
			data[27278] <= 8'h10 ;
			data[27279] <= 8'h10 ;
			data[27280] <= 8'h10 ;
			data[27281] <= 8'h10 ;
			data[27282] <= 8'h10 ;
			data[27283] <= 8'h10 ;
			data[27284] <= 8'h10 ;
			data[27285] <= 8'h10 ;
			data[27286] <= 8'h10 ;
			data[27287] <= 8'h10 ;
			data[27288] <= 8'h10 ;
			data[27289] <= 8'h10 ;
			data[27290] <= 8'h10 ;
			data[27291] <= 8'h10 ;
			data[27292] <= 8'h10 ;
			data[27293] <= 8'h10 ;
			data[27294] <= 8'h10 ;
			data[27295] <= 8'h10 ;
			data[27296] <= 8'h10 ;
			data[27297] <= 8'h10 ;
			data[27298] <= 8'h10 ;
			data[27299] <= 8'h10 ;
			data[27300] <= 8'h10 ;
			data[27301] <= 8'h10 ;
			data[27302] <= 8'h10 ;
			data[27303] <= 8'h10 ;
			data[27304] <= 8'h10 ;
			data[27305] <= 8'h10 ;
			data[27306] <= 8'h10 ;
			data[27307] <= 8'h10 ;
			data[27308] <= 8'h10 ;
			data[27309] <= 8'h10 ;
			data[27310] <= 8'h10 ;
			data[27311] <= 8'h10 ;
			data[27312] <= 8'h10 ;
			data[27313] <= 8'h10 ;
			data[27314] <= 8'h10 ;
			data[27315] <= 8'h10 ;
			data[27316] <= 8'h10 ;
			data[27317] <= 8'h10 ;
			data[27318] <= 8'h10 ;
			data[27319] <= 8'h10 ;
			data[27320] <= 8'h10 ;
			data[27321] <= 8'h10 ;
			data[27322] <= 8'h10 ;
			data[27323] <= 8'h10 ;
			data[27324] <= 8'h10 ;
			data[27325] <= 8'h10 ;
			data[27326] <= 8'h10 ;
			data[27327] <= 8'h10 ;
			data[27328] <= 8'h10 ;
			data[27329] <= 8'h10 ;
			data[27330] <= 8'h10 ;
			data[27331] <= 8'h10 ;
			data[27332] <= 8'h10 ;
			data[27333] <= 8'h10 ;
			data[27334] <= 8'h10 ;
			data[27335] <= 8'h10 ;
			data[27336] <= 8'h10 ;
			data[27337] <= 8'h10 ;
			data[27338] <= 8'h10 ;
			data[27339] <= 8'h10 ;
			data[27340] <= 8'h10 ;
			data[27341] <= 8'h10 ;
			data[27342] <= 8'h10 ;
			data[27343] <= 8'h10 ;
			data[27344] <= 8'h10 ;
			data[27345] <= 8'h10 ;
			data[27346] <= 8'h10 ;
			data[27347] <= 8'h10 ;
			data[27348] <= 8'h10 ;
			data[27349] <= 8'h10 ;
			data[27350] <= 8'h10 ;
			data[27351] <= 8'h10 ;
			data[27352] <= 8'h10 ;
			data[27353] <= 8'h10 ;
			data[27354] <= 8'h10 ;
			data[27355] <= 8'h10 ;
			data[27356] <= 8'h10 ;
			data[27357] <= 8'h10 ;
			data[27358] <= 8'h10 ;
			data[27359] <= 8'h10 ;
			data[27360] <= 8'h10 ;
			data[27361] <= 8'h10 ;
			data[27362] <= 8'h10 ;
			data[27363] <= 8'h10 ;
			data[27364] <= 8'h10 ;
			data[27365] <= 8'h10 ;
			data[27366] <= 8'h10 ;
			data[27367] <= 8'h10 ;
			data[27368] <= 8'h10 ;
			data[27369] <= 8'h10 ;
			data[27370] <= 8'h10 ;
			data[27371] <= 8'h10 ;
			data[27372] <= 8'h10 ;
			data[27373] <= 8'h10 ;
			data[27374] <= 8'h10 ;
			data[27375] <= 8'h10 ;
			data[27376] <= 8'h10 ;
			data[27377] <= 8'h10 ;
			data[27378] <= 8'h10 ;
			data[27379] <= 8'h10 ;
			data[27380] <= 8'h10 ;
			data[27381] <= 8'h10 ;
			data[27382] <= 8'h10 ;
			data[27383] <= 8'h10 ;
			data[27384] <= 8'h10 ;
			data[27385] <= 8'h10 ;
			data[27386] <= 8'h10 ;
			data[27387] <= 8'h10 ;
			data[27388] <= 8'h10 ;
			data[27389] <= 8'h10 ;
			data[27390] <= 8'h10 ;
			data[27391] <= 8'h10 ;
			data[27392] <= 8'h10 ;
			data[27393] <= 8'h10 ;
			data[27394] <= 8'h10 ;
			data[27395] <= 8'h10 ;
			data[27396] <= 8'h10 ;
			data[27397] <= 8'h10 ;
			data[27398] <= 8'h10 ;
			data[27399] <= 8'h10 ;
			data[27400] <= 8'h10 ;
			data[27401] <= 8'h10 ;
			data[27402] <= 8'h10 ;
			data[27403] <= 8'h10 ;
			data[27404] <= 8'h10 ;
			data[27405] <= 8'h10 ;
			data[27406] <= 8'h10 ;
			data[27407] <= 8'h10 ;
			data[27408] <= 8'h10 ;
			data[27409] <= 8'h10 ;
			data[27410] <= 8'h10 ;
			data[27411] <= 8'h10 ;
			data[27412] <= 8'h10 ;
			data[27413] <= 8'h10 ;
			data[27414] <= 8'h10 ;
			data[27415] <= 8'h10 ;
			data[27416] <= 8'h10 ;
			data[27417] <= 8'h10 ;
			data[27418] <= 8'h10 ;
			data[27419] <= 8'h10 ;
			data[27420] <= 8'h10 ;
			data[27421] <= 8'h10 ;
			data[27422] <= 8'h10 ;
			data[27423] <= 8'h10 ;
			data[27424] <= 8'h10 ;
			data[27425] <= 8'h10 ;
			data[27426] <= 8'h10 ;
			data[27427] <= 8'h10 ;
			data[27428] <= 8'h10 ;
			data[27429] <= 8'h10 ;
			data[27430] <= 8'h10 ;
			data[27431] <= 8'h10 ;
			data[27432] <= 8'h10 ;
			data[27433] <= 8'h10 ;
			data[27434] <= 8'h10 ;
			data[27435] <= 8'h10 ;
			data[27436] <= 8'h10 ;
			data[27437] <= 8'h10 ;
			data[27438] <= 8'h10 ;
			data[27439] <= 8'h10 ;
			data[27440] <= 8'h10 ;
			data[27441] <= 8'h10 ;
			data[27442] <= 8'h10 ;
			data[27443] <= 8'h10 ;
			data[27444] <= 8'h10 ;
			data[27445] <= 8'h10 ;
			data[27446] <= 8'h10 ;
			data[27447] <= 8'h10 ;
			data[27448] <= 8'h10 ;
			data[27449] <= 8'h10 ;
			data[27450] <= 8'h10 ;
			data[27451] <= 8'h10 ;
			data[27452] <= 8'h10 ;
			data[27453] <= 8'h10 ;
			data[27454] <= 8'h10 ;
			data[27455] <= 8'h10 ;
			data[27456] <= 8'h10 ;
			data[27457] <= 8'h10 ;
			data[27458] <= 8'h10 ;
			data[27459] <= 8'h10 ;
			data[27460] <= 8'h10 ;
			data[27461] <= 8'h10 ;
			data[27462] <= 8'h10 ;
			data[27463] <= 8'h10 ;
			data[27464] <= 8'h10 ;
			data[27465] <= 8'h10 ;
			data[27466] <= 8'h10 ;
			data[27467] <= 8'h10 ;
			data[27468] <= 8'h10 ;
			data[27469] <= 8'h10 ;
			data[27470] <= 8'h10 ;
			data[27471] <= 8'h10 ;
			data[27472] <= 8'h10 ;
			data[27473] <= 8'h10 ;
			data[27474] <= 8'h10 ;
			data[27475] <= 8'h10 ;
			data[27476] <= 8'h10 ;
			data[27477] <= 8'h10 ;
			data[27478] <= 8'h10 ;
			data[27479] <= 8'h10 ;
			data[27480] <= 8'h10 ;
			data[27481] <= 8'h10 ;
			data[27482] <= 8'h10 ;
			data[27483] <= 8'h10 ;
			data[27484] <= 8'h10 ;
			data[27485] <= 8'h10 ;
			data[27486] <= 8'h10 ;
			data[27487] <= 8'h10 ;
			data[27488] <= 8'h10 ;
			data[27489] <= 8'h10 ;
			data[27490] <= 8'h10 ;
			data[27491] <= 8'h10 ;
			data[27492] <= 8'h10 ;
			data[27493] <= 8'h10 ;
			data[27494] <= 8'h10 ;
			data[27495] <= 8'h10 ;
			data[27496] <= 8'h10 ;
			data[27497] <= 8'h10 ;
			data[27498] <= 8'h10 ;
			data[27499] <= 8'h10 ;
			data[27500] <= 8'h10 ;
			data[27501] <= 8'h10 ;
			data[27502] <= 8'h10 ;
			data[27503] <= 8'h10 ;
			data[27504] <= 8'h10 ;
			data[27505] <= 8'h10 ;
			data[27506] <= 8'h10 ;
			data[27507] <= 8'h10 ;
			data[27508] <= 8'h10 ;
			data[27509] <= 8'h10 ;
			data[27510] <= 8'h10 ;
			data[27511] <= 8'h10 ;
			data[27512] <= 8'h10 ;
			data[27513] <= 8'h10 ;
			data[27514] <= 8'h10 ;
			data[27515] <= 8'h10 ;
			data[27516] <= 8'h10 ;
			data[27517] <= 8'h10 ;
			data[27518] <= 8'h10 ;
			data[27519] <= 8'h10 ;
			data[27520] <= 8'h10 ;
			data[27521] <= 8'h10 ;
			data[27522] <= 8'h10 ;
			data[27523] <= 8'h10 ;
			data[27524] <= 8'h10 ;
			data[27525] <= 8'h10 ;
			data[27526] <= 8'h10 ;
			data[27527] <= 8'h10 ;
			data[27528] <= 8'h10 ;
			data[27529] <= 8'h10 ;
			data[27530] <= 8'h10 ;
			data[27531] <= 8'h10 ;
			data[27532] <= 8'h10 ;
			data[27533] <= 8'h10 ;
			data[27534] <= 8'h10 ;
			data[27535] <= 8'h10 ;
			data[27536] <= 8'h10 ;
			data[27537] <= 8'h10 ;
			data[27538] <= 8'h10 ;
			data[27539] <= 8'h10 ;
			data[27540] <= 8'h10 ;
			data[27541] <= 8'h10 ;
			data[27542] <= 8'h10 ;
			data[27543] <= 8'h10 ;
			data[27544] <= 8'h10 ;
			data[27545] <= 8'h10 ;
			data[27546] <= 8'h10 ;
			data[27547] <= 8'h10 ;
			data[27548] <= 8'h10 ;
			data[27549] <= 8'h10 ;
			data[27550] <= 8'h10 ;
			data[27551] <= 8'h10 ;
			data[27552] <= 8'h10 ;
			data[27553] <= 8'h10 ;
			data[27554] <= 8'h10 ;
			data[27555] <= 8'h10 ;
			data[27556] <= 8'h10 ;
			data[27557] <= 8'h10 ;
			data[27558] <= 8'h10 ;
			data[27559] <= 8'h10 ;
			data[27560] <= 8'h10 ;
			data[27561] <= 8'h10 ;
			data[27562] <= 8'h10 ;
			data[27563] <= 8'h10 ;
			data[27564] <= 8'h10 ;
			data[27565] <= 8'h10 ;
			data[27566] <= 8'h10 ;
			data[27567] <= 8'h10 ;
			data[27568] <= 8'h10 ;
			data[27569] <= 8'h10 ;
			data[27570] <= 8'h10 ;
			data[27571] <= 8'h10 ;
			data[27572] <= 8'h10 ;
			data[27573] <= 8'h10 ;
			data[27574] <= 8'h10 ;
			data[27575] <= 8'h10 ;
			data[27576] <= 8'h10 ;
			data[27577] <= 8'h10 ;
			data[27578] <= 8'h10 ;
			data[27579] <= 8'h10 ;
			data[27580] <= 8'h10 ;
			data[27581] <= 8'h10 ;
			data[27582] <= 8'h10 ;
			data[27583] <= 8'h10 ;
			data[27584] <= 8'h10 ;
			data[27585] <= 8'h10 ;
			data[27586] <= 8'h10 ;
			data[27587] <= 8'h10 ;
			data[27588] <= 8'h10 ;
			data[27589] <= 8'h10 ;
			data[27590] <= 8'h10 ;
			data[27591] <= 8'h10 ;
			data[27592] <= 8'h10 ;
			data[27593] <= 8'h10 ;
			data[27594] <= 8'h10 ;
			data[27595] <= 8'h10 ;
			data[27596] <= 8'h10 ;
			data[27597] <= 8'h10 ;
			data[27598] <= 8'h10 ;
			data[27599] <= 8'h10 ;
			data[27600] <= 8'h10 ;
			data[27601] <= 8'h10 ;
			data[27602] <= 8'h10 ;
			data[27603] <= 8'h10 ;
			data[27604] <= 8'h10 ;
			data[27605] <= 8'h10 ;
			data[27606] <= 8'h10 ;
			data[27607] <= 8'h10 ;
			data[27608] <= 8'h10 ;
			data[27609] <= 8'h10 ;
			data[27610] <= 8'h10 ;
			data[27611] <= 8'h10 ;
			data[27612] <= 8'h10 ;
			data[27613] <= 8'h10 ;
			data[27614] <= 8'h10 ;
			data[27615] <= 8'h10 ;
			data[27616] <= 8'h10 ;
			data[27617] <= 8'h10 ;
			data[27618] <= 8'h10 ;
			data[27619] <= 8'h10 ;
			data[27620] <= 8'h10 ;
			data[27621] <= 8'h10 ;
			data[27622] <= 8'h10 ;
			data[27623] <= 8'h10 ;
			data[27624] <= 8'h10 ;
			data[27625] <= 8'h10 ;
			data[27626] <= 8'h10 ;
			data[27627] <= 8'h10 ;
			data[27628] <= 8'h10 ;
			data[27629] <= 8'h10 ;
			data[27630] <= 8'h10 ;
			data[27631] <= 8'h10 ;
			data[27632] <= 8'h10 ;
			data[27633] <= 8'h10 ;
			data[27634] <= 8'h10 ;
			data[27635] <= 8'h10 ;
			data[27636] <= 8'h10 ;
			data[27637] <= 8'h10 ;
			data[27638] <= 8'h10 ;
			data[27639] <= 8'h10 ;
			data[27640] <= 8'h10 ;
			data[27641] <= 8'h10 ;
			data[27642] <= 8'h10 ;
			data[27643] <= 8'h10 ;
			data[27644] <= 8'h10 ;
			data[27645] <= 8'h10 ;
			data[27646] <= 8'h10 ;
			data[27647] <= 8'h10 ;
			data[27648] <= 8'h10 ;
			data[27649] <= 8'h10 ;
			data[27650] <= 8'h10 ;
			data[27651] <= 8'h10 ;
			data[27652] <= 8'h10 ;
			data[27653] <= 8'h10 ;
			data[27654] <= 8'h10 ;
			data[27655] <= 8'h10 ;
			data[27656] <= 8'h10 ;
			data[27657] <= 8'h10 ;
			data[27658] <= 8'h10 ;
			data[27659] <= 8'h10 ;
			data[27660] <= 8'h10 ;
			data[27661] <= 8'h10 ;
			data[27662] <= 8'h10 ;
			data[27663] <= 8'h10 ;
			data[27664] <= 8'h10 ;
			data[27665] <= 8'h10 ;
			data[27666] <= 8'h10 ;
			data[27667] <= 8'h10 ;
			data[27668] <= 8'h10 ;
			data[27669] <= 8'h10 ;
			data[27670] <= 8'h10 ;
			data[27671] <= 8'h10 ;
			data[27672] <= 8'h10 ;
			data[27673] <= 8'h10 ;
			data[27674] <= 8'h10 ;
			data[27675] <= 8'h10 ;
			data[27676] <= 8'h10 ;
			data[27677] <= 8'h10 ;
			data[27678] <= 8'h10 ;
			data[27679] <= 8'h10 ;
			data[27680] <= 8'h10 ;
			data[27681] <= 8'h10 ;
			data[27682] <= 8'h10 ;
			data[27683] <= 8'h10 ;
			data[27684] <= 8'h10 ;
			data[27685] <= 8'h10 ;
			data[27686] <= 8'h10 ;
			data[27687] <= 8'h10 ;
			data[27688] <= 8'h10 ;
			data[27689] <= 8'h10 ;
			data[27690] <= 8'h10 ;
			data[27691] <= 8'h10 ;
			data[27692] <= 8'h10 ;
			data[27693] <= 8'h10 ;
			data[27694] <= 8'h10 ;
			data[27695] <= 8'h10 ;
			data[27696] <= 8'h10 ;
			data[27697] <= 8'h10 ;
			data[27698] <= 8'h10 ;
			data[27699] <= 8'h10 ;
			data[27700] <= 8'h10 ;
			data[27701] <= 8'h10 ;
			data[27702] <= 8'h10 ;
			data[27703] <= 8'h10 ;
			data[27704] <= 8'h10 ;
			data[27705] <= 8'h10 ;
			data[27706] <= 8'h10 ;
			data[27707] <= 8'h10 ;
			data[27708] <= 8'h10 ;
			data[27709] <= 8'h10 ;
			data[27710] <= 8'h10 ;
			data[27711] <= 8'h10 ;
			data[27712] <= 8'h10 ;
			data[27713] <= 8'h10 ;
			data[27714] <= 8'h10 ;
			data[27715] <= 8'h10 ;
			data[27716] <= 8'h10 ;
			data[27717] <= 8'h10 ;
			data[27718] <= 8'h10 ;
			data[27719] <= 8'h10 ;
			data[27720] <= 8'h10 ;
			data[27721] <= 8'h10 ;
			data[27722] <= 8'h10 ;
			data[27723] <= 8'h10 ;
			data[27724] <= 8'h10 ;
			data[27725] <= 8'h10 ;
			data[27726] <= 8'h10 ;
			data[27727] <= 8'h10 ;
			data[27728] <= 8'h10 ;
			data[27729] <= 8'h10 ;
			data[27730] <= 8'h10 ;
			data[27731] <= 8'h10 ;
			data[27732] <= 8'h10 ;
			data[27733] <= 8'h10 ;
			data[27734] <= 8'h10 ;
			data[27735] <= 8'h10 ;
			data[27736] <= 8'h10 ;
			data[27737] <= 8'h10 ;
			data[27738] <= 8'h10 ;
			data[27739] <= 8'h10 ;
			data[27740] <= 8'h10 ;
			data[27741] <= 8'h10 ;
			data[27742] <= 8'h10 ;
			data[27743] <= 8'h10 ;
			data[27744] <= 8'h10 ;
			data[27745] <= 8'h10 ;
			data[27746] <= 8'h10 ;
			data[27747] <= 8'h10 ;
			data[27748] <= 8'h10 ;
			data[27749] <= 8'h10 ;
			data[27750] <= 8'h10 ;
			data[27751] <= 8'h10 ;
			data[27752] <= 8'h10 ;
			data[27753] <= 8'h10 ;
			data[27754] <= 8'h10 ;
			data[27755] <= 8'h10 ;
			data[27756] <= 8'h10 ;
			data[27757] <= 8'h10 ;
			data[27758] <= 8'h10 ;
			data[27759] <= 8'h10 ;
			data[27760] <= 8'h10 ;
			data[27761] <= 8'h10 ;
			data[27762] <= 8'h10 ;
			data[27763] <= 8'h10 ;
			data[27764] <= 8'h10 ;
			data[27765] <= 8'h10 ;
			data[27766] <= 8'h10 ;
			data[27767] <= 8'h10 ;
			data[27768] <= 8'h10 ;
			data[27769] <= 8'h10 ;
			data[27770] <= 8'h10 ;
			data[27771] <= 8'h10 ;
			data[27772] <= 8'h10 ;
			data[27773] <= 8'h10 ;
			data[27774] <= 8'h10 ;
			data[27775] <= 8'h10 ;
			data[27776] <= 8'h10 ;
			data[27777] <= 8'h10 ;
			data[27778] <= 8'h10 ;
			data[27779] <= 8'h10 ;
			data[27780] <= 8'h10 ;
			data[27781] <= 8'h10 ;
			data[27782] <= 8'h10 ;
			data[27783] <= 8'h10 ;
			data[27784] <= 8'h10 ;
			data[27785] <= 8'h10 ;
			data[27786] <= 8'h10 ;
			data[27787] <= 8'h10 ;
			data[27788] <= 8'h10 ;
			data[27789] <= 8'h10 ;
			data[27790] <= 8'h10 ;
			data[27791] <= 8'h10 ;
			data[27792] <= 8'h10 ;
			data[27793] <= 8'h10 ;
			data[27794] <= 8'h10 ;
			data[27795] <= 8'h10 ;
			data[27796] <= 8'h10 ;
			data[27797] <= 8'h10 ;
			data[27798] <= 8'h10 ;
			data[27799] <= 8'h10 ;
			data[27800] <= 8'h10 ;
			data[27801] <= 8'h10 ;
			data[27802] <= 8'h10 ;
			data[27803] <= 8'h10 ;
			data[27804] <= 8'h10 ;
			data[27805] <= 8'h10 ;
			data[27806] <= 8'h10 ;
			data[27807] <= 8'h10 ;
			data[27808] <= 8'h10 ;
			data[27809] <= 8'h10 ;
			data[27810] <= 8'h10 ;
			data[27811] <= 8'h10 ;
			data[27812] <= 8'h10 ;
			data[27813] <= 8'h10 ;
			data[27814] <= 8'h10 ;
			data[27815] <= 8'h10 ;
			data[27816] <= 8'h10 ;
			data[27817] <= 8'h10 ;
			data[27818] <= 8'h10 ;
			data[27819] <= 8'h10 ;
			data[27820] <= 8'h10 ;
			data[27821] <= 8'h10 ;
			data[27822] <= 8'h10 ;
			data[27823] <= 8'h10 ;
			data[27824] <= 8'h10 ;
			data[27825] <= 8'h10 ;
			data[27826] <= 8'h10 ;
			data[27827] <= 8'h10 ;
			data[27828] <= 8'h10 ;
			data[27829] <= 8'h10 ;
			data[27830] <= 8'h10 ;
			data[27831] <= 8'h10 ;
			data[27832] <= 8'h10 ;
			data[27833] <= 8'h10 ;
			data[27834] <= 8'h10 ;
			data[27835] <= 8'h10 ;
			data[27836] <= 8'h10 ;
			data[27837] <= 8'h10 ;
			data[27838] <= 8'h10 ;
			data[27839] <= 8'h10 ;
			data[27840] <= 8'h10 ;
			data[27841] <= 8'h10 ;
			data[27842] <= 8'h10 ;
			data[27843] <= 8'h10 ;
			data[27844] <= 8'h10 ;
			data[27845] <= 8'h10 ;
			data[27846] <= 8'h10 ;
			data[27847] <= 8'h10 ;
			data[27848] <= 8'h10 ;
			data[27849] <= 8'h10 ;
			data[27850] <= 8'h10 ;
			data[27851] <= 8'h10 ;
			data[27852] <= 8'h10 ;
			data[27853] <= 8'h10 ;
			data[27854] <= 8'h10 ;
			data[27855] <= 8'h10 ;
			data[27856] <= 8'h10 ;
			data[27857] <= 8'h10 ;
			data[27858] <= 8'h10 ;
			data[27859] <= 8'h10 ;
			data[27860] <= 8'h10 ;
			data[27861] <= 8'h10 ;
			data[27862] <= 8'h10 ;
			data[27863] <= 8'h10 ;
			data[27864] <= 8'h10 ;
			data[27865] <= 8'h10 ;
			data[27866] <= 8'h10 ;
			data[27867] <= 8'h10 ;
			data[27868] <= 8'h10 ;
			data[27869] <= 8'h10 ;
			data[27870] <= 8'h10 ;
			data[27871] <= 8'h10 ;
			data[27872] <= 8'h10 ;
			data[27873] <= 8'h10 ;
			data[27874] <= 8'h10 ;
			data[27875] <= 8'h10 ;
			data[27876] <= 8'h10 ;
			data[27877] <= 8'h10 ;
			data[27878] <= 8'h10 ;
			data[27879] <= 8'h10 ;
			data[27880] <= 8'h10 ;
			data[27881] <= 8'h10 ;
			data[27882] <= 8'h10 ;
			data[27883] <= 8'h10 ;
			data[27884] <= 8'h10 ;
			data[27885] <= 8'h10 ;
			data[27886] <= 8'h10 ;
			data[27887] <= 8'h10 ;
			data[27888] <= 8'h10 ;
			data[27889] <= 8'h10 ;
			data[27890] <= 8'h10 ;
			data[27891] <= 8'h10 ;
			data[27892] <= 8'h10 ;
			data[27893] <= 8'h10 ;
			data[27894] <= 8'h10 ;
			data[27895] <= 8'h10 ;
			data[27896] <= 8'h10 ;
			data[27897] <= 8'h10 ;
			data[27898] <= 8'h10 ;
			data[27899] <= 8'h10 ;
			data[27900] <= 8'h10 ;
			data[27901] <= 8'h10 ;
			data[27902] <= 8'h10 ;
			data[27903] <= 8'h10 ;
			data[27904] <= 8'h10 ;
			data[27905] <= 8'h10 ;
			data[27906] <= 8'h10 ;
			data[27907] <= 8'h10 ;
			data[27908] <= 8'h10 ;
			data[27909] <= 8'h10 ;
			data[27910] <= 8'h10 ;
			data[27911] <= 8'h10 ;
			data[27912] <= 8'h10 ;
			data[27913] <= 8'h10 ;
			data[27914] <= 8'h10 ;
			data[27915] <= 8'h10 ;
			data[27916] <= 8'h10 ;
			data[27917] <= 8'h10 ;
			data[27918] <= 8'h10 ;
			data[27919] <= 8'h10 ;
			data[27920] <= 8'h10 ;
			data[27921] <= 8'h10 ;
			data[27922] <= 8'h10 ;
			data[27923] <= 8'h10 ;
			data[27924] <= 8'h10 ;
			data[27925] <= 8'h10 ;
			data[27926] <= 8'h10 ;
			data[27927] <= 8'h10 ;
			data[27928] <= 8'h10 ;
			data[27929] <= 8'h10 ;
			data[27930] <= 8'h10 ;
			data[27931] <= 8'h10 ;
			data[27932] <= 8'h10 ;
			data[27933] <= 8'h10 ;
			data[27934] <= 8'h10 ;
			data[27935] <= 8'h10 ;
			data[27936] <= 8'h10 ;
			data[27937] <= 8'h10 ;
			data[27938] <= 8'h10 ;
			data[27939] <= 8'h10 ;
			data[27940] <= 8'h10 ;
			data[27941] <= 8'h10 ;
			data[27942] <= 8'h10 ;
			data[27943] <= 8'h10 ;
			data[27944] <= 8'h10 ;
			data[27945] <= 8'h10 ;
			data[27946] <= 8'h10 ;
			data[27947] <= 8'h10 ;
			data[27948] <= 8'h10 ;
			data[27949] <= 8'h10 ;
			data[27950] <= 8'h10 ;
			data[27951] <= 8'h10 ;
			data[27952] <= 8'h10 ;
			data[27953] <= 8'h10 ;
			data[27954] <= 8'h10 ;
			data[27955] <= 8'h10 ;
			data[27956] <= 8'h10 ;
			data[27957] <= 8'h10 ;
			data[27958] <= 8'h10 ;
			data[27959] <= 8'h10 ;
			data[27960] <= 8'h10 ;
			data[27961] <= 8'h10 ;
			data[27962] <= 8'h10 ;
			data[27963] <= 8'h10 ;
			data[27964] <= 8'h10 ;
			data[27965] <= 8'h10 ;
			data[27966] <= 8'h10 ;
			data[27967] <= 8'h10 ;
			data[27968] <= 8'h10 ;
			data[27969] <= 8'h10 ;
			data[27970] <= 8'h10 ;
			data[27971] <= 8'h10 ;
			data[27972] <= 8'h10 ;
			data[27973] <= 8'h10 ;
			data[27974] <= 8'h10 ;
			data[27975] <= 8'h10 ;
			data[27976] <= 8'h10 ;
			data[27977] <= 8'h10 ;
			data[27978] <= 8'h10 ;
			data[27979] <= 8'h10 ;
			data[27980] <= 8'h10 ;
			data[27981] <= 8'h10 ;
			data[27982] <= 8'h10 ;
			data[27983] <= 8'h10 ;
			data[27984] <= 8'h10 ;
			data[27985] <= 8'h10 ;
			data[27986] <= 8'h10 ;
			data[27987] <= 8'h10 ;
			data[27988] <= 8'h10 ;
			data[27989] <= 8'h10 ;
			data[27990] <= 8'h10 ;
			data[27991] <= 8'h10 ;
			data[27992] <= 8'h10 ;
			data[27993] <= 8'h10 ;
			data[27994] <= 8'h10 ;
			data[27995] <= 8'h10 ;
			data[27996] <= 8'h10 ;
			data[27997] <= 8'h10 ;
			data[27998] <= 8'h10 ;
			data[27999] <= 8'h10 ;
			data[28000] <= 8'h10 ;
			data[28001] <= 8'h10 ;
			data[28002] <= 8'h10 ;
			data[28003] <= 8'h10 ;
			data[28004] <= 8'h10 ;
			data[28005] <= 8'h10 ;
			data[28006] <= 8'h10 ;
			data[28007] <= 8'h10 ;
			data[28008] <= 8'h10 ;
			data[28009] <= 8'h10 ;
			data[28010] <= 8'h10 ;
			data[28011] <= 8'h10 ;
			data[28012] <= 8'h10 ;
			data[28013] <= 8'h10 ;
			data[28014] <= 8'h10 ;
			data[28015] <= 8'h10 ;
			data[28016] <= 8'h10 ;
			data[28017] <= 8'h10 ;
			data[28018] <= 8'h10 ;
			data[28019] <= 8'h10 ;
			data[28020] <= 8'h10 ;
			data[28021] <= 8'h10 ;
			data[28022] <= 8'h10 ;
			data[28023] <= 8'h10 ;
			data[28024] <= 8'h10 ;
			data[28025] <= 8'h10 ;
			data[28026] <= 8'h10 ;
			data[28027] <= 8'h10 ;
			data[28028] <= 8'h10 ;
			data[28029] <= 8'h10 ;
			data[28030] <= 8'h10 ;
			data[28031] <= 8'h10 ;
			data[28032] <= 8'h10 ;
			data[28033] <= 8'h10 ;
			data[28034] <= 8'h10 ;
			data[28035] <= 8'h10 ;
			data[28036] <= 8'h10 ;
			data[28037] <= 8'h10 ;
			data[28038] <= 8'h10 ;
			data[28039] <= 8'h10 ;
			data[28040] <= 8'h10 ;
			data[28041] <= 8'h10 ;
			data[28042] <= 8'h10 ;
			data[28043] <= 8'h10 ;
			data[28044] <= 8'h10 ;
			data[28045] <= 8'h10 ;
			data[28046] <= 8'h10 ;
			data[28047] <= 8'h10 ;
			data[28048] <= 8'h10 ;
			data[28049] <= 8'h10 ;
			data[28050] <= 8'h10 ;
			data[28051] <= 8'h10 ;
			data[28052] <= 8'h10 ;
			data[28053] <= 8'h10 ;
			data[28054] <= 8'h10 ;
			data[28055] <= 8'h10 ;
			data[28056] <= 8'h10 ;
			data[28057] <= 8'h10 ;
			data[28058] <= 8'h10 ;
			data[28059] <= 8'h10 ;
			data[28060] <= 8'h10 ;
			data[28061] <= 8'h10 ;
			data[28062] <= 8'h10 ;
			data[28063] <= 8'h10 ;
			data[28064] <= 8'h10 ;
			data[28065] <= 8'h10 ;
			data[28066] <= 8'h10 ;
			data[28067] <= 8'h10 ;
			data[28068] <= 8'h10 ;
			data[28069] <= 8'h10 ;
			data[28070] <= 8'h10 ;
			data[28071] <= 8'h10 ;
			data[28072] <= 8'h10 ;
			data[28073] <= 8'h10 ;
			data[28074] <= 8'h10 ;
			data[28075] <= 8'h10 ;
			data[28076] <= 8'h10 ;
			data[28077] <= 8'h10 ;
			data[28078] <= 8'h10 ;
			data[28079] <= 8'h10 ;
			data[28080] <= 8'h10 ;
			data[28081] <= 8'h10 ;
			data[28082] <= 8'h10 ;
			data[28083] <= 8'h10 ;
			data[28084] <= 8'h10 ;
			data[28085] <= 8'h10 ;
			data[28086] <= 8'h10 ;
			data[28087] <= 8'h10 ;
			data[28088] <= 8'h10 ;
			data[28089] <= 8'h10 ;
			data[28090] <= 8'h10 ;
			data[28091] <= 8'h10 ;
			data[28092] <= 8'h10 ;
			data[28093] <= 8'h10 ;
			data[28094] <= 8'h10 ;
			data[28095] <= 8'h10 ;
			data[28096] <= 8'h10 ;
			data[28097] <= 8'h10 ;
			data[28098] <= 8'h10 ;
			data[28099] <= 8'h10 ;
			data[28100] <= 8'h10 ;
			data[28101] <= 8'h10 ;
			data[28102] <= 8'h10 ;
			data[28103] <= 8'h10 ;
			data[28104] <= 8'h10 ;
			data[28105] <= 8'h10 ;
			data[28106] <= 8'h10 ;
			data[28107] <= 8'h10 ;
			data[28108] <= 8'h10 ;
			data[28109] <= 8'h10 ;
			data[28110] <= 8'h10 ;
			data[28111] <= 8'h10 ;
			data[28112] <= 8'h10 ;
			data[28113] <= 8'h10 ;
			data[28114] <= 8'h10 ;
			data[28115] <= 8'h10 ;
			data[28116] <= 8'h10 ;
			data[28117] <= 8'h10 ;
			data[28118] <= 8'h10 ;
			data[28119] <= 8'h10 ;
			data[28120] <= 8'h10 ;
			data[28121] <= 8'h10 ;
			data[28122] <= 8'h10 ;
			data[28123] <= 8'h10 ;
			data[28124] <= 8'h10 ;
			data[28125] <= 8'h10 ;
			data[28126] <= 8'h10 ;
			data[28127] <= 8'h10 ;
			data[28128] <= 8'h10 ;
			data[28129] <= 8'h10 ;
			data[28130] <= 8'h10 ;
			data[28131] <= 8'h10 ;
			data[28132] <= 8'h10 ;
			data[28133] <= 8'h10 ;
			data[28134] <= 8'h10 ;
			data[28135] <= 8'h10 ;
			data[28136] <= 8'h10 ;
			data[28137] <= 8'h10 ;
			data[28138] <= 8'h10 ;
			data[28139] <= 8'h10 ;
			data[28140] <= 8'h10 ;
			data[28141] <= 8'h10 ;
			data[28142] <= 8'h10 ;
			data[28143] <= 8'h10 ;
			data[28144] <= 8'h10 ;
			data[28145] <= 8'h10 ;
			data[28146] <= 8'h10 ;
			data[28147] <= 8'h10 ;
			data[28148] <= 8'h10 ;
			data[28149] <= 8'h10 ;
			data[28150] <= 8'h10 ;
			data[28151] <= 8'h10 ;
			data[28152] <= 8'h10 ;
			data[28153] <= 8'h10 ;
			data[28154] <= 8'h10 ;
			data[28155] <= 8'h10 ;
			data[28156] <= 8'h10 ;
			data[28157] <= 8'h10 ;
			data[28158] <= 8'h10 ;
			data[28159] <= 8'h10 ;
			data[28160] <= 8'h10 ;
			data[28161] <= 8'h10 ;
			data[28162] <= 8'h10 ;
			data[28163] <= 8'h10 ;
			data[28164] <= 8'h10 ;
			data[28165] <= 8'h10 ;
			data[28166] <= 8'h10 ;
			data[28167] <= 8'h10 ;
			data[28168] <= 8'h10 ;
			data[28169] <= 8'h10 ;
			data[28170] <= 8'h10 ;
			data[28171] <= 8'h10 ;
			data[28172] <= 8'h10 ;
			data[28173] <= 8'h10 ;
			data[28174] <= 8'h10 ;
			data[28175] <= 8'h10 ;
			data[28176] <= 8'h10 ;
			data[28177] <= 8'h10 ;
			data[28178] <= 8'h10 ;
			data[28179] <= 8'h10 ;
			data[28180] <= 8'h10 ;
			data[28181] <= 8'h10 ;
			data[28182] <= 8'h10 ;
			data[28183] <= 8'h10 ;
			data[28184] <= 8'h10 ;
			data[28185] <= 8'h10 ;
			data[28186] <= 8'h10 ;
			data[28187] <= 8'h10 ;
			data[28188] <= 8'h10 ;
			data[28189] <= 8'h10 ;
			data[28190] <= 8'h10 ;
			data[28191] <= 8'h10 ;
			data[28192] <= 8'h10 ;
			data[28193] <= 8'h10 ;
			data[28194] <= 8'h10 ;
			data[28195] <= 8'h10 ;
			data[28196] <= 8'h10 ;
			data[28197] <= 8'h10 ;
			data[28198] <= 8'h10 ;
			data[28199] <= 8'h10 ;
			data[28200] <= 8'h10 ;
			data[28201] <= 8'h10 ;
			data[28202] <= 8'h10 ;
			data[28203] <= 8'h10 ;
			data[28204] <= 8'h10 ;
			data[28205] <= 8'h10 ;
			data[28206] <= 8'h10 ;
			data[28207] <= 8'h10 ;
			data[28208] <= 8'h10 ;
			data[28209] <= 8'h10 ;
			data[28210] <= 8'h10 ;
			data[28211] <= 8'h10 ;
			data[28212] <= 8'h10 ;
			data[28213] <= 8'h10 ;
			data[28214] <= 8'h10 ;
			data[28215] <= 8'h10 ;
			data[28216] <= 8'h10 ;
			data[28217] <= 8'h10 ;
			data[28218] <= 8'h10 ;
			data[28219] <= 8'h10 ;
			data[28220] <= 8'h10 ;
			data[28221] <= 8'h10 ;
			data[28222] <= 8'h10 ;
			data[28223] <= 8'h10 ;
			data[28224] <= 8'h10 ;
			data[28225] <= 8'h10 ;
			data[28226] <= 8'h10 ;
			data[28227] <= 8'h10 ;
			data[28228] <= 8'h10 ;
			data[28229] <= 8'h10 ;
			data[28230] <= 8'h10 ;
			data[28231] <= 8'h10 ;
			data[28232] <= 8'h10 ;
			data[28233] <= 8'h10 ;
			data[28234] <= 8'h10 ;
			data[28235] <= 8'h10 ;
			data[28236] <= 8'h10 ;
			data[28237] <= 8'h10 ;
			data[28238] <= 8'h10 ;
			data[28239] <= 8'h10 ;
			data[28240] <= 8'h10 ;
			data[28241] <= 8'h10 ;
			data[28242] <= 8'h10 ;
			data[28243] <= 8'h10 ;
			data[28244] <= 8'h10 ;
			data[28245] <= 8'h10 ;
			data[28246] <= 8'h10 ;
			data[28247] <= 8'h10 ;
			data[28248] <= 8'h10 ;
			data[28249] <= 8'h10 ;
			data[28250] <= 8'h10 ;
			data[28251] <= 8'h10 ;
			data[28252] <= 8'h10 ;
			data[28253] <= 8'h10 ;
			data[28254] <= 8'h10 ;
			data[28255] <= 8'h10 ;
			data[28256] <= 8'h10 ;
			data[28257] <= 8'h10 ;
			data[28258] <= 8'h10 ;
			data[28259] <= 8'h10 ;
			data[28260] <= 8'h10 ;
			data[28261] <= 8'h10 ;
			data[28262] <= 8'h10 ;
			data[28263] <= 8'h10 ;
			data[28264] <= 8'h10 ;
			data[28265] <= 8'h10 ;
			data[28266] <= 8'h10 ;
			data[28267] <= 8'h10 ;
			data[28268] <= 8'h10 ;
			data[28269] <= 8'h10 ;
			data[28270] <= 8'h10 ;
			data[28271] <= 8'h10 ;
			data[28272] <= 8'h10 ;
			data[28273] <= 8'h10 ;
			data[28274] <= 8'h10 ;
			data[28275] <= 8'h10 ;
			data[28276] <= 8'h10 ;
			data[28277] <= 8'h10 ;
			data[28278] <= 8'h10 ;
			data[28279] <= 8'h10 ;
			data[28280] <= 8'h10 ;
			data[28281] <= 8'h10 ;
			data[28282] <= 8'h10 ;
			data[28283] <= 8'h10 ;
			data[28284] <= 8'h10 ;
			data[28285] <= 8'h10 ;
			data[28286] <= 8'h10 ;
			data[28287] <= 8'h10 ;
			data[28288] <= 8'h10 ;
			data[28289] <= 8'h10 ;
			data[28290] <= 8'h10 ;
			data[28291] <= 8'h10 ;
			data[28292] <= 8'h10 ;
			data[28293] <= 8'h10 ;
			data[28294] <= 8'h10 ;
			data[28295] <= 8'h10 ;
			data[28296] <= 8'h10 ;
			data[28297] <= 8'h10 ;
			data[28298] <= 8'h10 ;
			data[28299] <= 8'h10 ;
			data[28300] <= 8'h10 ;
			data[28301] <= 8'h10 ;
			data[28302] <= 8'h10 ;
			data[28303] <= 8'h10 ;
			data[28304] <= 8'h10 ;
			data[28305] <= 8'h10 ;
			data[28306] <= 8'h10 ;
			data[28307] <= 8'h10 ;
			data[28308] <= 8'h10 ;
			data[28309] <= 8'h10 ;
			data[28310] <= 8'h10 ;
			data[28311] <= 8'h10 ;
			data[28312] <= 8'h10 ;
			data[28313] <= 8'h10 ;
			data[28314] <= 8'h10 ;
			data[28315] <= 8'h10 ;
			data[28316] <= 8'h10 ;
			data[28317] <= 8'h10 ;
			data[28318] <= 8'h10 ;
			data[28319] <= 8'h10 ;
			data[28320] <= 8'h10 ;
			data[28321] <= 8'h10 ;
			data[28322] <= 8'h10 ;
			data[28323] <= 8'h10 ;
			data[28324] <= 8'h10 ;
			data[28325] <= 8'h10 ;
			data[28326] <= 8'h10 ;
			data[28327] <= 8'h10 ;
			data[28328] <= 8'h10 ;
			data[28329] <= 8'h10 ;
			data[28330] <= 8'h10 ;
			data[28331] <= 8'h10 ;
			data[28332] <= 8'h10 ;
			data[28333] <= 8'h10 ;
			data[28334] <= 8'h10 ;
			data[28335] <= 8'h10 ;
			data[28336] <= 8'h10 ;
			data[28337] <= 8'h10 ;
			data[28338] <= 8'h10 ;
			data[28339] <= 8'h10 ;
			data[28340] <= 8'h10 ;
			data[28341] <= 8'h10 ;
			data[28342] <= 8'h10 ;
			data[28343] <= 8'h10 ;
			data[28344] <= 8'h10 ;
			data[28345] <= 8'h10 ;
			data[28346] <= 8'h10 ;
			data[28347] <= 8'h10 ;
			data[28348] <= 8'h10 ;
			data[28349] <= 8'h10 ;
			data[28350] <= 8'h10 ;
			data[28351] <= 8'h10 ;
			data[28352] <= 8'h10 ;
			data[28353] <= 8'h10 ;
			data[28354] <= 8'h10 ;
			data[28355] <= 8'h10 ;
			data[28356] <= 8'h10 ;
			data[28357] <= 8'h10 ;
			data[28358] <= 8'h10 ;
			data[28359] <= 8'h10 ;
			data[28360] <= 8'h10 ;
			data[28361] <= 8'h10 ;
			data[28362] <= 8'h10 ;
			data[28363] <= 8'h10 ;
			data[28364] <= 8'h10 ;
			data[28365] <= 8'h10 ;
			data[28366] <= 8'h10 ;
			data[28367] <= 8'h10 ;
			data[28368] <= 8'h10 ;
			data[28369] <= 8'h10 ;
			data[28370] <= 8'h10 ;
			data[28371] <= 8'h10 ;
			data[28372] <= 8'h10 ;
			data[28373] <= 8'h10 ;
			data[28374] <= 8'h10 ;
			data[28375] <= 8'h10 ;
			data[28376] <= 8'h10 ;
			data[28377] <= 8'h10 ;
			data[28378] <= 8'h10 ;
			data[28379] <= 8'h10 ;
			data[28380] <= 8'h10 ;
			data[28381] <= 8'h10 ;
			data[28382] <= 8'h10 ;
			data[28383] <= 8'h10 ;
			data[28384] <= 8'h10 ;
			data[28385] <= 8'h10 ;
			data[28386] <= 8'h10 ;
			data[28387] <= 8'h10 ;
			data[28388] <= 8'h10 ;
			data[28389] <= 8'h10 ;
			data[28390] <= 8'h10 ;
			data[28391] <= 8'h10 ;
			data[28392] <= 8'h10 ;
			data[28393] <= 8'h10 ;
			data[28394] <= 8'h10 ;
			data[28395] <= 8'h10 ;
			data[28396] <= 8'h10 ;
			data[28397] <= 8'h10 ;
			data[28398] <= 8'h10 ;
			data[28399] <= 8'h10 ;
			data[28400] <= 8'h10 ;
			data[28401] <= 8'h10 ;
			data[28402] <= 8'h10 ;
			data[28403] <= 8'h10 ;
			data[28404] <= 8'h10 ;
			data[28405] <= 8'h10 ;
			data[28406] <= 8'h10 ;
			data[28407] <= 8'h10 ;
			data[28408] <= 8'h10 ;
			data[28409] <= 8'h10 ;
			data[28410] <= 8'h10 ;
			data[28411] <= 8'h10 ;
			data[28412] <= 8'h10 ;
			data[28413] <= 8'h10 ;
			data[28414] <= 8'h10 ;
			data[28415] <= 8'h10 ;
			data[28416] <= 8'h10 ;
			data[28417] <= 8'h10 ;
			data[28418] <= 8'h10 ;
			data[28419] <= 8'h10 ;
			data[28420] <= 8'h10 ;
			data[28421] <= 8'h10 ;
			data[28422] <= 8'h10 ;
			data[28423] <= 8'h10 ;
			data[28424] <= 8'h10 ;
			data[28425] <= 8'h10 ;
			data[28426] <= 8'h10 ;
			data[28427] <= 8'h10 ;
			data[28428] <= 8'h10 ;
			data[28429] <= 8'h10 ;
			data[28430] <= 8'h10 ;
			data[28431] <= 8'h10 ;
			data[28432] <= 8'h10 ;
			data[28433] <= 8'h10 ;
			data[28434] <= 8'h10 ;
			data[28435] <= 8'h10 ;
			data[28436] <= 8'h10 ;
			data[28437] <= 8'h10 ;
			data[28438] <= 8'h10 ;
			data[28439] <= 8'h10 ;
			data[28440] <= 8'h10 ;
			data[28441] <= 8'h10 ;
			data[28442] <= 8'h10 ;
			data[28443] <= 8'h10 ;
			data[28444] <= 8'h10 ;
			data[28445] <= 8'h10 ;
			data[28446] <= 8'h10 ;
			data[28447] <= 8'h10 ;
			data[28448] <= 8'h10 ;
			data[28449] <= 8'h10 ;
			data[28450] <= 8'h10 ;
			data[28451] <= 8'h10 ;
			data[28452] <= 8'h10 ;
			data[28453] <= 8'h10 ;
			data[28454] <= 8'h10 ;
			data[28455] <= 8'h10 ;
			data[28456] <= 8'h10 ;
			data[28457] <= 8'h10 ;
			data[28458] <= 8'h10 ;
			data[28459] <= 8'h10 ;
			data[28460] <= 8'h10 ;
			data[28461] <= 8'h10 ;
			data[28462] <= 8'h10 ;
			data[28463] <= 8'h10 ;
			data[28464] <= 8'h10 ;
			data[28465] <= 8'h10 ;
			data[28466] <= 8'h10 ;
			data[28467] <= 8'h10 ;
			data[28468] <= 8'h10 ;
			data[28469] <= 8'h10 ;
			data[28470] <= 8'h10 ;
			data[28471] <= 8'h10 ;
			data[28472] <= 8'h10 ;
			data[28473] <= 8'h10 ;
			data[28474] <= 8'h10 ;
			data[28475] <= 8'h10 ;
			data[28476] <= 8'h10 ;
			data[28477] <= 8'h10 ;
			data[28478] <= 8'h10 ;
			data[28479] <= 8'h10 ;
			data[28480] <= 8'h10 ;
			data[28481] <= 8'h10 ;
			data[28482] <= 8'h10 ;
			data[28483] <= 8'h10 ;
			data[28484] <= 8'h10 ;
			data[28485] <= 8'h10 ;
			data[28486] <= 8'h10 ;
			data[28487] <= 8'h10 ;
			data[28488] <= 8'h10 ;
			data[28489] <= 8'h10 ;
			data[28490] <= 8'h10 ;
			data[28491] <= 8'h10 ;
			data[28492] <= 8'h10 ;
			data[28493] <= 8'h10 ;
			data[28494] <= 8'h10 ;
			data[28495] <= 8'h10 ;
			data[28496] <= 8'h10 ;
			data[28497] <= 8'h10 ;
			data[28498] <= 8'h10 ;
			data[28499] <= 8'h10 ;
			data[28500] <= 8'h10 ;
			data[28501] <= 8'h10 ;
			data[28502] <= 8'h10 ;
			data[28503] <= 8'h10 ;
			data[28504] <= 8'h10 ;
			data[28505] <= 8'h10 ;
			data[28506] <= 8'h10 ;
			data[28507] <= 8'h10 ;
			data[28508] <= 8'h10 ;
			data[28509] <= 8'h10 ;
			data[28510] <= 8'h10 ;
			data[28511] <= 8'h10 ;
			data[28512] <= 8'h10 ;
			data[28513] <= 8'h10 ;
			data[28514] <= 8'h10 ;
			data[28515] <= 8'h10 ;
			data[28516] <= 8'h10 ;
			data[28517] <= 8'h10 ;
			data[28518] <= 8'h10 ;
			data[28519] <= 8'h10 ;
			data[28520] <= 8'h10 ;
			data[28521] <= 8'h10 ;
			data[28522] <= 8'h10 ;
			data[28523] <= 8'h10 ;
			data[28524] <= 8'h10 ;
			data[28525] <= 8'h10 ;
			data[28526] <= 8'h10 ;
			data[28527] <= 8'h10 ;
			data[28528] <= 8'h10 ;
			data[28529] <= 8'h10 ;
			data[28530] <= 8'h10 ;
			data[28531] <= 8'h10 ;
			data[28532] <= 8'h10 ;
			data[28533] <= 8'h10 ;
			data[28534] <= 8'h10 ;
			data[28535] <= 8'h10 ;
			data[28536] <= 8'h10 ;
			data[28537] <= 8'h10 ;
			data[28538] <= 8'h10 ;
			data[28539] <= 8'h10 ;
			data[28540] <= 8'h10 ;
			data[28541] <= 8'h10 ;
			data[28542] <= 8'h10 ;
			data[28543] <= 8'h10 ;
			data[28544] <= 8'h10 ;
			data[28545] <= 8'h10 ;
			data[28546] <= 8'h10 ;
			data[28547] <= 8'h10 ;
			data[28548] <= 8'h10 ;
			data[28549] <= 8'h10 ;
			data[28550] <= 8'h10 ;
			data[28551] <= 8'h10 ;
			data[28552] <= 8'h10 ;
			data[28553] <= 8'h10 ;
			data[28554] <= 8'h10 ;
			data[28555] <= 8'h10 ;
			data[28556] <= 8'h10 ;
			data[28557] <= 8'h10 ;
			data[28558] <= 8'h10 ;
			data[28559] <= 8'h10 ;
			data[28560] <= 8'h10 ;
			data[28561] <= 8'h10 ;
			data[28562] <= 8'h10 ;
			data[28563] <= 8'h10 ;
			data[28564] <= 8'h10 ;
			data[28565] <= 8'h10 ;
			data[28566] <= 8'h10 ;
			data[28567] <= 8'h10 ;
			data[28568] <= 8'h10 ;
			data[28569] <= 8'h10 ;
			data[28570] <= 8'h10 ;
			data[28571] <= 8'h10 ;
			data[28572] <= 8'h10 ;
			data[28573] <= 8'h10 ;
			data[28574] <= 8'h10 ;
			data[28575] <= 8'h10 ;
			data[28576] <= 8'h10 ;
			data[28577] <= 8'h10 ;
			data[28578] <= 8'h10 ;
			data[28579] <= 8'h10 ;
			data[28580] <= 8'h10 ;
			data[28581] <= 8'h10 ;
			data[28582] <= 8'h10 ;
			data[28583] <= 8'h10 ;
			data[28584] <= 8'h10 ;
			data[28585] <= 8'h10 ;
			data[28586] <= 8'h10 ;
			data[28587] <= 8'h10 ;
			data[28588] <= 8'h10 ;
			data[28589] <= 8'h10 ;
			data[28590] <= 8'h10 ;
			data[28591] <= 8'h10 ;
			data[28592] <= 8'h10 ;
			data[28593] <= 8'h10 ;
			data[28594] <= 8'h10 ;
			data[28595] <= 8'h10 ;
			data[28596] <= 8'h10 ;
			data[28597] <= 8'h10 ;
			data[28598] <= 8'h10 ;
			data[28599] <= 8'h10 ;
			data[28600] <= 8'h10 ;
			data[28601] <= 8'h10 ;
			data[28602] <= 8'h10 ;
			data[28603] <= 8'h10 ;
			data[28604] <= 8'h10 ;
			data[28605] <= 8'h10 ;
			data[28606] <= 8'h10 ;
			data[28607] <= 8'h10 ;
			data[28608] <= 8'h10 ;
			data[28609] <= 8'h10 ;
			data[28610] <= 8'h10 ;
			data[28611] <= 8'h10 ;
			data[28612] <= 8'h10 ;
			data[28613] <= 8'h10 ;
			data[28614] <= 8'h10 ;
			data[28615] <= 8'h10 ;
			data[28616] <= 8'h10 ;
			data[28617] <= 8'h10 ;
			data[28618] <= 8'h10 ;
			data[28619] <= 8'h10 ;
			data[28620] <= 8'h10 ;
			data[28621] <= 8'h10 ;
			data[28622] <= 8'h10 ;
			data[28623] <= 8'h10 ;
			data[28624] <= 8'h10 ;
			data[28625] <= 8'h10 ;
			data[28626] <= 8'h10 ;
			data[28627] <= 8'h10 ;
			data[28628] <= 8'h10 ;
			data[28629] <= 8'h10 ;
			data[28630] <= 8'h10 ;
			data[28631] <= 8'h10 ;
			data[28632] <= 8'h10 ;
			data[28633] <= 8'h10 ;
			data[28634] <= 8'h10 ;
			data[28635] <= 8'h10 ;
			data[28636] <= 8'h10 ;
			data[28637] <= 8'h10 ;
			data[28638] <= 8'h10 ;
			data[28639] <= 8'h10 ;
			data[28640] <= 8'h10 ;
			data[28641] <= 8'h10 ;
			data[28642] <= 8'h10 ;
			data[28643] <= 8'h10 ;
			data[28644] <= 8'h10 ;
			data[28645] <= 8'h10 ;
			data[28646] <= 8'h10 ;
			data[28647] <= 8'h10 ;
			data[28648] <= 8'h10 ;
			data[28649] <= 8'h10 ;
			data[28650] <= 8'h10 ;
			data[28651] <= 8'h10 ;
			data[28652] <= 8'h10 ;
			data[28653] <= 8'h10 ;
			data[28654] <= 8'h10 ;
			data[28655] <= 8'h10 ;
			data[28656] <= 8'h10 ;
			data[28657] <= 8'h10 ;
			data[28658] <= 8'h10 ;
			data[28659] <= 8'h10 ;
			data[28660] <= 8'h10 ;
			data[28661] <= 8'h10 ;
			data[28662] <= 8'h10 ;
			data[28663] <= 8'h10 ;
			data[28664] <= 8'h10 ;
			data[28665] <= 8'h10 ;
			data[28666] <= 8'h10 ;
			data[28667] <= 8'h10 ;
			data[28668] <= 8'h10 ;
			data[28669] <= 8'h10 ;
			data[28670] <= 8'h10 ;
			data[28671] <= 8'h10 ;
			data[28672] <= 8'h10 ;
			data[28673] <= 8'h10 ;
			data[28674] <= 8'h10 ;
			data[28675] <= 8'h10 ;
			data[28676] <= 8'h10 ;
			data[28677] <= 8'h10 ;
			data[28678] <= 8'h10 ;
			data[28679] <= 8'h10 ;
			data[28680] <= 8'h10 ;
			data[28681] <= 8'h10 ;
			data[28682] <= 8'h10 ;
			data[28683] <= 8'h10 ;
			data[28684] <= 8'h10 ;
			data[28685] <= 8'h10 ;
			data[28686] <= 8'h10 ;
			data[28687] <= 8'h10 ;
			data[28688] <= 8'h10 ;
			data[28689] <= 8'h10 ;
			data[28690] <= 8'h10 ;
			data[28691] <= 8'h10 ;
			data[28692] <= 8'h10 ;
			data[28693] <= 8'h10 ;
			data[28694] <= 8'h10 ;
			data[28695] <= 8'h10 ;
			data[28696] <= 8'h10 ;
			data[28697] <= 8'h10 ;
			data[28698] <= 8'h10 ;
			data[28699] <= 8'h10 ;
			data[28700] <= 8'h10 ;
			data[28701] <= 8'h10 ;
			data[28702] <= 8'h10 ;
			data[28703] <= 8'h10 ;
			data[28704] <= 8'h10 ;
			data[28705] <= 8'h10 ;
			data[28706] <= 8'h10 ;
			data[28707] <= 8'h10 ;
			data[28708] <= 8'h10 ;
			data[28709] <= 8'h10 ;
			data[28710] <= 8'h10 ;
			data[28711] <= 8'h10 ;
			data[28712] <= 8'h10 ;
			data[28713] <= 8'h10 ;
			data[28714] <= 8'h10 ;
			data[28715] <= 8'h10 ;
			data[28716] <= 8'h10 ;
			data[28717] <= 8'h10 ;
			data[28718] <= 8'h10 ;
			data[28719] <= 8'h10 ;
			data[28720] <= 8'h10 ;
			data[28721] <= 8'h10 ;
			data[28722] <= 8'h10 ;
			data[28723] <= 8'h10 ;
			data[28724] <= 8'h10 ;
			data[28725] <= 8'h10 ;
			data[28726] <= 8'h10 ;
			data[28727] <= 8'h10 ;
			data[28728] <= 8'h10 ;
			data[28729] <= 8'h10 ;
			data[28730] <= 8'h10 ;
			data[28731] <= 8'h10 ;
			data[28732] <= 8'h10 ;
			data[28733] <= 8'h10 ;
			data[28734] <= 8'h10 ;
			data[28735] <= 8'h10 ;
			data[28736] <= 8'h10 ;
			data[28737] <= 8'h10 ;
			data[28738] <= 8'h10 ;
			data[28739] <= 8'h10 ;
			data[28740] <= 8'h10 ;
			data[28741] <= 8'h10 ;
			data[28742] <= 8'h10 ;
			data[28743] <= 8'h10 ;
			data[28744] <= 8'h10 ;
			data[28745] <= 8'h10 ;
			data[28746] <= 8'h10 ;
			data[28747] <= 8'h10 ;
			data[28748] <= 8'h10 ;
			data[28749] <= 8'h10 ;
			data[28750] <= 8'h10 ;
			data[28751] <= 8'h10 ;
			data[28752] <= 8'h10 ;
			data[28753] <= 8'h10 ;
			data[28754] <= 8'h10 ;
			data[28755] <= 8'h10 ;
			data[28756] <= 8'h10 ;
			data[28757] <= 8'h10 ;
			data[28758] <= 8'h10 ;
			data[28759] <= 8'h10 ;
			data[28760] <= 8'h10 ;
			data[28761] <= 8'h10 ;
			data[28762] <= 8'h10 ;
			data[28763] <= 8'h10 ;
			data[28764] <= 8'h10 ;
			data[28765] <= 8'h10 ;
			data[28766] <= 8'h10 ;
			data[28767] <= 8'h10 ;
			data[28768] <= 8'h10 ;
			data[28769] <= 8'h10 ;
			data[28770] <= 8'h10 ;
			data[28771] <= 8'h10 ;
			data[28772] <= 8'h10 ;
			data[28773] <= 8'h10 ;
			data[28774] <= 8'h10 ;
			data[28775] <= 8'h10 ;
			data[28776] <= 8'h10 ;
			data[28777] <= 8'h10 ;
			data[28778] <= 8'h10 ;
			data[28779] <= 8'h10 ;
			data[28780] <= 8'h10 ;
			data[28781] <= 8'h10 ;
			data[28782] <= 8'h10 ;
			data[28783] <= 8'h10 ;
			data[28784] <= 8'h10 ;
			data[28785] <= 8'h10 ;
			data[28786] <= 8'h10 ;
			data[28787] <= 8'h10 ;
			data[28788] <= 8'h10 ;
			data[28789] <= 8'h10 ;
			data[28790] <= 8'h10 ;
			data[28791] <= 8'h10 ;
			data[28792] <= 8'h10 ;
			data[28793] <= 8'h10 ;
			data[28794] <= 8'h10 ;
			data[28795] <= 8'h10 ;
			data[28796] <= 8'h10 ;
			data[28797] <= 8'h10 ;
			data[28798] <= 8'h10 ;
			data[28799] <= 8'h10 ;
			data[28800] <= 8'h10 ;
			data[28801] <= 8'h10 ;
			data[28802] <= 8'h10 ;
			data[28803] <= 8'h10 ;
			data[28804] <= 8'h10 ;
			data[28805] <= 8'h10 ;
			data[28806] <= 8'h10 ;
			data[28807] <= 8'h10 ;
			data[28808] <= 8'h10 ;
			data[28809] <= 8'h10 ;
			data[28810] <= 8'h10 ;
			data[28811] <= 8'h10 ;
			data[28812] <= 8'h10 ;
			data[28813] <= 8'h10 ;
			data[28814] <= 8'h10 ;
			data[28815] <= 8'h10 ;
			data[28816] <= 8'h10 ;
			data[28817] <= 8'h10 ;
			data[28818] <= 8'h10 ;
			data[28819] <= 8'h10 ;
			data[28820] <= 8'h10 ;
			data[28821] <= 8'h10 ;
			data[28822] <= 8'h10 ;
			data[28823] <= 8'h10 ;
			data[28824] <= 8'h10 ;
			data[28825] <= 8'h10 ;
			data[28826] <= 8'h10 ;
			data[28827] <= 8'h10 ;
			data[28828] <= 8'h10 ;
			data[28829] <= 8'h10 ;
			data[28830] <= 8'h10 ;
			data[28831] <= 8'h10 ;
			data[28832] <= 8'h10 ;
			data[28833] <= 8'h10 ;
			data[28834] <= 8'h10 ;
			data[28835] <= 8'h10 ;
			data[28836] <= 8'h10 ;
			data[28837] <= 8'h10 ;
			data[28838] <= 8'h10 ;
			data[28839] <= 8'h10 ;
			data[28840] <= 8'h10 ;
			data[28841] <= 8'h10 ;
			data[28842] <= 8'h10 ;
			data[28843] <= 8'h10 ;
			data[28844] <= 8'h10 ;
			data[28845] <= 8'h10 ;
			data[28846] <= 8'h10 ;
			data[28847] <= 8'h10 ;
			data[28848] <= 8'h10 ;
			data[28849] <= 8'h10 ;
			data[28850] <= 8'h10 ;
			data[28851] <= 8'h10 ;
			data[28852] <= 8'h10 ;
			data[28853] <= 8'h10 ;
			data[28854] <= 8'h10 ;
			data[28855] <= 8'h10 ;
			data[28856] <= 8'h10 ;
			data[28857] <= 8'h10 ;
			data[28858] <= 8'h10 ;
			data[28859] <= 8'h10 ;
			data[28860] <= 8'h10 ;
			data[28861] <= 8'h10 ;
			data[28862] <= 8'h10 ;
			data[28863] <= 8'h10 ;
			data[28864] <= 8'h10 ;
			data[28865] <= 8'h10 ;
			data[28866] <= 8'h10 ;
			data[28867] <= 8'h10 ;
			data[28868] <= 8'h10 ;
			data[28869] <= 8'h10 ;
			data[28870] <= 8'h10 ;
			data[28871] <= 8'h10 ;
			data[28872] <= 8'h10 ;
			data[28873] <= 8'h10 ;
			data[28874] <= 8'h10 ;
			data[28875] <= 8'h10 ;
			data[28876] <= 8'h10 ;
			data[28877] <= 8'h10 ;
			data[28878] <= 8'h10 ;
			data[28879] <= 8'h10 ;
			data[28880] <= 8'h10 ;
			data[28881] <= 8'h10 ;
			data[28882] <= 8'h10 ;
			data[28883] <= 8'h10 ;
			data[28884] <= 8'h10 ;
			data[28885] <= 8'h10 ;
			data[28886] <= 8'h10 ;
			data[28887] <= 8'h10 ;
			data[28888] <= 8'h10 ;
			data[28889] <= 8'h10 ;
			data[28890] <= 8'h10 ;
			data[28891] <= 8'h10 ;
			data[28892] <= 8'h10 ;
			data[28893] <= 8'h10 ;
			data[28894] <= 8'h10 ;
			data[28895] <= 8'h10 ;
			data[28896] <= 8'h10 ;
			data[28897] <= 8'h10 ;
			data[28898] <= 8'h10 ;
			data[28899] <= 8'h10 ;
			data[28900] <= 8'h10 ;
			data[28901] <= 8'h10 ;
			data[28902] <= 8'h10 ;
			data[28903] <= 8'h10 ;
			data[28904] <= 8'h10 ;
			data[28905] <= 8'h10 ;
			data[28906] <= 8'h10 ;
			data[28907] <= 8'h10 ;
			data[28908] <= 8'h10 ;
			data[28909] <= 8'h10 ;
			data[28910] <= 8'h10 ;
			data[28911] <= 8'h10 ;
			data[28912] <= 8'h10 ;
			data[28913] <= 8'h10 ;
			data[28914] <= 8'h10 ;
			data[28915] <= 8'h10 ;
			data[28916] <= 8'h10 ;
			data[28917] <= 8'h10 ;
			data[28918] <= 8'h10 ;
			data[28919] <= 8'h10 ;
			data[28920] <= 8'h10 ;
			data[28921] <= 8'h10 ;
			data[28922] <= 8'h10 ;
			data[28923] <= 8'h10 ;
			data[28924] <= 8'h10 ;
			data[28925] <= 8'h10 ;
			data[28926] <= 8'h10 ;
			data[28927] <= 8'h10 ;
			data[28928] <= 8'h10 ;
			data[28929] <= 8'h10 ;
			data[28930] <= 8'h10 ;
			data[28931] <= 8'h10 ;
			data[28932] <= 8'h10 ;
			data[28933] <= 8'h10 ;
			data[28934] <= 8'h10 ;
			data[28935] <= 8'h10 ;
			data[28936] <= 8'h10 ;
			data[28937] <= 8'h10 ;
			data[28938] <= 8'h10 ;
			data[28939] <= 8'h10 ;
			data[28940] <= 8'h10 ;
			data[28941] <= 8'h10 ;
			data[28942] <= 8'h10 ;
			data[28943] <= 8'h10 ;
			data[28944] <= 8'h10 ;
			data[28945] <= 8'h10 ;
			data[28946] <= 8'h10 ;
			data[28947] <= 8'h10 ;
			data[28948] <= 8'h10 ;
			data[28949] <= 8'h10 ;
			data[28950] <= 8'h10 ;
			data[28951] <= 8'h10 ;
			data[28952] <= 8'h10 ;
			data[28953] <= 8'h10 ;
			data[28954] <= 8'h10 ;
			data[28955] <= 8'h10 ;
			data[28956] <= 8'h10 ;
			data[28957] <= 8'h10 ;
			data[28958] <= 8'h10 ;
			data[28959] <= 8'h10 ;
			data[28960] <= 8'h10 ;
			data[28961] <= 8'h10 ;
			data[28962] <= 8'h10 ;
			data[28963] <= 8'h10 ;
			data[28964] <= 8'h10 ;
			data[28965] <= 8'h10 ;
			data[28966] <= 8'h10 ;
			data[28967] <= 8'h10 ;
			data[28968] <= 8'h10 ;
			data[28969] <= 8'h10 ;
			data[28970] <= 8'h10 ;
			data[28971] <= 8'h10 ;
			data[28972] <= 8'h10 ;
			data[28973] <= 8'h10 ;
			data[28974] <= 8'h10 ;
			data[28975] <= 8'h10 ;
			data[28976] <= 8'h10 ;
			data[28977] <= 8'h10 ;
			data[28978] <= 8'h10 ;
			data[28979] <= 8'h10 ;
			data[28980] <= 8'h10 ;
			data[28981] <= 8'h10 ;
			data[28982] <= 8'h10 ;
			data[28983] <= 8'h10 ;
			data[28984] <= 8'h10 ;
			data[28985] <= 8'h10 ;
			data[28986] <= 8'h10 ;
			data[28987] <= 8'h10 ;
			data[28988] <= 8'h10 ;
			data[28989] <= 8'h10 ;
			data[28990] <= 8'h10 ;
			data[28991] <= 8'h10 ;
			data[28992] <= 8'h10 ;
			data[28993] <= 8'h10 ;
			data[28994] <= 8'h10 ;
			data[28995] <= 8'h10 ;
			data[28996] <= 8'h10 ;
			data[28997] <= 8'h10 ;
			data[28998] <= 8'h10 ;
			data[28999] <= 8'h10 ;
			data[29000] <= 8'h10 ;
			data[29001] <= 8'h10 ;
			data[29002] <= 8'h10 ;
			data[29003] <= 8'h10 ;
			data[29004] <= 8'h10 ;
			data[29005] <= 8'h10 ;
			data[29006] <= 8'h10 ;
			data[29007] <= 8'h10 ;
			data[29008] <= 8'h10 ;
			data[29009] <= 8'h10 ;
			data[29010] <= 8'h10 ;
			data[29011] <= 8'h10 ;
			data[29012] <= 8'h10 ;
			data[29013] <= 8'h10 ;
			data[29014] <= 8'h10 ;
			data[29015] <= 8'h10 ;
			data[29016] <= 8'h10 ;
			data[29017] <= 8'h10 ;
			data[29018] <= 8'h10 ;
			data[29019] <= 8'h10 ;
			data[29020] <= 8'h10 ;
			data[29021] <= 8'h10 ;
			data[29022] <= 8'h10 ;
			data[29023] <= 8'h10 ;
			data[29024] <= 8'h10 ;
			data[29025] <= 8'h10 ;
			data[29026] <= 8'h10 ;
			data[29027] <= 8'h10 ;
			data[29028] <= 8'h10 ;
			data[29029] <= 8'h10 ;
			data[29030] <= 8'h10 ;
			data[29031] <= 8'h10 ;
			data[29032] <= 8'h10 ;
			data[29033] <= 8'h10 ;
			data[29034] <= 8'h10 ;
			data[29035] <= 8'h10 ;
			data[29036] <= 8'h10 ;
			data[29037] <= 8'h10 ;
			data[29038] <= 8'h10 ;
			data[29039] <= 8'h10 ;
			data[29040] <= 8'h10 ;
			data[29041] <= 8'h10 ;
			data[29042] <= 8'h10 ;
			data[29043] <= 8'h10 ;
			data[29044] <= 8'h10 ;
			data[29045] <= 8'h10 ;
			data[29046] <= 8'h10 ;
			data[29047] <= 8'h10 ;
			data[29048] <= 8'h10 ;
			data[29049] <= 8'h10 ;
			data[29050] <= 8'h10 ;
			data[29051] <= 8'h10 ;
			data[29052] <= 8'h10 ;
			data[29053] <= 8'h10 ;
			data[29054] <= 8'h10 ;
			data[29055] <= 8'h10 ;
			data[29056] <= 8'h10 ;
			data[29057] <= 8'h10 ;
			data[29058] <= 8'h10 ;
			data[29059] <= 8'h10 ;
			data[29060] <= 8'h10 ;
			data[29061] <= 8'h10 ;
			data[29062] <= 8'h10 ;
			data[29063] <= 8'h10 ;
			data[29064] <= 8'h10 ;
			data[29065] <= 8'h10 ;
			data[29066] <= 8'h10 ;
			data[29067] <= 8'h10 ;
			data[29068] <= 8'h10 ;
			data[29069] <= 8'h10 ;
			data[29070] <= 8'h10 ;
			data[29071] <= 8'h10 ;
			data[29072] <= 8'h10 ;
			data[29073] <= 8'h10 ;
			data[29074] <= 8'h10 ;
			data[29075] <= 8'h10 ;
			data[29076] <= 8'h10 ;
			data[29077] <= 8'h10 ;
			data[29078] <= 8'h10 ;
			data[29079] <= 8'h10 ;
			data[29080] <= 8'h10 ;
			data[29081] <= 8'h10 ;
			data[29082] <= 8'h10 ;
			data[29083] <= 8'h10 ;
			data[29084] <= 8'h10 ;
			data[29085] <= 8'h10 ;
			data[29086] <= 8'h10 ;
			data[29087] <= 8'h10 ;
			data[29088] <= 8'h10 ;
			data[29089] <= 8'h10 ;
			data[29090] <= 8'h10 ;
			data[29091] <= 8'h10 ;
			data[29092] <= 8'h10 ;
			data[29093] <= 8'h10 ;
			data[29094] <= 8'h10 ;
			data[29095] <= 8'h10 ;
			data[29096] <= 8'h10 ;
			data[29097] <= 8'h10 ;
			data[29098] <= 8'h10 ;
			data[29099] <= 8'h10 ;
			data[29100] <= 8'h10 ;
			data[29101] <= 8'h10 ;
			data[29102] <= 8'h10 ;
			data[29103] <= 8'h10 ;
			data[29104] <= 8'h10 ;
			data[29105] <= 8'h10 ;
			data[29106] <= 8'h10 ;
			data[29107] <= 8'h10 ;
			data[29108] <= 8'h10 ;
			data[29109] <= 8'h10 ;
			data[29110] <= 8'h10 ;
			data[29111] <= 8'h10 ;
			data[29112] <= 8'h10 ;
			data[29113] <= 8'h10 ;
			data[29114] <= 8'h10 ;
			data[29115] <= 8'h10 ;
			data[29116] <= 8'h10 ;
			data[29117] <= 8'h10 ;
			data[29118] <= 8'h10 ;
			data[29119] <= 8'h10 ;
			data[29120] <= 8'h10 ;
			data[29121] <= 8'h10 ;
			data[29122] <= 8'h10 ;
			data[29123] <= 8'h10 ;
			data[29124] <= 8'h10 ;
			data[29125] <= 8'h10 ;
			data[29126] <= 8'h10 ;
			data[29127] <= 8'h10 ;
			data[29128] <= 8'h10 ;
			data[29129] <= 8'h10 ;
			data[29130] <= 8'h10 ;
			data[29131] <= 8'h10 ;
			data[29132] <= 8'h10 ;
			data[29133] <= 8'h10 ;
			data[29134] <= 8'h10 ;
			data[29135] <= 8'h10 ;
			data[29136] <= 8'h10 ;
			data[29137] <= 8'h10 ;
			data[29138] <= 8'h10 ;
			data[29139] <= 8'h10 ;
			data[29140] <= 8'h10 ;
			data[29141] <= 8'h10 ;
			data[29142] <= 8'h10 ;
			data[29143] <= 8'h10 ;
			data[29144] <= 8'h10 ;
			data[29145] <= 8'h10 ;
			data[29146] <= 8'h10 ;
			data[29147] <= 8'h10 ;
			data[29148] <= 8'h10 ;
			data[29149] <= 8'h10 ;
			data[29150] <= 8'h10 ;
			data[29151] <= 8'h10 ;
			data[29152] <= 8'h10 ;
			data[29153] <= 8'h10 ;
			data[29154] <= 8'h10 ;
			data[29155] <= 8'h10 ;
			data[29156] <= 8'h10 ;
			data[29157] <= 8'h10 ;
			data[29158] <= 8'h10 ;
			data[29159] <= 8'h10 ;
			data[29160] <= 8'h10 ;
			data[29161] <= 8'h10 ;
			data[29162] <= 8'h10 ;
			data[29163] <= 8'h10 ;
			data[29164] <= 8'h10 ;
			data[29165] <= 8'h10 ;
			data[29166] <= 8'h10 ;
			data[29167] <= 8'h10 ;
			data[29168] <= 8'h10 ;
			data[29169] <= 8'h10 ;
			data[29170] <= 8'h10 ;
			data[29171] <= 8'h10 ;
			data[29172] <= 8'h10 ;
			data[29173] <= 8'h10 ;
			data[29174] <= 8'h10 ;
			data[29175] <= 8'h10 ;
			data[29176] <= 8'h10 ;
			data[29177] <= 8'h10 ;
			data[29178] <= 8'h10 ;
			data[29179] <= 8'h10 ;
			data[29180] <= 8'h10 ;
			data[29181] <= 8'h10 ;
			data[29182] <= 8'h10 ;
			data[29183] <= 8'h10 ;
			data[29184] <= 8'h10 ;
			data[29185] <= 8'h10 ;
			data[29186] <= 8'h10 ;
			data[29187] <= 8'h10 ;
			data[29188] <= 8'h10 ;
			data[29189] <= 8'h10 ;
			data[29190] <= 8'h10 ;
			data[29191] <= 8'h10 ;
			data[29192] <= 8'h10 ;
			data[29193] <= 8'h10 ;
			data[29194] <= 8'h10 ;
			data[29195] <= 8'h10 ;
			data[29196] <= 8'h10 ;
			data[29197] <= 8'h10 ;
			data[29198] <= 8'h10 ;
			data[29199] <= 8'h10 ;
			data[29200] <= 8'h10 ;
			data[29201] <= 8'h10 ;
			data[29202] <= 8'h10 ;
			data[29203] <= 8'h10 ;
			data[29204] <= 8'h10 ;
			data[29205] <= 8'h10 ;
			data[29206] <= 8'h10 ;
			data[29207] <= 8'h10 ;
			data[29208] <= 8'h10 ;
			data[29209] <= 8'h10 ;
			data[29210] <= 8'h10 ;
			data[29211] <= 8'h10 ;
			data[29212] <= 8'h10 ;
			data[29213] <= 8'h10 ;
			data[29214] <= 8'h10 ;
			data[29215] <= 8'h10 ;
			data[29216] <= 8'h10 ;
			data[29217] <= 8'h10 ;
			data[29218] <= 8'h10 ;
			data[29219] <= 8'h10 ;
			data[29220] <= 8'h10 ;
			data[29221] <= 8'h10 ;
			data[29222] <= 8'h10 ;
			data[29223] <= 8'h10 ;
			data[29224] <= 8'h10 ;
			data[29225] <= 8'h10 ;
			data[29226] <= 8'h10 ;
			data[29227] <= 8'h10 ;
			data[29228] <= 8'h10 ;
			data[29229] <= 8'h10 ;
			data[29230] <= 8'h10 ;
			data[29231] <= 8'h10 ;
			data[29232] <= 8'h10 ;
			data[29233] <= 8'h10 ;
			data[29234] <= 8'h10 ;
			data[29235] <= 8'h10 ;
			data[29236] <= 8'h10 ;
			data[29237] <= 8'h10 ;
			data[29238] <= 8'h10 ;
			data[29239] <= 8'h10 ;
			data[29240] <= 8'h10 ;
			data[29241] <= 8'h10 ;
			data[29242] <= 8'h10 ;
			data[29243] <= 8'h10 ;
			data[29244] <= 8'h10 ;
			data[29245] <= 8'h10 ;
			data[29246] <= 8'h10 ;
			data[29247] <= 8'h10 ;
			data[29248] <= 8'h10 ;
			data[29249] <= 8'h10 ;
			data[29250] <= 8'h10 ;
			data[29251] <= 8'h10 ;
			data[29252] <= 8'h10 ;
			data[29253] <= 8'h10 ;
			data[29254] <= 8'h10 ;
			data[29255] <= 8'h10 ;
			data[29256] <= 8'h10 ;
			data[29257] <= 8'h10 ;
			data[29258] <= 8'h10 ;
			data[29259] <= 8'h10 ;
			data[29260] <= 8'h10 ;
			data[29261] <= 8'h10 ;
			data[29262] <= 8'h10 ;
			data[29263] <= 8'h10 ;
			data[29264] <= 8'h10 ;
			data[29265] <= 8'h10 ;
			data[29266] <= 8'h10 ;
			data[29267] <= 8'h10 ;
			data[29268] <= 8'h10 ;
			data[29269] <= 8'h10 ;
			data[29270] <= 8'h10 ;
			data[29271] <= 8'h10 ;
			data[29272] <= 8'h10 ;
			data[29273] <= 8'h10 ;
			data[29274] <= 8'h10 ;
			data[29275] <= 8'h10 ;
			data[29276] <= 8'h10 ;
			data[29277] <= 8'h10 ;
			data[29278] <= 8'h10 ;
			data[29279] <= 8'h10 ;
			data[29280] <= 8'h10 ;
			data[29281] <= 8'h10 ;
			data[29282] <= 8'h10 ;
			data[29283] <= 8'h10 ;
			data[29284] <= 8'h10 ;
			data[29285] <= 8'h10 ;
			data[29286] <= 8'h10 ;
			data[29287] <= 8'h10 ;
			data[29288] <= 8'h10 ;
			data[29289] <= 8'h10 ;
			data[29290] <= 8'h10 ;
			data[29291] <= 8'h10 ;
			data[29292] <= 8'h10 ;
			data[29293] <= 8'h10 ;
			data[29294] <= 8'h10 ;
			data[29295] <= 8'h10 ;
			data[29296] <= 8'h10 ;
			data[29297] <= 8'h10 ;
			data[29298] <= 8'h10 ;
			data[29299] <= 8'h10 ;
			data[29300] <= 8'h10 ;
			data[29301] <= 8'h10 ;
			data[29302] <= 8'h10 ;
			data[29303] <= 8'h10 ;
			data[29304] <= 8'h10 ;
			data[29305] <= 8'h10 ;
			data[29306] <= 8'h10 ;
			data[29307] <= 8'h10 ;
			data[29308] <= 8'h10 ;
			data[29309] <= 8'h10 ;
			data[29310] <= 8'h10 ;
			data[29311] <= 8'h10 ;
			data[29312] <= 8'h10 ;
			data[29313] <= 8'h10 ;
			data[29314] <= 8'h10 ;
			data[29315] <= 8'h10 ;
			data[29316] <= 8'h10 ;
			data[29317] <= 8'h10 ;
			data[29318] <= 8'h10 ;
			data[29319] <= 8'h10 ;
			data[29320] <= 8'h10 ;
			data[29321] <= 8'h10 ;
			data[29322] <= 8'h10 ;
			data[29323] <= 8'h10 ;
			data[29324] <= 8'h10 ;
			data[29325] <= 8'h10 ;
			data[29326] <= 8'h10 ;
			data[29327] <= 8'h10 ;
			data[29328] <= 8'h10 ;
			data[29329] <= 8'h10 ;
			data[29330] <= 8'h10 ;
			data[29331] <= 8'h10 ;
			data[29332] <= 8'h10 ;
			data[29333] <= 8'h10 ;
			data[29334] <= 8'h10 ;
			data[29335] <= 8'h10 ;
			data[29336] <= 8'h10 ;
			data[29337] <= 8'h10 ;
			data[29338] <= 8'h10 ;
			data[29339] <= 8'h10 ;
			data[29340] <= 8'h10 ;
			data[29341] <= 8'h10 ;
			data[29342] <= 8'h10 ;
			data[29343] <= 8'h10 ;
			data[29344] <= 8'h10 ;
			data[29345] <= 8'h10 ;
			data[29346] <= 8'h10 ;
			data[29347] <= 8'h10 ;
			data[29348] <= 8'h10 ;
			data[29349] <= 8'h10 ;
			data[29350] <= 8'h10 ;
			data[29351] <= 8'h10 ;
			data[29352] <= 8'h10 ;
			data[29353] <= 8'h10 ;
			data[29354] <= 8'h10 ;
			data[29355] <= 8'h10 ;
			data[29356] <= 8'h10 ;
			data[29357] <= 8'h10 ;
			data[29358] <= 8'h10 ;
			data[29359] <= 8'h10 ;
			data[29360] <= 8'h10 ;
			data[29361] <= 8'h10 ;
			data[29362] <= 8'h10 ;
			data[29363] <= 8'h10 ;
			data[29364] <= 8'h10 ;
			data[29365] <= 8'h10 ;
			data[29366] <= 8'h10 ;
			data[29367] <= 8'h10 ;
			data[29368] <= 8'h10 ;
			data[29369] <= 8'h10 ;
			data[29370] <= 8'h10 ;
			data[29371] <= 8'h10 ;
			data[29372] <= 8'h10 ;
			data[29373] <= 8'h10 ;
			data[29374] <= 8'h10 ;
			data[29375] <= 8'h10 ;
			data[29376] <= 8'h10 ;
			data[29377] <= 8'h10 ;
			data[29378] <= 8'h10 ;
			data[29379] <= 8'h10 ;
			data[29380] <= 8'h10 ;
			data[29381] <= 8'h10 ;
			data[29382] <= 8'h10 ;
			data[29383] <= 8'h10 ;
			data[29384] <= 8'h10 ;
			data[29385] <= 8'h10 ;
			data[29386] <= 8'h10 ;
			data[29387] <= 8'h10 ;
			data[29388] <= 8'h10 ;
			data[29389] <= 8'h10 ;
			data[29390] <= 8'h10 ;
			data[29391] <= 8'h10 ;
			data[29392] <= 8'h10 ;
			data[29393] <= 8'h10 ;
			data[29394] <= 8'h10 ;
			data[29395] <= 8'h10 ;
			data[29396] <= 8'h10 ;
			data[29397] <= 8'h10 ;
			data[29398] <= 8'h10 ;
			data[29399] <= 8'h10 ;
			data[29400] <= 8'h10 ;
			data[29401] <= 8'h10 ;
			data[29402] <= 8'h10 ;
			data[29403] <= 8'h10 ;
			data[29404] <= 8'h10 ;
			data[29405] <= 8'h10 ;
			data[29406] <= 8'h10 ;
			data[29407] <= 8'h10 ;
			data[29408] <= 8'h10 ;
			data[29409] <= 8'h10 ;
			data[29410] <= 8'h10 ;
			data[29411] <= 8'h10 ;
			data[29412] <= 8'h10 ;
			data[29413] <= 8'h10 ;
			data[29414] <= 8'h10 ;
			data[29415] <= 8'h10 ;
			data[29416] <= 8'h10 ;
			data[29417] <= 8'h10 ;
			data[29418] <= 8'h10 ;
			data[29419] <= 8'h10 ;
			data[29420] <= 8'h10 ;
			data[29421] <= 8'h10 ;
			data[29422] <= 8'h10 ;
			data[29423] <= 8'h10 ;
			data[29424] <= 8'h10 ;
			data[29425] <= 8'h10 ;
			data[29426] <= 8'h10 ;
			data[29427] <= 8'h10 ;
			data[29428] <= 8'h10 ;
			data[29429] <= 8'h10 ;
			data[29430] <= 8'h10 ;
			data[29431] <= 8'h10 ;
			data[29432] <= 8'h10 ;
			data[29433] <= 8'h10 ;
			data[29434] <= 8'h10 ;
			data[29435] <= 8'h10 ;
			data[29436] <= 8'h10 ;
			data[29437] <= 8'h10 ;
			data[29438] <= 8'h10 ;
			data[29439] <= 8'h10 ;
			data[29440] <= 8'h10 ;
			data[29441] <= 8'h10 ;
			data[29442] <= 8'h10 ;
			data[29443] <= 8'h10 ;
			data[29444] <= 8'h10 ;
			data[29445] <= 8'h10 ;
			data[29446] <= 8'h10 ;
			data[29447] <= 8'h10 ;
			data[29448] <= 8'h10 ;
			data[29449] <= 8'h10 ;
			data[29450] <= 8'h10 ;
			data[29451] <= 8'h10 ;
			data[29452] <= 8'h10 ;
			data[29453] <= 8'h10 ;
			data[29454] <= 8'h10 ;
			data[29455] <= 8'h10 ;
			data[29456] <= 8'h10 ;
			data[29457] <= 8'h10 ;
			data[29458] <= 8'h10 ;
			data[29459] <= 8'h10 ;
			data[29460] <= 8'h10 ;
			data[29461] <= 8'h10 ;
			data[29462] <= 8'h10 ;
			data[29463] <= 8'h10 ;
			data[29464] <= 8'h10 ;
			data[29465] <= 8'h10 ;
			data[29466] <= 8'h10 ;
			data[29467] <= 8'h10 ;
			data[29468] <= 8'h10 ;
			data[29469] <= 8'h10 ;
			data[29470] <= 8'h10 ;
			data[29471] <= 8'h10 ;
			data[29472] <= 8'h10 ;
			data[29473] <= 8'h10 ;
			data[29474] <= 8'h10 ;
			data[29475] <= 8'h10 ;
			data[29476] <= 8'h10 ;
			data[29477] <= 8'h10 ;
			data[29478] <= 8'h10 ;
			data[29479] <= 8'h10 ;
			data[29480] <= 8'h10 ;
			data[29481] <= 8'h10 ;
			data[29482] <= 8'h10 ;
			data[29483] <= 8'h10 ;
			data[29484] <= 8'h10 ;
			data[29485] <= 8'h10 ;
			data[29486] <= 8'h10 ;
			data[29487] <= 8'h10 ;
			data[29488] <= 8'h10 ;
			data[29489] <= 8'h10 ;
			data[29490] <= 8'h10 ;
			data[29491] <= 8'h10 ;
			data[29492] <= 8'h10 ;
			data[29493] <= 8'h10 ;
			data[29494] <= 8'h10 ;
			data[29495] <= 8'h10 ;
			data[29496] <= 8'h10 ;
			data[29497] <= 8'h10 ;
			data[29498] <= 8'h10 ;
			data[29499] <= 8'h10 ;
			data[29500] <= 8'h10 ;
			data[29501] <= 8'h10 ;
			data[29502] <= 8'h10 ;
			data[29503] <= 8'h10 ;
			data[29504] <= 8'h10 ;
			data[29505] <= 8'h10 ;
			data[29506] <= 8'h10 ;
			data[29507] <= 8'h10 ;
			data[29508] <= 8'h10 ;
			data[29509] <= 8'h10 ;
			data[29510] <= 8'h10 ;
			data[29511] <= 8'h10 ;
			data[29512] <= 8'h10 ;
			data[29513] <= 8'h10 ;
			data[29514] <= 8'h10 ;
			data[29515] <= 8'h10 ;
			data[29516] <= 8'h10 ;
			data[29517] <= 8'h10 ;
			data[29518] <= 8'h10 ;
			data[29519] <= 8'h10 ;
			data[29520] <= 8'h10 ;
			data[29521] <= 8'h10 ;
			data[29522] <= 8'h10 ;
			data[29523] <= 8'h10 ;
			data[29524] <= 8'h10 ;
			data[29525] <= 8'h10 ;
			data[29526] <= 8'h10 ;
			data[29527] <= 8'h10 ;
			data[29528] <= 8'h10 ;
			data[29529] <= 8'h10 ;
			data[29530] <= 8'h10 ;
			data[29531] <= 8'h10 ;
			data[29532] <= 8'h10 ;
			data[29533] <= 8'h10 ;
			data[29534] <= 8'h10 ;
			data[29535] <= 8'h10 ;
			data[29536] <= 8'h10 ;
			data[29537] <= 8'h10 ;
			data[29538] <= 8'h10 ;
			data[29539] <= 8'h10 ;
			data[29540] <= 8'h10 ;
			data[29541] <= 8'h10 ;
			data[29542] <= 8'h10 ;
			data[29543] <= 8'h10 ;
			data[29544] <= 8'h10 ;
			data[29545] <= 8'h10 ;
			data[29546] <= 8'h10 ;
			data[29547] <= 8'h10 ;
			data[29548] <= 8'h10 ;
			data[29549] <= 8'h10 ;
			data[29550] <= 8'h10 ;
			data[29551] <= 8'h10 ;
			data[29552] <= 8'h10 ;
			data[29553] <= 8'h10 ;
			data[29554] <= 8'h10 ;
			data[29555] <= 8'h10 ;
			data[29556] <= 8'h10 ;
			data[29557] <= 8'h10 ;
			data[29558] <= 8'h10 ;
			data[29559] <= 8'h10 ;
			data[29560] <= 8'h10 ;
			data[29561] <= 8'h10 ;
			data[29562] <= 8'h10 ;
			data[29563] <= 8'h10 ;
			data[29564] <= 8'h10 ;
			data[29565] <= 8'h10 ;
			data[29566] <= 8'h10 ;
			data[29567] <= 8'h10 ;
			data[29568] <= 8'h10 ;
			data[29569] <= 8'h10 ;
			data[29570] <= 8'h10 ;
			data[29571] <= 8'h10 ;
			data[29572] <= 8'h10 ;
			data[29573] <= 8'h10 ;
			data[29574] <= 8'h10 ;
			data[29575] <= 8'h10 ;
			data[29576] <= 8'h10 ;
			data[29577] <= 8'h10 ;
			data[29578] <= 8'h10 ;
			data[29579] <= 8'h10 ;
			data[29580] <= 8'h10 ;
			data[29581] <= 8'h10 ;
			data[29582] <= 8'h10 ;
			data[29583] <= 8'h10 ;
			data[29584] <= 8'h10 ;
			data[29585] <= 8'h10 ;
			data[29586] <= 8'h10 ;
			data[29587] <= 8'h10 ;
			data[29588] <= 8'h10 ;
			data[29589] <= 8'h10 ;
			data[29590] <= 8'h10 ;
			data[29591] <= 8'h10 ;
			data[29592] <= 8'h10 ;
			data[29593] <= 8'h10 ;
			data[29594] <= 8'h10 ;
			data[29595] <= 8'h10 ;
			data[29596] <= 8'h10 ;
			data[29597] <= 8'h10 ;
			data[29598] <= 8'h10 ;
			data[29599] <= 8'h10 ;
			data[29600] <= 8'h10 ;
			data[29601] <= 8'h10 ;
			data[29602] <= 8'h10 ;
			data[29603] <= 8'h10 ;
			data[29604] <= 8'h10 ;
			data[29605] <= 8'h10 ;
			data[29606] <= 8'h10 ;
			data[29607] <= 8'h10 ;
			data[29608] <= 8'h10 ;
			data[29609] <= 8'h10 ;
			data[29610] <= 8'h10 ;
			data[29611] <= 8'h10 ;
			data[29612] <= 8'h10 ;
			data[29613] <= 8'h10 ;
			data[29614] <= 8'h10 ;
			data[29615] <= 8'h10 ;
			data[29616] <= 8'h10 ;
			data[29617] <= 8'h10 ;
			data[29618] <= 8'h10 ;
			data[29619] <= 8'h10 ;
			data[29620] <= 8'h10 ;
			data[29621] <= 8'h10 ;
			data[29622] <= 8'h10 ;
			data[29623] <= 8'h10 ;
			data[29624] <= 8'h10 ;
			data[29625] <= 8'h10 ;
			data[29626] <= 8'h10 ;
			data[29627] <= 8'h10 ;
			data[29628] <= 8'h10 ;
			data[29629] <= 8'h10 ;
			data[29630] <= 8'h10 ;
			data[29631] <= 8'h10 ;
			data[29632] <= 8'h10 ;
			data[29633] <= 8'h10 ;
			data[29634] <= 8'h10 ;
			data[29635] <= 8'h10 ;
			data[29636] <= 8'h10 ;
			data[29637] <= 8'h10 ;
			data[29638] <= 8'h10 ;
			data[29639] <= 8'h10 ;
			data[29640] <= 8'h10 ;
			data[29641] <= 8'h10 ;
			data[29642] <= 8'h10 ;
			data[29643] <= 8'h10 ;
			data[29644] <= 8'h10 ;
			data[29645] <= 8'h10 ;
			data[29646] <= 8'h10 ;
			data[29647] <= 8'h10 ;
			data[29648] <= 8'h10 ;
			data[29649] <= 8'h10 ;
			data[29650] <= 8'h10 ;
			data[29651] <= 8'h10 ;
			data[29652] <= 8'h10 ;
			data[29653] <= 8'h10 ;
			data[29654] <= 8'h10 ;
			data[29655] <= 8'h10 ;
			data[29656] <= 8'h10 ;
			data[29657] <= 8'h10 ;
			data[29658] <= 8'h10 ;
			data[29659] <= 8'h10 ;
			data[29660] <= 8'h10 ;
			data[29661] <= 8'h10 ;
			data[29662] <= 8'h10 ;
			data[29663] <= 8'h10 ;
			data[29664] <= 8'h10 ;
			data[29665] <= 8'h10 ;
			data[29666] <= 8'h10 ;
			data[29667] <= 8'h10 ;
			data[29668] <= 8'h10 ;
			data[29669] <= 8'h10 ;
			data[29670] <= 8'h10 ;
			data[29671] <= 8'h10 ;
			data[29672] <= 8'h10 ;
			data[29673] <= 8'h10 ;
			data[29674] <= 8'h10 ;
			data[29675] <= 8'h10 ;
			data[29676] <= 8'h10 ;
			data[29677] <= 8'h10 ;
			data[29678] <= 8'h10 ;
			data[29679] <= 8'h10 ;
			data[29680] <= 8'h10 ;
			data[29681] <= 8'h10 ;
			data[29682] <= 8'h10 ;
			data[29683] <= 8'h10 ;
			data[29684] <= 8'h10 ;
			data[29685] <= 8'h10 ;
			data[29686] <= 8'h10 ;
			data[29687] <= 8'h10 ;
			data[29688] <= 8'h10 ;
			data[29689] <= 8'h10 ;
			data[29690] <= 8'h10 ;
			data[29691] <= 8'h10 ;
			data[29692] <= 8'h10 ;
			data[29693] <= 8'h10 ;
			data[29694] <= 8'h10 ;
			data[29695] <= 8'h10 ;
			data[29696] <= 8'h10 ;
			data[29697] <= 8'h10 ;
			data[29698] <= 8'h10 ;
			data[29699] <= 8'h10 ;
			data[29700] <= 8'h10 ;
			data[29701] <= 8'h10 ;
			data[29702] <= 8'h10 ;
			data[29703] <= 8'h10 ;
			data[29704] <= 8'h10 ;
			data[29705] <= 8'h10 ;
			data[29706] <= 8'h10 ;
			data[29707] <= 8'h10 ;
			data[29708] <= 8'h10 ;
			data[29709] <= 8'h10 ;
			data[29710] <= 8'h10 ;
			data[29711] <= 8'h10 ;
			data[29712] <= 8'h10 ;
			data[29713] <= 8'h10 ;
			data[29714] <= 8'h10 ;
			data[29715] <= 8'h10 ;
			data[29716] <= 8'h10 ;
			data[29717] <= 8'h10 ;
			data[29718] <= 8'h10 ;
			data[29719] <= 8'h10 ;
			data[29720] <= 8'h10 ;
			data[29721] <= 8'h10 ;
			data[29722] <= 8'h10 ;
			data[29723] <= 8'h10 ;
			data[29724] <= 8'h10 ;
			data[29725] <= 8'h10 ;
			data[29726] <= 8'h10 ;
			data[29727] <= 8'h10 ;
			data[29728] <= 8'h10 ;
			data[29729] <= 8'h10 ;
			data[29730] <= 8'h10 ;
			data[29731] <= 8'h10 ;
			data[29732] <= 8'h10 ;
			data[29733] <= 8'h10 ;
			data[29734] <= 8'h10 ;
			data[29735] <= 8'h10 ;
			data[29736] <= 8'h10 ;
			data[29737] <= 8'h10 ;
			data[29738] <= 8'h10 ;
			data[29739] <= 8'h10 ;
			data[29740] <= 8'h10 ;
			data[29741] <= 8'h10 ;
			data[29742] <= 8'h10 ;
			data[29743] <= 8'h10 ;
			data[29744] <= 8'h10 ;
			data[29745] <= 8'h10 ;
			data[29746] <= 8'h10 ;
			data[29747] <= 8'h10 ;
			data[29748] <= 8'h10 ;
			data[29749] <= 8'h10 ;
			data[29750] <= 8'h10 ;
			data[29751] <= 8'h10 ;
			data[29752] <= 8'h10 ;
			data[29753] <= 8'h10 ;
			data[29754] <= 8'h10 ;
			data[29755] <= 8'h10 ;
			data[29756] <= 8'h10 ;
			data[29757] <= 8'h10 ;
			data[29758] <= 8'h10 ;
			data[29759] <= 8'h10 ;
			data[29760] <= 8'h10 ;
			data[29761] <= 8'h10 ;
			data[29762] <= 8'h10 ;
			data[29763] <= 8'h10 ;
			data[29764] <= 8'h10 ;
			data[29765] <= 8'h10 ;
			data[29766] <= 8'h10 ;
			data[29767] <= 8'h10 ;
			data[29768] <= 8'h10 ;
			data[29769] <= 8'h10 ;
			data[29770] <= 8'h10 ;
			data[29771] <= 8'h10 ;
			data[29772] <= 8'h10 ;
			data[29773] <= 8'h10 ;
			data[29774] <= 8'h10 ;
			data[29775] <= 8'h10 ;
			data[29776] <= 8'h10 ;
			data[29777] <= 8'h10 ;
			data[29778] <= 8'h10 ;
			data[29779] <= 8'h10 ;
			data[29780] <= 8'h10 ;
			data[29781] <= 8'h10 ;
			data[29782] <= 8'h10 ;
			data[29783] <= 8'h10 ;
			data[29784] <= 8'h10 ;
			data[29785] <= 8'h10 ;
			data[29786] <= 8'h10 ;
			data[29787] <= 8'h10 ;
			data[29788] <= 8'h10 ;
			data[29789] <= 8'h10 ;
			data[29790] <= 8'h10 ;
			data[29791] <= 8'h10 ;
			data[29792] <= 8'h10 ;
			data[29793] <= 8'h10 ;
			data[29794] <= 8'h10 ;
			data[29795] <= 8'h10 ;
			data[29796] <= 8'h10 ;
			data[29797] <= 8'h10 ;
			data[29798] <= 8'h10 ;
			data[29799] <= 8'h10 ;
			data[29800] <= 8'h10 ;
			data[29801] <= 8'h10 ;
			data[29802] <= 8'h10 ;
			data[29803] <= 8'h10 ;
			data[29804] <= 8'h10 ;
			data[29805] <= 8'h10 ;
			data[29806] <= 8'h10 ;
			data[29807] <= 8'h10 ;
			data[29808] <= 8'h10 ;
			data[29809] <= 8'h10 ;
			data[29810] <= 8'h10 ;
			data[29811] <= 8'h10 ;
			data[29812] <= 8'h10 ;
			data[29813] <= 8'h10 ;
			data[29814] <= 8'h10 ;
			data[29815] <= 8'h10 ;
			data[29816] <= 8'h10 ;
			data[29817] <= 8'h10 ;
			data[29818] <= 8'h10 ;
			data[29819] <= 8'h10 ;
			data[29820] <= 8'h10 ;
			data[29821] <= 8'h10 ;
			data[29822] <= 8'h10 ;
			data[29823] <= 8'h10 ;
			data[29824] <= 8'h10 ;
			data[29825] <= 8'h10 ;
			data[29826] <= 8'h10 ;
			data[29827] <= 8'h10 ;
			data[29828] <= 8'h10 ;
			data[29829] <= 8'h10 ;
			data[29830] <= 8'h10 ;
			data[29831] <= 8'h10 ;
			data[29832] <= 8'h10 ;
			data[29833] <= 8'h10 ;
			data[29834] <= 8'h10 ;
			data[29835] <= 8'h10 ;
			data[29836] <= 8'h10 ;
			data[29837] <= 8'h10 ;
			data[29838] <= 8'h10 ;
			data[29839] <= 8'h10 ;
			data[29840] <= 8'h10 ;
			data[29841] <= 8'h10 ;
			data[29842] <= 8'h10 ;
			data[29843] <= 8'h10 ;
			data[29844] <= 8'h10 ;
			data[29845] <= 8'h10 ;
			data[29846] <= 8'h10 ;
			data[29847] <= 8'h10 ;
			data[29848] <= 8'h10 ;
			data[29849] <= 8'h10 ;
			data[29850] <= 8'h10 ;
			data[29851] <= 8'h10 ;
			data[29852] <= 8'h10 ;
			data[29853] <= 8'h10 ;
			data[29854] <= 8'h10 ;
			data[29855] <= 8'h10 ;
			data[29856] <= 8'h10 ;
			data[29857] <= 8'h10 ;
			data[29858] <= 8'h10 ;
			data[29859] <= 8'h10 ;
			data[29860] <= 8'h10 ;
			data[29861] <= 8'h10 ;
			data[29862] <= 8'h10 ;
			data[29863] <= 8'h10 ;
			data[29864] <= 8'h10 ;
			data[29865] <= 8'h10 ;
			data[29866] <= 8'h10 ;
			data[29867] <= 8'h10 ;
			data[29868] <= 8'h10 ;
			data[29869] <= 8'h10 ;
			data[29870] <= 8'h10 ;
			data[29871] <= 8'h10 ;
			data[29872] <= 8'h10 ;
			data[29873] <= 8'h10 ;
			data[29874] <= 8'h10 ;
			data[29875] <= 8'h10 ;
			data[29876] <= 8'h10 ;
			data[29877] <= 8'h10 ;
			data[29878] <= 8'h10 ;
			data[29879] <= 8'h10 ;
			data[29880] <= 8'h10 ;
			data[29881] <= 8'h10 ;
			data[29882] <= 8'h10 ;
			data[29883] <= 8'h10 ;
			data[29884] <= 8'h10 ;
			data[29885] <= 8'h10 ;
			data[29886] <= 8'h10 ;
			data[29887] <= 8'h10 ;
			data[29888] <= 8'h10 ;
			data[29889] <= 8'h10 ;
			data[29890] <= 8'h10 ;
			data[29891] <= 8'h10 ;
			data[29892] <= 8'h10 ;
			data[29893] <= 8'h10 ;
			data[29894] <= 8'h10 ;
			data[29895] <= 8'h10 ;
			data[29896] <= 8'h10 ;
			data[29897] <= 8'h10 ;
			data[29898] <= 8'h10 ;
			data[29899] <= 8'h10 ;
			data[29900] <= 8'h10 ;
			data[29901] <= 8'h10 ;
			data[29902] <= 8'h10 ;
			data[29903] <= 8'h10 ;
			data[29904] <= 8'h10 ;
			data[29905] <= 8'h10 ;
			data[29906] <= 8'h10 ;
			data[29907] <= 8'h10 ;
			data[29908] <= 8'h10 ;
			data[29909] <= 8'h10 ;
			data[29910] <= 8'h10 ;
			data[29911] <= 8'h10 ;
			data[29912] <= 8'h10 ;
			data[29913] <= 8'h10 ;
			data[29914] <= 8'h10 ;
			data[29915] <= 8'h10 ;
			data[29916] <= 8'h10 ;
			data[29917] <= 8'h10 ;
			data[29918] <= 8'h10 ;
			data[29919] <= 8'h10 ;
			data[29920] <= 8'h10 ;
			data[29921] <= 8'h10 ;
			data[29922] <= 8'h10 ;
			data[29923] <= 8'h10 ;
			data[29924] <= 8'h10 ;
			data[29925] <= 8'h10 ;
			data[29926] <= 8'h10 ;
			data[29927] <= 8'h10 ;
			data[29928] <= 8'h10 ;
			data[29929] <= 8'h10 ;
			data[29930] <= 8'h10 ;
			data[29931] <= 8'h10 ;
			data[29932] <= 8'h10 ;
			data[29933] <= 8'h10 ;
			data[29934] <= 8'h10 ;
			data[29935] <= 8'h10 ;
			data[29936] <= 8'h10 ;
			data[29937] <= 8'h10 ;
			data[29938] <= 8'h10 ;
			data[29939] <= 8'h10 ;
			data[29940] <= 8'h10 ;
			data[29941] <= 8'h10 ;
			data[29942] <= 8'h10 ;
			data[29943] <= 8'h10 ;
			data[29944] <= 8'h10 ;
			data[29945] <= 8'h10 ;
			data[29946] <= 8'h10 ;
			data[29947] <= 8'h10 ;
			data[29948] <= 8'h10 ;
			data[29949] <= 8'h10 ;
			data[29950] <= 8'h10 ;
			data[29951] <= 8'h10 ;
			data[29952] <= 8'h10 ;
			data[29953] <= 8'h10 ;
			data[29954] <= 8'h10 ;
			data[29955] <= 8'h10 ;
			data[29956] <= 8'h10 ;
			data[29957] <= 8'h10 ;
			data[29958] <= 8'h10 ;
			data[29959] <= 8'h10 ;
			data[29960] <= 8'h10 ;
			data[29961] <= 8'h10 ;
			data[29962] <= 8'h10 ;
			data[29963] <= 8'h10 ;
			data[29964] <= 8'h10 ;
			data[29965] <= 8'h10 ;
			data[29966] <= 8'h10 ;
			data[29967] <= 8'h10 ;
			data[29968] <= 8'h10 ;
			data[29969] <= 8'h10 ;
			data[29970] <= 8'h10 ;
			data[29971] <= 8'h10 ;
			data[29972] <= 8'h10 ;
			data[29973] <= 8'h10 ;
			data[29974] <= 8'h10 ;
			data[29975] <= 8'h10 ;
			data[29976] <= 8'h10 ;
			data[29977] <= 8'h10 ;
			data[29978] <= 8'h10 ;
			data[29979] <= 8'h10 ;
			data[29980] <= 8'h10 ;
			data[29981] <= 8'h10 ;
			data[29982] <= 8'h10 ;
			data[29983] <= 8'h10 ;
			data[29984] <= 8'h10 ;
			data[29985] <= 8'h10 ;
			data[29986] <= 8'h10 ;
			data[29987] <= 8'h10 ;
			data[29988] <= 8'h10 ;
			data[29989] <= 8'h10 ;
			data[29990] <= 8'h10 ;
			data[29991] <= 8'h10 ;
			data[29992] <= 8'h10 ;
			data[29993] <= 8'h10 ;
			data[29994] <= 8'h10 ;
			data[29995] <= 8'h10 ;
			data[29996] <= 8'h10 ;
			data[29997] <= 8'h10 ;
			data[29998] <= 8'h10 ;
			data[29999] <= 8'h10 ;
			data[30000] <= 8'h10 ;
			data[30001] <= 8'h10 ;
			data[30002] <= 8'h10 ;
			data[30003] <= 8'h10 ;
			data[30004] <= 8'h10 ;
			data[30005] <= 8'h10 ;
			data[30006] <= 8'h10 ;
			data[30007] <= 8'h10 ;
			data[30008] <= 8'h10 ;
			data[30009] <= 8'h10 ;
			data[30010] <= 8'h10 ;
			data[30011] <= 8'h10 ;
			data[30012] <= 8'h10 ;
			data[30013] <= 8'h10 ;
			data[30014] <= 8'h10 ;
			data[30015] <= 8'h10 ;
			data[30016] <= 8'h10 ;
			data[30017] <= 8'h10 ;
			data[30018] <= 8'h10 ;
			data[30019] <= 8'h10 ;
			data[30020] <= 8'h10 ;
			data[30021] <= 8'h10 ;
			data[30022] <= 8'h10 ;
			data[30023] <= 8'h10 ;
			data[30024] <= 8'h10 ;
			data[30025] <= 8'h10 ;
			data[30026] <= 8'h10 ;
			data[30027] <= 8'h10 ;
			data[30028] <= 8'h10 ;
			data[30029] <= 8'h10 ;
			data[30030] <= 8'h10 ;
			data[30031] <= 8'h10 ;
			data[30032] <= 8'h10 ;
			data[30033] <= 8'h10 ;
			data[30034] <= 8'h10 ;
			data[30035] <= 8'h10 ;
			data[30036] <= 8'h10 ;
			data[30037] <= 8'h10 ;
			data[30038] <= 8'h10 ;
			data[30039] <= 8'h10 ;
			data[30040] <= 8'h10 ;
			data[30041] <= 8'h10 ;
			data[30042] <= 8'h10 ;
			data[30043] <= 8'h10 ;
			data[30044] <= 8'h10 ;
			data[30045] <= 8'h10 ;
			data[30046] <= 8'h10 ;
			data[30047] <= 8'h10 ;
			data[30048] <= 8'h10 ;
			data[30049] <= 8'h10 ;
			data[30050] <= 8'h10 ;
			data[30051] <= 8'h10 ;
			data[30052] <= 8'h10 ;
			data[30053] <= 8'h10 ;
			data[30054] <= 8'h10 ;
			data[30055] <= 8'h10 ;
			data[30056] <= 8'h10 ;
			data[30057] <= 8'h10 ;
			data[30058] <= 8'h10 ;
			data[30059] <= 8'h10 ;
			data[30060] <= 8'h10 ;
			data[30061] <= 8'h10 ;
			data[30062] <= 8'h10 ;
			data[30063] <= 8'h10 ;
			data[30064] <= 8'h10 ;
			data[30065] <= 8'h10 ;
			data[30066] <= 8'h10 ;
			data[30067] <= 8'h10 ;
			data[30068] <= 8'h10 ;
			data[30069] <= 8'h10 ;
			data[30070] <= 8'h10 ;
			data[30071] <= 8'h10 ;
			data[30072] <= 8'h10 ;
			data[30073] <= 8'h10 ;
			data[30074] <= 8'h10 ;
			data[30075] <= 8'h10 ;
			data[30076] <= 8'h10 ;
			data[30077] <= 8'h10 ;
			data[30078] <= 8'h10 ;
			data[30079] <= 8'h10 ;
			data[30080] <= 8'h10 ;
			data[30081] <= 8'h10 ;
			data[30082] <= 8'h10 ;
			data[30083] <= 8'h10 ;
			data[30084] <= 8'h10 ;
			data[30085] <= 8'h10 ;
			data[30086] <= 8'h10 ;
			data[30087] <= 8'h10 ;
			data[30088] <= 8'h10 ;
			data[30089] <= 8'h10 ;
			data[30090] <= 8'h10 ;
			data[30091] <= 8'h10 ;
			data[30092] <= 8'h10 ;
			data[30093] <= 8'h10 ;
			data[30094] <= 8'h10 ;
			data[30095] <= 8'h10 ;
			data[30096] <= 8'h10 ;
			data[30097] <= 8'h10 ;
			data[30098] <= 8'h10 ;
			data[30099] <= 8'h10 ;
			data[30100] <= 8'h10 ;
			data[30101] <= 8'h10 ;
			data[30102] <= 8'h10 ;
			data[30103] <= 8'h10 ;
			data[30104] <= 8'h10 ;
			data[30105] <= 8'h10 ;
			data[30106] <= 8'h10 ;
			data[30107] <= 8'h10 ;
			data[30108] <= 8'h10 ;
			data[30109] <= 8'h10 ;
			data[30110] <= 8'h10 ;
			data[30111] <= 8'h10 ;
			data[30112] <= 8'h10 ;
			data[30113] <= 8'h10 ;
			data[30114] <= 8'h10 ;
			data[30115] <= 8'h10 ;
			data[30116] <= 8'h10 ;
			data[30117] <= 8'h10 ;
			data[30118] <= 8'h10 ;
			data[30119] <= 8'h10 ;
			data[30120] <= 8'h10 ;
			data[30121] <= 8'h10 ;
			data[30122] <= 8'h10 ;
			data[30123] <= 8'h10 ;
			data[30124] <= 8'h10 ;
			data[30125] <= 8'h10 ;
			data[30126] <= 8'h10 ;
			data[30127] <= 8'h10 ;
			data[30128] <= 8'h10 ;
			data[30129] <= 8'h10 ;
			data[30130] <= 8'h10 ;
			data[30131] <= 8'h10 ;
			data[30132] <= 8'h10 ;
			data[30133] <= 8'h10 ;
			data[30134] <= 8'h10 ;
			data[30135] <= 8'h10 ;
			data[30136] <= 8'h10 ;
			data[30137] <= 8'h10 ;
			data[30138] <= 8'h10 ;
			data[30139] <= 8'h10 ;
			data[30140] <= 8'h10 ;
			data[30141] <= 8'h10 ;
			data[30142] <= 8'h10 ;
			data[30143] <= 8'h10 ;
			data[30144] <= 8'h10 ;
			data[30145] <= 8'h10 ;
			data[30146] <= 8'h10 ;
			data[30147] <= 8'h10 ;
			data[30148] <= 8'h10 ;
			data[30149] <= 8'h10 ;
			data[30150] <= 8'h10 ;
			data[30151] <= 8'h10 ;
			data[30152] <= 8'h10 ;
			data[30153] <= 8'h10 ;
			data[30154] <= 8'h10 ;
			data[30155] <= 8'h10 ;
			data[30156] <= 8'h10 ;
			data[30157] <= 8'h10 ;
			data[30158] <= 8'h10 ;
			data[30159] <= 8'h10 ;
			data[30160] <= 8'h10 ;
			data[30161] <= 8'h10 ;
			data[30162] <= 8'h10 ;
			data[30163] <= 8'h10 ;
			data[30164] <= 8'h10 ;
			data[30165] <= 8'h10 ;
			data[30166] <= 8'h10 ;
			data[30167] <= 8'h10 ;
			data[30168] <= 8'h10 ;
			data[30169] <= 8'h10 ;
			data[30170] <= 8'h10 ;
			data[30171] <= 8'h10 ;
			data[30172] <= 8'h10 ;
			data[30173] <= 8'h10 ;
			data[30174] <= 8'h10 ;
			data[30175] <= 8'h10 ;
			data[30176] <= 8'h10 ;
			data[30177] <= 8'h10 ;
			data[30178] <= 8'h10 ;
			data[30179] <= 8'h10 ;
			data[30180] <= 8'h10 ;
			data[30181] <= 8'h10 ;
			data[30182] <= 8'h10 ;
			data[30183] <= 8'h10 ;
			data[30184] <= 8'h10 ;
			data[30185] <= 8'h10 ;
			data[30186] <= 8'h10 ;
			data[30187] <= 8'h10 ;
			data[30188] <= 8'h10 ;
			data[30189] <= 8'h10 ;
			data[30190] <= 8'h10 ;
			data[30191] <= 8'h10 ;
			data[30192] <= 8'h10 ;
			data[30193] <= 8'h10 ;
			data[30194] <= 8'h10 ;
			data[30195] <= 8'h10 ;
			data[30196] <= 8'h10 ;
			data[30197] <= 8'h10 ;
			data[30198] <= 8'h10 ;
			data[30199] <= 8'h10 ;
			data[30200] <= 8'h10 ;
			data[30201] <= 8'h10 ;
			data[30202] <= 8'h10 ;
			data[30203] <= 8'h10 ;
			data[30204] <= 8'h10 ;
			data[30205] <= 8'h10 ;
			data[30206] <= 8'h10 ;
			data[30207] <= 8'h10 ;
			data[30208] <= 8'h10 ;
			data[30209] <= 8'h10 ;
			data[30210] <= 8'h10 ;
			data[30211] <= 8'h10 ;
			data[30212] <= 8'h10 ;
			data[30213] <= 8'h10 ;
			data[30214] <= 8'h10 ;
			data[30215] <= 8'h10 ;
			data[30216] <= 8'h10 ;
			data[30217] <= 8'h10 ;
			data[30218] <= 8'h10 ;
			data[30219] <= 8'h10 ;
			data[30220] <= 8'h10 ;
			data[30221] <= 8'h10 ;
			data[30222] <= 8'h10 ;
			data[30223] <= 8'h10 ;
			data[30224] <= 8'h10 ;
			data[30225] <= 8'h10 ;
			data[30226] <= 8'h10 ;
			data[30227] <= 8'h10 ;
			data[30228] <= 8'h10 ;
			data[30229] <= 8'h10 ;
			data[30230] <= 8'h10 ;
			data[30231] <= 8'h10 ;
			data[30232] <= 8'h10 ;
			data[30233] <= 8'h10 ;
			data[30234] <= 8'h10 ;
			data[30235] <= 8'h10 ;
			data[30236] <= 8'h10 ;
			data[30237] <= 8'h10 ;
			data[30238] <= 8'h10 ;
			data[30239] <= 8'h10 ;
			data[30240] <= 8'h10 ;
			data[30241] <= 8'h10 ;
			data[30242] <= 8'h10 ;
			data[30243] <= 8'h10 ;
			data[30244] <= 8'h10 ;
			data[30245] <= 8'h10 ;
			data[30246] <= 8'h10 ;
			data[30247] <= 8'h10 ;
			data[30248] <= 8'h10 ;
			data[30249] <= 8'h10 ;
			data[30250] <= 8'h10 ;
			data[30251] <= 8'h10 ;
			data[30252] <= 8'h10 ;
			data[30253] <= 8'h10 ;
			data[30254] <= 8'h10 ;
			data[30255] <= 8'h10 ;
			data[30256] <= 8'h10 ;
			data[30257] <= 8'h10 ;
			data[30258] <= 8'h10 ;
			data[30259] <= 8'h10 ;
			data[30260] <= 8'h10 ;
			data[30261] <= 8'h10 ;
			data[30262] <= 8'h10 ;
			data[30263] <= 8'h10 ;
			data[30264] <= 8'h10 ;
			data[30265] <= 8'h10 ;
			data[30266] <= 8'h10 ;
			data[30267] <= 8'h10 ;
			data[30268] <= 8'h10 ;
			data[30269] <= 8'h10 ;
			data[30270] <= 8'h10 ;
			data[30271] <= 8'h10 ;
			data[30272] <= 8'h10 ;
			data[30273] <= 8'h10 ;
			data[30274] <= 8'h10 ;
			data[30275] <= 8'h10 ;
			data[30276] <= 8'h10 ;
			data[30277] <= 8'h10 ;
			data[30278] <= 8'h10 ;
			data[30279] <= 8'h10 ;
			data[30280] <= 8'h10 ;
			data[30281] <= 8'h10 ;
			data[30282] <= 8'h10 ;
			data[30283] <= 8'h10 ;
			data[30284] <= 8'h10 ;
			data[30285] <= 8'h10 ;
			data[30286] <= 8'h10 ;
			data[30287] <= 8'h10 ;
			data[30288] <= 8'h10 ;
			data[30289] <= 8'h10 ;
			data[30290] <= 8'h10 ;
			data[30291] <= 8'h10 ;
			data[30292] <= 8'h10 ;
			data[30293] <= 8'h10 ;
			data[30294] <= 8'h10 ;
			data[30295] <= 8'h10 ;
			data[30296] <= 8'h10 ;
			data[30297] <= 8'h10 ;
			data[30298] <= 8'h10 ;
			data[30299] <= 8'h10 ;
			data[30300] <= 8'h10 ;
			data[30301] <= 8'h10 ;
			data[30302] <= 8'h10 ;
			data[30303] <= 8'h10 ;
			data[30304] <= 8'h10 ;
			data[30305] <= 8'h10 ;
			data[30306] <= 8'h10 ;
			data[30307] <= 8'h10 ;
			data[30308] <= 8'h10 ;
			data[30309] <= 8'h10 ;
			data[30310] <= 8'h10 ;
			data[30311] <= 8'h10 ;
			data[30312] <= 8'h10 ;
			data[30313] <= 8'h10 ;
			data[30314] <= 8'h10 ;
			data[30315] <= 8'h10 ;
			data[30316] <= 8'h10 ;
			data[30317] <= 8'h10 ;
			data[30318] <= 8'h10 ;
			data[30319] <= 8'h10 ;
			data[30320] <= 8'h10 ;
			data[30321] <= 8'h10 ;
			data[30322] <= 8'h10 ;
			data[30323] <= 8'h10 ;
			data[30324] <= 8'h10 ;
			data[30325] <= 8'h10 ;
			data[30326] <= 8'h10 ;
			data[30327] <= 8'h10 ;
			data[30328] <= 8'h10 ;
			data[30329] <= 8'h10 ;
			data[30330] <= 8'h10 ;
			data[30331] <= 8'h10 ;
			data[30332] <= 8'h10 ;
			data[30333] <= 8'h10 ;
			data[30334] <= 8'h10 ;
			data[30335] <= 8'h10 ;
			data[30336] <= 8'h10 ;
			data[30337] <= 8'h10 ;
			data[30338] <= 8'h10 ;
			data[30339] <= 8'h10 ;
			data[30340] <= 8'h10 ;
			data[30341] <= 8'h10 ;
			data[30342] <= 8'h10 ;
			data[30343] <= 8'h10 ;
			data[30344] <= 8'h10 ;
			data[30345] <= 8'h10 ;
			data[30346] <= 8'h10 ;
			data[30347] <= 8'h10 ;
			data[30348] <= 8'h10 ;
			data[30349] <= 8'h10 ;
			data[30350] <= 8'h10 ;
			data[30351] <= 8'h10 ;
			data[30352] <= 8'h10 ;
			data[30353] <= 8'h10 ;
			data[30354] <= 8'h10 ;
			data[30355] <= 8'h10 ;
			data[30356] <= 8'h10 ;
			data[30357] <= 8'h10 ;
			data[30358] <= 8'h10 ;
			data[30359] <= 8'h10 ;
			data[30360] <= 8'h10 ;
			data[30361] <= 8'h10 ;
			data[30362] <= 8'h10 ;
			data[30363] <= 8'h10 ;
			data[30364] <= 8'h10 ;
			data[30365] <= 8'h10 ;
			data[30366] <= 8'h10 ;
			data[30367] <= 8'h10 ;
			data[30368] <= 8'h10 ;
			data[30369] <= 8'h10 ;
			data[30370] <= 8'h10 ;
			data[30371] <= 8'h10 ;
			data[30372] <= 8'h10 ;
			data[30373] <= 8'h10 ;
			data[30374] <= 8'h10 ;
			data[30375] <= 8'h10 ;
			data[30376] <= 8'h10 ;
			data[30377] <= 8'h10 ;
			data[30378] <= 8'h10 ;
			data[30379] <= 8'h10 ;
			data[30380] <= 8'h10 ;
			data[30381] <= 8'h10 ;
			data[30382] <= 8'h10 ;
			data[30383] <= 8'h10 ;
			data[30384] <= 8'h10 ;
			data[30385] <= 8'h10 ;
			data[30386] <= 8'h10 ;
			data[30387] <= 8'h10 ;
			data[30388] <= 8'h10 ;
			data[30389] <= 8'h10 ;
			data[30390] <= 8'h10 ;
			data[30391] <= 8'h10 ;
			data[30392] <= 8'h10 ;
			data[30393] <= 8'h10 ;
			data[30394] <= 8'h10 ;
			data[30395] <= 8'h10 ;
			data[30396] <= 8'h10 ;
			data[30397] <= 8'h10 ;
			data[30398] <= 8'h10 ;
			data[30399] <= 8'h10 ;
			data[30400] <= 8'h10 ;
			data[30401] <= 8'h10 ;
			data[30402] <= 8'h10 ;
			data[30403] <= 8'h10 ;
			data[30404] <= 8'h10 ;
			data[30405] <= 8'h10 ;
			data[30406] <= 8'h10 ;
			data[30407] <= 8'h10 ;
			data[30408] <= 8'h10 ;
			data[30409] <= 8'h10 ;
			data[30410] <= 8'h10 ;
			data[30411] <= 8'h10 ;
			data[30412] <= 8'h10 ;
			data[30413] <= 8'h10 ;
			data[30414] <= 8'h10 ;
			data[30415] <= 8'h10 ;
			data[30416] <= 8'h10 ;
			data[30417] <= 8'h10 ;
			data[30418] <= 8'h10 ;
			data[30419] <= 8'h10 ;
			data[30420] <= 8'h10 ;
			data[30421] <= 8'h10 ;
			data[30422] <= 8'h10 ;
			data[30423] <= 8'h10 ;
			data[30424] <= 8'h10 ;
			data[30425] <= 8'h10 ;
			data[30426] <= 8'h10 ;
			data[30427] <= 8'h10 ;
			data[30428] <= 8'h10 ;
			data[30429] <= 8'h10 ;
			data[30430] <= 8'h10 ;
			data[30431] <= 8'h10 ;
			data[30432] <= 8'h10 ;
			data[30433] <= 8'h10 ;
			data[30434] <= 8'h10 ;
			data[30435] <= 8'h10 ;
			data[30436] <= 8'h10 ;
			data[30437] <= 8'h10 ;
			data[30438] <= 8'h10 ;
			data[30439] <= 8'h10 ;
			data[30440] <= 8'h10 ;
			data[30441] <= 8'h10 ;
			data[30442] <= 8'h10 ;
			data[30443] <= 8'h10 ;
			data[30444] <= 8'h10 ;
			data[30445] <= 8'h10 ;
			data[30446] <= 8'h10 ;
			data[30447] <= 8'h10 ;
			data[30448] <= 8'h10 ;
			data[30449] <= 8'h10 ;
			data[30450] <= 8'h10 ;
			data[30451] <= 8'h10 ;
			data[30452] <= 8'h10 ;
			data[30453] <= 8'h10 ;
			data[30454] <= 8'h10 ;
			data[30455] <= 8'h10 ;
			data[30456] <= 8'h10 ;
			data[30457] <= 8'h10 ;
			data[30458] <= 8'h10 ;
			data[30459] <= 8'h10 ;
			data[30460] <= 8'h10 ;
			data[30461] <= 8'h10 ;
			data[30462] <= 8'h10 ;
			data[30463] <= 8'h10 ;
			data[30464] <= 8'h10 ;
			data[30465] <= 8'h10 ;
			data[30466] <= 8'h10 ;
			data[30467] <= 8'h10 ;
			data[30468] <= 8'h10 ;
			data[30469] <= 8'h10 ;
			data[30470] <= 8'h10 ;
			data[30471] <= 8'h10 ;
			data[30472] <= 8'h10 ;
			data[30473] <= 8'h10 ;
			data[30474] <= 8'h10 ;
			data[30475] <= 8'h10 ;
			data[30476] <= 8'h10 ;
			data[30477] <= 8'h10 ;
			data[30478] <= 8'h10 ;
			data[30479] <= 8'h10 ;
			data[30480] <= 8'h10 ;
			data[30481] <= 8'h10 ;
			data[30482] <= 8'h10 ;
			data[30483] <= 8'h10 ;
			data[30484] <= 8'h10 ;
			data[30485] <= 8'h10 ;
			data[30486] <= 8'h10 ;
			data[30487] <= 8'h10 ;
			data[30488] <= 8'h10 ;
			data[30489] <= 8'h10 ;
			data[30490] <= 8'h10 ;
			data[30491] <= 8'h10 ;
			data[30492] <= 8'h10 ;
			data[30493] <= 8'h10 ;
			data[30494] <= 8'h10 ;
			data[30495] <= 8'h10 ;
			data[30496] <= 8'h10 ;
			data[30497] <= 8'h10 ;
			data[30498] <= 8'h10 ;
			data[30499] <= 8'h10 ;
			data[30500] <= 8'h10 ;
			data[30501] <= 8'h10 ;
			data[30502] <= 8'h10 ;
			data[30503] <= 8'h10 ;
			data[30504] <= 8'h10 ;
			data[30505] <= 8'h10 ;
			data[30506] <= 8'h10 ;
			data[30507] <= 8'h10 ;
			data[30508] <= 8'h10 ;
			data[30509] <= 8'h10 ;
			data[30510] <= 8'h10 ;
			data[30511] <= 8'h10 ;
			data[30512] <= 8'h10 ;
			data[30513] <= 8'h10 ;
			data[30514] <= 8'h10 ;
			data[30515] <= 8'h10 ;
			data[30516] <= 8'h10 ;
			data[30517] <= 8'h10 ;
			data[30518] <= 8'h10 ;
			data[30519] <= 8'h10 ;
			data[30520] <= 8'h10 ;
			data[30521] <= 8'h10 ;
			data[30522] <= 8'h10 ;
			data[30523] <= 8'h10 ;
			data[30524] <= 8'h10 ;
			data[30525] <= 8'h10 ;
			data[30526] <= 8'h10 ;
			data[30527] <= 8'h10 ;
			data[30528] <= 8'h10 ;
			data[30529] <= 8'h10 ;
			data[30530] <= 8'h10 ;
			data[30531] <= 8'h10 ;
			data[30532] <= 8'h10 ;
			data[30533] <= 8'h10 ;
			data[30534] <= 8'h10 ;
			data[30535] <= 8'h10 ;
			data[30536] <= 8'h10 ;
			data[30537] <= 8'h10 ;
			data[30538] <= 8'h10 ;
			data[30539] <= 8'h10 ;
			data[30540] <= 8'h10 ;
			data[30541] <= 8'h10 ;
			data[30542] <= 8'h10 ;
			data[30543] <= 8'h10 ;
			data[30544] <= 8'h10 ;
			data[30545] <= 8'h10 ;
			data[30546] <= 8'h10 ;
			data[30547] <= 8'h10 ;
			data[30548] <= 8'h10 ;
			data[30549] <= 8'h10 ;
			data[30550] <= 8'h10 ;
			data[30551] <= 8'h10 ;
			data[30552] <= 8'h10 ;
			data[30553] <= 8'h10 ;
			data[30554] <= 8'h10 ;
			data[30555] <= 8'h10 ;
			data[30556] <= 8'h10 ;
			data[30557] <= 8'h10 ;
			data[30558] <= 8'h10 ;
			data[30559] <= 8'h10 ;
			data[30560] <= 8'h10 ;
			data[30561] <= 8'h10 ;
			data[30562] <= 8'h10 ;
			data[30563] <= 8'h10 ;
			data[30564] <= 8'h10 ;
			data[30565] <= 8'h10 ;
			data[30566] <= 8'h10 ;
			data[30567] <= 8'h10 ;
			data[30568] <= 8'h10 ;
			data[30569] <= 8'h10 ;
			data[30570] <= 8'h10 ;
			data[30571] <= 8'h10 ;
			data[30572] <= 8'h10 ;
			data[30573] <= 8'h10 ;
			data[30574] <= 8'h10 ;
			data[30575] <= 8'h10 ;
			data[30576] <= 8'h10 ;
			data[30577] <= 8'h10 ;
			data[30578] <= 8'h10 ;
			data[30579] <= 8'h10 ;
			data[30580] <= 8'h10 ;
			data[30581] <= 8'h10 ;
			data[30582] <= 8'h10 ;
			data[30583] <= 8'h10 ;
			data[30584] <= 8'h10 ;
			data[30585] <= 8'h10 ;
			data[30586] <= 8'h10 ;
			data[30587] <= 8'h10 ;
			data[30588] <= 8'h10 ;
			data[30589] <= 8'h10 ;
			data[30590] <= 8'h10 ;
			data[30591] <= 8'h10 ;
			data[30592] <= 8'h10 ;
			data[30593] <= 8'h10 ;
			data[30594] <= 8'h10 ;
			data[30595] <= 8'h10 ;
			data[30596] <= 8'h10 ;
			data[30597] <= 8'h10 ;
			data[30598] <= 8'h10 ;
			data[30599] <= 8'h10 ;
			data[30600] <= 8'h10 ;
			data[30601] <= 8'h10 ;
			data[30602] <= 8'h10 ;
			data[30603] <= 8'h10 ;
			data[30604] <= 8'h10 ;
			data[30605] <= 8'h10 ;
			data[30606] <= 8'h10 ;
			data[30607] <= 8'h10 ;
			data[30608] <= 8'h10 ;
			data[30609] <= 8'h10 ;
			data[30610] <= 8'h10 ;
			data[30611] <= 8'h10 ;
			data[30612] <= 8'h10 ;
			data[30613] <= 8'h10 ;
			data[30614] <= 8'h10 ;
			data[30615] <= 8'h10 ;
			data[30616] <= 8'h10 ;
			data[30617] <= 8'h10 ;
			data[30618] <= 8'h10 ;
			data[30619] <= 8'h10 ;
			data[30620] <= 8'h10 ;
			data[30621] <= 8'h10 ;
			data[30622] <= 8'h10 ;
			data[30623] <= 8'h10 ;
			data[30624] <= 8'h10 ;
			data[30625] <= 8'h10 ;
			data[30626] <= 8'h10 ;
			data[30627] <= 8'h10 ;
			data[30628] <= 8'h10 ;
			data[30629] <= 8'h10 ;
			data[30630] <= 8'h10 ;
			data[30631] <= 8'h10 ;
			data[30632] <= 8'h10 ;
			data[30633] <= 8'h10 ;
			data[30634] <= 8'h10 ;
			data[30635] <= 8'h10 ;
			data[30636] <= 8'h10 ;
			data[30637] <= 8'h10 ;
			data[30638] <= 8'h10 ;
			data[30639] <= 8'h10 ;
			data[30640] <= 8'h10 ;
			data[30641] <= 8'h10 ;
			data[30642] <= 8'h10 ;
			data[30643] <= 8'h10 ;
			data[30644] <= 8'h10 ;
			data[30645] <= 8'h10 ;
			data[30646] <= 8'h10 ;
			data[30647] <= 8'h10 ;
			data[30648] <= 8'h10 ;
			data[30649] <= 8'h10 ;
			data[30650] <= 8'h10 ;
			data[30651] <= 8'h10 ;
			data[30652] <= 8'h10 ;
			data[30653] <= 8'h10 ;
			data[30654] <= 8'h10 ;
			data[30655] <= 8'h10 ;
			data[30656] <= 8'h10 ;
			data[30657] <= 8'h10 ;
			data[30658] <= 8'h10 ;
			data[30659] <= 8'h10 ;
			data[30660] <= 8'h10 ;
			data[30661] <= 8'h10 ;
			data[30662] <= 8'h10 ;
			data[30663] <= 8'h10 ;
			data[30664] <= 8'h10 ;
			data[30665] <= 8'h10 ;
			data[30666] <= 8'h10 ;
			data[30667] <= 8'h10 ;
			data[30668] <= 8'h10 ;
			data[30669] <= 8'h10 ;
			data[30670] <= 8'h10 ;
			data[30671] <= 8'h10 ;
			data[30672] <= 8'h10 ;
			data[30673] <= 8'h10 ;
			data[30674] <= 8'h10 ;
			data[30675] <= 8'h10 ;
			data[30676] <= 8'h10 ;
			data[30677] <= 8'h10 ;
			data[30678] <= 8'h10 ;
			data[30679] <= 8'h10 ;
			data[30680] <= 8'h10 ;
			data[30681] <= 8'h10 ;
			data[30682] <= 8'h10 ;
			data[30683] <= 8'h10 ;
			data[30684] <= 8'h10 ;
			data[30685] <= 8'h10 ;
			data[30686] <= 8'h10 ;
			data[30687] <= 8'h10 ;
			data[30688] <= 8'h10 ;
			data[30689] <= 8'h10 ;
			data[30690] <= 8'h10 ;
			data[30691] <= 8'h10 ;
			data[30692] <= 8'h10 ;
			data[30693] <= 8'h10 ;
			data[30694] <= 8'h10 ;
			data[30695] <= 8'h10 ;
			data[30696] <= 8'h10 ;
			data[30697] <= 8'h10 ;
			data[30698] <= 8'h10 ;
			data[30699] <= 8'h10 ;
			data[30700] <= 8'h10 ;
			data[30701] <= 8'h10 ;
			data[30702] <= 8'h10 ;
			data[30703] <= 8'h10 ;
			data[30704] <= 8'h10 ;
			data[30705] <= 8'h10 ;
			data[30706] <= 8'h10 ;
			data[30707] <= 8'h10 ;
			data[30708] <= 8'h10 ;
			data[30709] <= 8'h10 ;
			data[30710] <= 8'h10 ;
			data[30711] <= 8'h10 ;
			data[30712] <= 8'h10 ;
			data[30713] <= 8'h10 ;
			data[30714] <= 8'h10 ;
			data[30715] <= 8'h10 ;
			data[30716] <= 8'h10 ;
			data[30717] <= 8'h10 ;
			data[30718] <= 8'h10 ;
			data[30719] <= 8'h10 ;
			data[30720] <= 8'h10 ;
			data[30721] <= 8'h10 ;
			data[30722] <= 8'h10 ;
			data[30723] <= 8'h10 ;
			data[30724] <= 8'h10 ;
			data[30725] <= 8'h10 ;
			data[30726] <= 8'h10 ;
			data[30727] <= 8'h10 ;
			data[30728] <= 8'h10 ;
			data[30729] <= 8'h10 ;
			data[30730] <= 8'h10 ;
			data[30731] <= 8'h10 ;
			data[30732] <= 8'h10 ;
			data[30733] <= 8'h10 ;
			data[30734] <= 8'h10 ;
			data[30735] <= 8'h10 ;
			data[30736] <= 8'h10 ;
			data[30737] <= 8'h10 ;
			data[30738] <= 8'h10 ;
			data[30739] <= 8'h10 ;
			data[30740] <= 8'h10 ;
			data[30741] <= 8'h10 ;
			data[30742] <= 8'h10 ;
			data[30743] <= 8'h10 ;
			data[30744] <= 8'h10 ;
			data[30745] <= 8'h10 ;
			data[30746] <= 8'h10 ;
			data[30747] <= 8'h10 ;
			data[30748] <= 8'h10 ;
			data[30749] <= 8'h10 ;
			data[30750] <= 8'h10 ;
			data[30751] <= 8'h10 ;
			data[30752] <= 8'h10 ;
			data[30753] <= 8'h10 ;
			data[30754] <= 8'h10 ;
			data[30755] <= 8'h10 ;
			data[30756] <= 8'h10 ;
			data[30757] <= 8'h10 ;
			data[30758] <= 8'h10 ;
			data[30759] <= 8'h10 ;
			data[30760] <= 8'h10 ;
			data[30761] <= 8'h10 ;
			data[30762] <= 8'h10 ;
			data[30763] <= 8'h10 ;
			data[30764] <= 8'h10 ;
			data[30765] <= 8'h10 ;
			data[30766] <= 8'h10 ;
			data[30767] <= 8'h10 ;
			data[30768] <= 8'h10 ;
			data[30769] <= 8'h10 ;
			data[30770] <= 8'h10 ;
			data[30771] <= 8'h10 ;
			data[30772] <= 8'h10 ;
			data[30773] <= 8'h10 ;
			data[30774] <= 8'h10 ;
			data[30775] <= 8'h10 ;
			data[30776] <= 8'h10 ;
			data[30777] <= 8'h10 ;
			data[30778] <= 8'h10 ;
			data[30779] <= 8'h10 ;
			data[30780] <= 8'h10 ;
			data[30781] <= 8'h10 ;
			data[30782] <= 8'h10 ;
			data[30783] <= 8'h10 ;
			data[30784] <= 8'h10 ;
			data[30785] <= 8'h10 ;
			data[30786] <= 8'h10 ;
			data[30787] <= 8'h10 ;
			data[30788] <= 8'h10 ;
			data[30789] <= 8'h10 ;
			data[30790] <= 8'h10 ;
			data[30791] <= 8'h10 ;
			data[30792] <= 8'h10 ;
			data[30793] <= 8'h10 ;
			data[30794] <= 8'h10 ;
			data[30795] <= 8'h10 ;
			data[30796] <= 8'h10 ;
			data[30797] <= 8'h10 ;
			data[30798] <= 8'h10 ;
			data[30799] <= 8'h10 ;
			data[30800] <= 8'h10 ;
			data[30801] <= 8'h10 ;
			data[30802] <= 8'h10 ;
			data[30803] <= 8'h10 ;
			data[30804] <= 8'h10 ;
			data[30805] <= 8'h10 ;
			data[30806] <= 8'h10 ;
			data[30807] <= 8'h10 ;
			data[30808] <= 8'h10 ;
			data[30809] <= 8'h10 ;
			data[30810] <= 8'h10 ;
			data[30811] <= 8'h10 ;
			data[30812] <= 8'h10 ;
			data[30813] <= 8'h10 ;
			data[30814] <= 8'h10 ;
			data[30815] <= 8'h10 ;
			data[30816] <= 8'h10 ;
			data[30817] <= 8'h10 ;
			data[30818] <= 8'h10 ;
			data[30819] <= 8'h10 ;
			data[30820] <= 8'h10 ;
			data[30821] <= 8'h10 ;
			data[30822] <= 8'h10 ;
			data[30823] <= 8'h10 ;
			data[30824] <= 8'h10 ;
			data[30825] <= 8'h10 ;
			data[30826] <= 8'h10 ;
			data[30827] <= 8'h10 ;
			data[30828] <= 8'h10 ;
			data[30829] <= 8'h10 ;
			data[30830] <= 8'h10 ;
			data[30831] <= 8'h10 ;
			data[30832] <= 8'h10 ;
			data[30833] <= 8'h10 ;
			data[30834] <= 8'h10 ;
			data[30835] <= 8'h10 ;
			data[30836] <= 8'h10 ;
			data[30837] <= 8'h10 ;
			data[30838] <= 8'h10 ;
			data[30839] <= 8'h10 ;
			data[30840] <= 8'h10 ;
			data[30841] <= 8'h10 ;
			data[30842] <= 8'h10 ;
			data[30843] <= 8'h10 ;
			data[30844] <= 8'h10 ;
			data[30845] <= 8'h10 ;
			data[30846] <= 8'h10 ;
			data[30847] <= 8'h10 ;
			data[30848] <= 8'h10 ;
			data[30849] <= 8'h10 ;
			data[30850] <= 8'h10 ;
			data[30851] <= 8'h10 ;
			data[30852] <= 8'h10 ;
			data[30853] <= 8'h10 ;
			data[30854] <= 8'h10 ;
			data[30855] <= 8'h10 ;
			data[30856] <= 8'h10 ;
			data[30857] <= 8'h10 ;
			data[30858] <= 8'h10 ;
			data[30859] <= 8'h10 ;
			data[30860] <= 8'h10 ;
			data[30861] <= 8'h10 ;
			data[30862] <= 8'h10 ;
			data[30863] <= 8'h10 ;
			data[30864] <= 8'h10 ;
			data[30865] <= 8'h10 ;
			data[30866] <= 8'h10 ;
			data[30867] <= 8'h10 ;
			data[30868] <= 8'h10 ;
			data[30869] <= 8'h10 ;
			data[30870] <= 8'h10 ;
			data[30871] <= 8'h10 ;
			data[30872] <= 8'h10 ;
			data[30873] <= 8'h10 ;
			data[30874] <= 8'h10 ;
			data[30875] <= 8'h10 ;
			data[30876] <= 8'h10 ;
			data[30877] <= 8'h10 ;
			data[30878] <= 8'h10 ;
			data[30879] <= 8'h10 ;
			data[30880] <= 8'h10 ;
			data[30881] <= 8'h10 ;
			data[30882] <= 8'h10 ;
			data[30883] <= 8'h10 ;
			data[30884] <= 8'h10 ;
			data[30885] <= 8'h10 ;
			data[30886] <= 8'h10 ;
			data[30887] <= 8'h10 ;
			data[30888] <= 8'h10 ;
			data[30889] <= 8'h10 ;
			data[30890] <= 8'h10 ;
			data[30891] <= 8'h10 ;
			data[30892] <= 8'h10 ;
			data[30893] <= 8'h10 ;
			data[30894] <= 8'h10 ;
			data[30895] <= 8'h10 ;
			data[30896] <= 8'h10 ;
			data[30897] <= 8'h10 ;
			data[30898] <= 8'h10 ;
			data[30899] <= 8'h10 ;
			data[30900] <= 8'h10 ;
			data[30901] <= 8'h10 ;
			data[30902] <= 8'h10 ;
			data[30903] <= 8'h10 ;
			data[30904] <= 8'h10 ;
			data[30905] <= 8'h10 ;
			data[30906] <= 8'h10 ;
			data[30907] <= 8'h10 ;
			data[30908] <= 8'h10 ;
			data[30909] <= 8'h10 ;
			data[30910] <= 8'h10 ;
			data[30911] <= 8'h10 ;
			data[30912] <= 8'h10 ;
			data[30913] <= 8'h10 ;
			data[30914] <= 8'h10 ;
			data[30915] <= 8'h10 ;
			data[30916] <= 8'h10 ;
			data[30917] <= 8'h10 ;
			data[30918] <= 8'h10 ;
			data[30919] <= 8'h10 ;
			data[30920] <= 8'h10 ;
			data[30921] <= 8'h10 ;
			data[30922] <= 8'h10 ;
			data[30923] <= 8'h10 ;
			data[30924] <= 8'h10 ;
			data[30925] <= 8'h10 ;
			data[30926] <= 8'h10 ;
			data[30927] <= 8'h10 ;
			data[30928] <= 8'h10 ;
			data[30929] <= 8'h10 ;
			data[30930] <= 8'h10 ;
			data[30931] <= 8'h10 ;
			data[30932] <= 8'h10 ;
			data[30933] <= 8'h10 ;
			data[30934] <= 8'h10 ;
			data[30935] <= 8'h10 ;
			data[30936] <= 8'h10 ;
			data[30937] <= 8'h10 ;
			data[30938] <= 8'h10 ;
			data[30939] <= 8'h10 ;
			data[30940] <= 8'h10 ;
			data[30941] <= 8'h10 ;
			data[30942] <= 8'h10 ;
			data[30943] <= 8'h10 ;
			data[30944] <= 8'h10 ;
			data[30945] <= 8'h10 ;
			data[30946] <= 8'h10 ;
			data[30947] <= 8'h10 ;
			data[30948] <= 8'h10 ;
			data[30949] <= 8'h10 ;
			data[30950] <= 8'h10 ;
			data[30951] <= 8'h10 ;
			data[30952] <= 8'h10 ;
			data[30953] <= 8'h10 ;
			data[30954] <= 8'h10 ;
			data[30955] <= 8'h10 ;
			data[30956] <= 8'h10 ;
			data[30957] <= 8'h10 ;
			data[30958] <= 8'h10 ;
			data[30959] <= 8'h10 ;
			data[30960] <= 8'h10 ;
			data[30961] <= 8'h10 ;
			data[30962] <= 8'h10 ;
			data[30963] <= 8'h10 ;
			data[30964] <= 8'h10 ;
			data[30965] <= 8'h10 ;
			data[30966] <= 8'h10 ;
			data[30967] <= 8'h10 ;
			data[30968] <= 8'h10 ;
			data[30969] <= 8'h10 ;
			data[30970] <= 8'h10 ;
			data[30971] <= 8'h10 ;
			data[30972] <= 8'h10 ;
			data[30973] <= 8'h10 ;
			data[30974] <= 8'h10 ;
			data[30975] <= 8'h10 ;
			data[30976] <= 8'h10 ;
			data[30977] <= 8'h10 ;
			data[30978] <= 8'h10 ;
			data[30979] <= 8'h10 ;
			data[30980] <= 8'h10 ;
			data[30981] <= 8'h10 ;
			data[30982] <= 8'h10 ;
			data[30983] <= 8'h10 ;
			data[30984] <= 8'h10 ;
			data[30985] <= 8'h10 ;
			data[30986] <= 8'h10 ;
			data[30987] <= 8'h10 ;
			data[30988] <= 8'h10 ;
			data[30989] <= 8'h10 ;
			data[30990] <= 8'h10 ;
			data[30991] <= 8'h10 ;
			data[30992] <= 8'h10 ;
			data[30993] <= 8'h10 ;
			data[30994] <= 8'h10 ;
			data[30995] <= 8'h10 ;
			data[30996] <= 8'h10 ;
			data[30997] <= 8'h10 ;
			data[30998] <= 8'h10 ;
			data[30999] <= 8'h10 ;
			data[31000] <= 8'h10 ;
			data[31001] <= 8'h10 ;
			data[31002] <= 8'h10 ;
			data[31003] <= 8'h10 ;
			data[31004] <= 8'h10 ;
			data[31005] <= 8'h10 ;
			data[31006] <= 8'h10 ;
			data[31007] <= 8'h10 ;
			data[31008] <= 8'h10 ;
			data[31009] <= 8'h10 ;
			data[31010] <= 8'h10 ;
			data[31011] <= 8'h10 ;
			data[31012] <= 8'h10 ;
			data[31013] <= 8'h10 ;
			data[31014] <= 8'h10 ;
			data[31015] <= 8'h10 ;
			data[31016] <= 8'h10 ;
			data[31017] <= 8'h10 ;
			data[31018] <= 8'h10 ;
			data[31019] <= 8'h10 ;
			data[31020] <= 8'h10 ;
			data[31021] <= 8'h10 ;
			data[31022] <= 8'h10 ;
			data[31023] <= 8'h10 ;
			data[31024] <= 8'h10 ;
			data[31025] <= 8'h10 ;
			data[31026] <= 8'h10 ;
			data[31027] <= 8'h10 ;
			data[31028] <= 8'h10 ;
			data[31029] <= 8'h10 ;
			data[31030] <= 8'h10 ;
			data[31031] <= 8'h10 ;
			data[31032] <= 8'h10 ;
			data[31033] <= 8'h10 ;
			data[31034] <= 8'h10 ;
			data[31035] <= 8'h10 ;
			data[31036] <= 8'h10 ;
			data[31037] <= 8'h10 ;
			data[31038] <= 8'h10 ;
			data[31039] <= 8'h10 ;
			data[31040] <= 8'h10 ;
			data[31041] <= 8'h10 ;
			data[31042] <= 8'h10 ;
			data[31043] <= 8'h10 ;
			data[31044] <= 8'h10 ;
			data[31045] <= 8'h10 ;
			data[31046] <= 8'h10 ;
			data[31047] <= 8'h10 ;
			data[31048] <= 8'h10 ;
			data[31049] <= 8'h10 ;
			data[31050] <= 8'h10 ;
			data[31051] <= 8'h10 ;
			data[31052] <= 8'h10 ;
			data[31053] <= 8'h10 ;
			data[31054] <= 8'h10 ;
			data[31055] <= 8'h10 ;
			data[31056] <= 8'h10 ;
			data[31057] <= 8'h10 ;
			data[31058] <= 8'h10 ;
			data[31059] <= 8'h10 ;
			data[31060] <= 8'h10 ;
			data[31061] <= 8'h10 ;
			data[31062] <= 8'h10 ;
			data[31063] <= 8'h10 ;
			data[31064] <= 8'h10 ;
			data[31065] <= 8'h10 ;
			data[31066] <= 8'h10 ;
			data[31067] <= 8'h10 ;
			data[31068] <= 8'h10 ;
			data[31069] <= 8'h10 ;
			data[31070] <= 8'h10 ;
			data[31071] <= 8'h10 ;
			data[31072] <= 8'h10 ;
			data[31073] <= 8'h10 ;
			data[31074] <= 8'h10 ;
			data[31075] <= 8'h10 ;
			data[31076] <= 8'h10 ;
			data[31077] <= 8'h10 ;
			data[31078] <= 8'h10 ;
			data[31079] <= 8'h10 ;
			data[31080] <= 8'h10 ;
			data[31081] <= 8'h10 ;
			data[31082] <= 8'h10 ;
			data[31083] <= 8'h10 ;
			data[31084] <= 8'h10 ;
			data[31085] <= 8'h10 ;
			data[31086] <= 8'h10 ;
			data[31087] <= 8'h10 ;
			data[31088] <= 8'h10 ;
			data[31089] <= 8'h10 ;
			data[31090] <= 8'h10 ;
			data[31091] <= 8'h10 ;
			data[31092] <= 8'h10 ;
			data[31093] <= 8'h10 ;
			data[31094] <= 8'h10 ;
			data[31095] <= 8'h10 ;
			data[31096] <= 8'h10 ;
			data[31097] <= 8'h10 ;
			data[31098] <= 8'h10 ;
			data[31099] <= 8'h10 ;
			data[31100] <= 8'h10 ;
			data[31101] <= 8'h10 ;
			data[31102] <= 8'h10 ;
			data[31103] <= 8'h10 ;
			data[31104] <= 8'h10 ;
			data[31105] <= 8'h10 ;
			data[31106] <= 8'h10 ;
			data[31107] <= 8'h10 ;
			data[31108] <= 8'h10 ;
			data[31109] <= 8'h10 ;
			data[31110] <= 8'h10 ;
			data[31111] <= 8'h10 ;
			data[31112] <= 8'h10 ;
			data[31113] <= 8'h10 ;
			data[31114] <= 8'h10 ;
			data[31115] <= 8'h10 ;
			data[31116] <= 8'h10 ;
			data[31117] <= 8'h10 ;
			data[31118] <= 8'h10 ;
			data[31119] <= 8'h10 ;
			data[31120] <= 8'h10 ;
			data[31121] <= 8'h10 ;
			data[31122] <= 8'h10 ;
			data[31123] <= 8'h10 ;
			data[31124] <= 8'h10 ;
			data[31125] <= 8'h10 ;
			data[31126] <= 8'h10 ;
			data[31127] <= 8'h10 ;
			data[31128] <= 8'h10 ;
			data[31129] <= 8'h10 ;
			data[31130] <= 8'h10 ;
			data[31131] <= 8'h10 ;
			data[31132] <= 8'h10 ;
			data[31133] <= 8'h10 ;
			data[31134] <= 8'h10 ;
			data[31135] <= 8'h10 ;
			data[31136] <= 8'h10 ;
			data[31137] <= 8'h10 ;
			data[31138] <= 8'h10 ;
			data[31139] <= 8'h10 ;
			data[31140] <= 8'h10 ;
			data[31141] <= 8'h10 ;
			data[31142] <= 8'h10 ;
			data[31143] <= 8'h10 ;
			data[31144] <= 8'h10 ;
			data[31145] <= 8'h10 ;
			data[31146] <= 8'h10 ;
			data[31147] <= 8'h10 ;
			data[31148] <= 8'h10 ;
			data[31149] <= 8'h10 ;
			data[31150] <= 8'h10 ;
			data[31151] <= 8'h10 ;
			data[31152] <= 8'h10 ;
			data[31153] <= 8'h10 ;
			data[31154] <= 8'h10 ;
			data[31155] <= 8'h10 ;
			data[31156] <= 8'h10 ;
			data[31157] <= 8'h10 ;
			data[31158] <= 8'h10 ;
			data[31159] <= 8'h10 ;
			data[31160] <= 8'h10 ;
			data[31161] <= 8'h10 ;
			data[31162] <= 8'h10 ;
			data[31163] <= 8'h10 ;
			data[31164] <= 8'h10 ;
			data[31165] <= 8'h10 ;
			data[31166] <= 8'h10 ;
			data[31167] <= 8'h10 ;
			data[31168] <= 8'h10 ;
			data[31169] <= 8'h10 ;
			data[31170] <= 8'h10 ;
			data[31171] <= 8'h10 ;
			data[31172] <= 8'h10 ;
			data[31173] <= 8'h10 ;
			data[31174] <= 8'h10 ;
			data[31175] <= 8'h10 ;
			data[31176] <= 8'h10 ;
			data[31177] <= 8'h10 ;
			data[31178] <= 8'h10 ;
			data[31179] <= 8'h10 ;
			data[31180] <= 8'h10 ;
			data[31181] <= 8'h10 ;
			data[31182] <= 8'h10 ;
			data[31183] <= 8'h10 ;
			data[31184] <= 8'h10 ;
			data[31185] <= 8'h10 ;
			data[31186] <= 8'h10 ;
			data[31187] <= 8'h10 ;
			data[31188] <= 8'h10 ;
			data[31189] <= 8'h10 ;
			data[31190] <= 8'h10 ;
			data[31191] <= 8'h10 ;
			data[31192] <= 8'h10 ;
			data[31193] <= 8'h10 ;
			data[31194] <= 8'h10 ;
			data[31195] <= 8'h10 ;
			data[31196] <= 8'h10 ;
			data[31197] <= 8'h10 ;
			data[31198] <= 8'h10 ;
			data[31199] <= 8'h10 ;
			data[31200] <= 8'h10 ;
			data[31201] <= 8'h10 ;
			data[31202] <= 8'h10 ;
			data[31203] <= 8'h10 ;
			data[31204] <= 8'h10 ;
			data[31205] <= 8'h10 ;
			data[31206] <= 8'h10 ;
			data[31207] <= 8'h10 ;
			data[31208] <= 8'h10 ;
			data[31209] <= 8'h10 ;
			data[31210] <= 8'h10 ;
			data[31211] <= 8'h10 ;
			data[31212] <= 8'h10 ;
			data[31213] <= 8'h10 ;
			data[31214] <= 8'h10 ;
			data[31215] <= 8'h10 ;
			data[31216] <= 8'h10 ;
			data[31217] <= 8'h10 ;
			data[31218] <= 8'h10 ;
			data[31219] <= 8'h10 ;
			data[31220] <= 8'h10 ;
			data[31221] <= 8'h10 ;
			data[31222] <= 8'h10 ;
			data[31223] <= 8'h10 ;
			data[31224] <= 8'h10 ;
			data[31225] <= 8'h10 ;
			data[31226] <= 8'h10 ;
			data[31227] <= 8'h10 ;
			data[31228] <= 8'h10 ;
			data[31229] <= 8'h10 ;
			data[31230] <= 8'h10 ;
			data[31231] <= 8'h10 ;
			data[31232] <= 8'h10 ;
			data[31233] <= 8'h10 ;
			data[31234] <= 8'h10 ;
			data[31235] <= 8'h10 ;
			data[31236] <= 8'h10 ;
			data[31237] <= 8'h10 ;
			data[31238] <= 8'h10 ;
			data[31239] <= 8'h10 ;
			data[31240] <= 8'h10 ;
			data[31241] <= 8'h10 ;
			data[31242] <= 8'h10 ;
			data[31243] <= 8'h10 ;
			data[31244] <= 8'h10 ;
			data[31245] <= 8'h10 ;
			data[31246] <= 8'h10 ;
			data[31247] <= 8'h10 ;
			data[31248] <= 8'h10 ;
			data[31249] <= 8'h10 ;
			data[31250] <= 8'h10 ;
			data[31251] <= 8'h10 ;
			data[31252] <= 8'h10 ;
			data[31253] <= 8'h10 ;
			data[31254] <= 8'h10 ;
			data[31255] <= 8'h10 ;
			data[31256] <= 8'h10 ;
			data[31257] <= 8'h10 ;
			data[31258] <= 8'h10 ;
			data[31259] <= 8'h10 ;
			data[31260] <= 8'h10 ;
			data[31261] <= 8'h10 ;
			data[31262] <= 8'h10 ;
			data[31263] <= 8'h10 ;
			data[31264] <= 8'h10 ;
			data[31265] <= 8'h10 ;
			data[31266] <= 8'h10 ;
			data[31267] <= 8'h10 ;
			data[31268] <= 8'h10 ;
			data[31269] <= 8'h10 ;
			data[31270] <= 8'h10 ;
			data[31271] <= 8'h10 ;
			data[31272] <= 8'h10 ;
			data[31273] <= 8'h10 ;
			data[31274] <= 8'h10 ;
			data[31275] <= 8'h10 ;
			data[31276] <= 8'h10 ;
			data[31277] <= 8'h10 ;
			data[31278] <= 8'h10 ;
			data[31279] <= 8'h10 ;
			data[31280] <= 8'h10 ;
			data[31281] <= 8'h10 ;
			data[31282] <= 8'h10 ;
			data[31283] <= 8'h10 ;
			data[31284] <= 8'h10 ;
			data[31285] <= 8'h10 ;
			data[31286] <= 8'h10 ;
			data[31287] <= 8'h10 ;
			data[31288] <= 8'h10 ;
			data[31289] <= 8'h10 ;
			data[31290] <= 8'h10 ;
			data[31291] <= 8'h10 ;
			data[31292] <= 8'h10 ;
			data[31293] <= 8'h10 ;
			data[31294] <= 8'h10 ;
			data[31295] <= 8'h10 ;
			data[31296] <= 8'h10 ;
			data[31297] <= 8'h10 ;
			data[31298] <= 8'h10 ;
			data[31299] <= 8'h10 ;
			data[31300] <= 8'h10 ;
			data[31301] <= 8'h10 ;
			data[31302] <= 8'h10 ;
			data[31303] <= 8'h10 ;
			data[31304] <= 8'h10 ;
			data[31305] <= 8'h10 ;
			data[31306] <= 8'h10 ;
			data[31307] <= 8'h10 ;
			data[31308] <= 8'h10 ;
			data[31309] <= 8'h10 ;
			data[31310] <= 8'h10 ;
			data[31311] <= 8'h10 ;
			data[31312] <= 8'h10 ;
			data[31313] <= 8'h10 ;
			data[31314] <= 8'h10 ;
			data[31315] <= 8'h10 ;
			data[31316] <= 8'h10 ;
			data[31317] <= 8'h10 ;
			data[31318] <= 8'h10 ;
			data[31319] <= 8'h10 ;
			data[31320] <= 8'h10 ;
			data[31321] <= 8'h10 ;
			data[31322] <= 8'h10 ;
			data[31323] <= 8'h10 ;
			data[31324] <= 8'h10 ;
			data[31325] <= 8'h10 ;
			data[31326] <= 8'h10 ;
			data[31327] <= 8'h10 ;
			data[31328] <= 8'h10 ;
			data[31329] <= 8'h10 ;
			data[31330] <= 8'h10 ;
			data[31331] <= 8'h10 ;
			data[31332] <= 8'h10 ;
			data[31333] <= 8'h10 ;
			data[31334] <= 8'h10 ;
			data[31335] <= 8'h10 ;
			data[31336] <= 8'h10 ;
			data[31337] <= 8'h10 ;
			data[31338] <= 8'h10 ;
			data[31339] <= 8'h10 ;
			data[31340] <= 8'h10 ;
			data[31341] <= 8'h10 ;
			data[31342] <= 8'h10 ;
			data[31343] <= 8'h10 ;
			data[31344] <= 8'h10 ;
			data[31345] <= 8'h10 ;
			data[31346] <= 8'h10 ;
			data[31347] <= 8'h10 ;
			data[31348] <= 8'h10 ;
			data[31349] <= 8'h10 ;
			data[31350] <= 8'h10 ;
			data[31351] <= 8'h10 ;
			data[31352] <= 8'h10 ;
			data[31353] <= 8'h10 ;
			data[31354] <= 8'h10 ;
			data[31355] <= 8'h10 ;
			data[31356] <= 8'h10 ;
			data[31357] <= 8'h10 ;
			data[31358] <= 8'h10 ;
			data[31359] <= 8'h10 ;
			data[31360] <= 8'h10 ;
			data[31361] <= 8'h10 ;
			data[31362] <= 8'h10 ;
			data[31363] <= 8'h10 ;
			data[31364] <= 8'h10 ;
			data[31365] <= 8'h10 ;
			data[31366] <= 8'h10 ;
			data[31367] <= 8'h10 ;
			data[31368] <= 8'h10 ;
			data[31369] <= 8'h10 ;
			data[31370] <= 8'h10 ;
			data[31371] <= 8'h10 ;
			data[31372] <= 8'h10 ;
			data[31373] <= 8'h10 ;
			data[31374] <= 8'h10 ;
			data[31375] <= 8'h10 ;
			data[31376] <= 8'h10 ;
			data[31377] <= 8'h10 ;
			data[31378] <= 8'h10 ;
			data[31379] <= 8'h10 ;
			data[31380] <= 8'h10 ;
			data[31381] <= 8'h10 ;
			data[31382] <= 8'h10 ;
			data[31383] <= 8'h10 ;
			data[31384] <= 8'h10 ;
			data[31385] <= 8'h10 ;
			data[31386] <= 8'h10 ;
			data[31387] <= 8'h10 ;
			data[31388] <= 8'h10 ;
			data[31389] <= 8'h10 ;
			data[31390] <= 8'h10 ;
			data[31391] <= 8'h10 ;
			data[31392] <= 8'h10 ;
			data[31393] <= 8'h10 ;
			data[31394] <= 8'h10 ;
			data[31395] <= 8'h10 ;
			data[31396] <= 8'h10 ;
			data[31397] <= 8'h10 ;
			data[31398] <= 8'h10 ;
			data[31399] <= 8'h10 ;
			data[31400] <= 8'h10 ;
			data[31401] <= 8'h10 ;
			data[31402] <= 8'h10 ;
			data[31403] <= 8'h10 ;
			data[31404] <= 8'h10 ;
			data[31405] <= 8'h10 ;
			data[31406] <= 8'h10 ;
			data[31407] <= 8'h10 ;
			data[31408] <= 8'h10 ;
			data[31409] <= 8'h10 ;
			data[31410] <= 8'h10 ;
			data[31411] <= 8'h10 ;
			data[31412] <= 8'h10 ;
			data[31413] <= 8'h10 ;
			data[31414] <= 8'h10 ;
			data[31415] <= 8'h10 ;
			data[31416] <= 8'h10 ;
			data[31417] <= 8'h10 ;
			data[31418] <= 8'h10 ;
			data[31419] <= 8'h10 ;
			data[31420] <= 8'h10 ;
			data[31421] <= 8'h10 ;
			data[31422] <= 8'h10 ;
			data[31423] <= 8'h10 ;
			data[31424] <= 8'h10 ;
			data[31425] <= 8'h10 ;
			data[31426] <= 8'h10 ;
			data[31427] <= 8'h10 ;
			data[31428] <= 8'h10 ;
			data[31429] <= 8'h10 ;
			data[31430] <= 8'h10 ;
			data[31431] <= 8'h10 ;
			data[31432] <= 8'h10 ;
			data[31433] <= 8'h10 ;
			data[31434] <= 8'h10 ;
			data[31435] <= 8'h10 ;
			data[31436] <= 8'h10 ;
			data[31437] <= 8'h10 ;
			data[31438] <= 8'h10 ;
			data[31439] <= 8'h10 ;
			data[31440] <= 8'h10 ;
			data[31441] <= 8'h10 ;
			data[31442] <= 8'h10 ;
			data[31443] <= 8'h10 ;
			data[31444] <= 8'h10 ;
			data[31445] <= 8'h10 ;
			data[31446] <= 8'h10 ;
			data[31447] <= 8'h10 ;
			data[31448] <= 8'h10 ;
			data[31449] <= 8'h10 ;
			data[31450] <= 8'h10 ;
			data[31451] <= 8'h10 ;
			data[31452] <= 8'h10 ;
			data[31453] <= 8'h10 ;
			data[31454] <= 8'h10 ;
			data[31455] <= 8'h10 ;
			data[31456] <= 8'h10 ;
			data[31457] <= 8'h10 ;
			data[31458] <= 8'h10 ;
			data[31459] <= 8'h10 ;
			data[31460] <= 8'h10 ;
			data[31461] <= 8'h10 ;
			data[31462] <= 8'h10 ;
			data[31463] <= 8'h10 ;
			data[31464] <= 8'h10 ;
			data[31465] <= 8'h10 ;
			data[31466] <= 8'h10 ;
			data[31467] <= 8'h10 ;
			data[31468] <= 8'h10 ;
			data[31469] <= 8'h10 ;
			data[31470] <= 8'h10 ;
			data[31471] <= 8'h10 ;
			data[31472] <= 8'h10 ;
			data[31473] <= 8'h10 ;
			data[31474] <= 8'h10 ;
			data[31475] <= 8'h10 ;
			data[31476] <= 8'h10 ;
			data[31477] <= 8'h10 ;
			data[31478] <= 8'h10 ;
			data[31479] <= 8'h10 ;
			data[31480] <= 8'h10 ;
			data[31481] <= 8'h10 ;
			data[31482] <= 8'h10 ;
			data[31483] <= 8'h10 ;
			data[31484] <= 8'h10 ;
			data[31485] <= 8'h10 ;
			data[31486] <= 8'h10 ;
			data[31487] <= 8'h10 ;
			data[31488] <= 8'h10 ;
			data[31489] <= 8'h10 ;
			data[31490] <= 8'h10 ;
			data[31491] <= 8'h10 ;
			data[31492] <= 8'h10 ;
			data[31493] <= 8'h10 ;
			data[31494] <= 8'h10 ;
			data[31495] <= 8'h10 ;
			data[31496] <= 8'h10 ;
			data[31497] <= 8'h10 ;
			data[31498] <= 8'h10 ;
			data[31499] <= 8'h10 ;
			data[31500] <= 8'h10 ;
			data[31501] <= 8'h10 ;
			data[31502] <= 8'h10 ;
			data[31503] <= 8'h10 ;
			data[31504] <= 8'h10 ;
			data[31505] <= 8'h10 ;
			data[31506] <= 8'h10 ;
			data[31507] <= 8'h10 ;
			data[31508] <= 8'h10 ;
			data[31509] <= 8'h10 ;
			data[31510] <= 8'h10 ;
			data[31511] <= 8'h10 ;
			data[31512] <= 8'h10 ;
			data[31513] <= 8'h10 ;
			data[31514] <= 8'h10 ;
			data[31515] <= 8'h10 ;
			data[31516] <= 8'h10 ;
			data[31517] <= 8'h10 ;
			data[31518] <= 8'h10 ;
			data[31519] <= 8'h10 ;
			data[31520] <= 8'h10 ;
			data[31521] <= 8'h10 ;
			data[31522] <= 8'h10 ;
			data[31523] <= 8'h10 ;
			data[31524] <= 8'h10 ;
			data[31525] <= 8'h10 ;
			data[31526] <= 8'h10 ;
			data[31527] <= 8'h10 ;
			data[31528] <= 8'h10 ;
			data[31529] <= 8'h10 ;
			data[31530] <= 8'h10 ;
			data[31531] <= 8'h10 ;
			data[31532] <= 8'h10 ;
			data[31533] <= 8'h10 ;
			data[31534] <= 8'h10 ;
			data[31535] <= 8'h10 ;
			data[31536] <= 8'h10 ;
			data[31537] <= 8'h10 ;
			data[31538] <= 8'h10 ;
			data[31539] <= 8'h10 ;
			data[31540] <= 8'h10 ;
			data[31541] <= 8'h10 ;
			data[31542] <= 8'h10 ;
			data[31543] <= 8'h10 ;
			data[31544] <= 8'h10 ;
			data[31545] <= 8'h10 ;
			data[31546] <= 8'h10 ;
			data[31547] <= 8'h10 ;
			data[31548] <= 8'h10 ;
			data[31549] <= 8'h10 ;
			data[31550] <= 8'h10 ;
			data[31551] <= 8'h10 ;
			data[31552] <= 8'h10 ;
			data[31553] <= 8'h10 ;
			data[31554] <= 8'h10 ;
			data[31555] <= 8'h10 ;
			data[31556] <= 8'h10 ;
			data[31557] <= 8'h10 ;
			data[31558] <= 8'h10 ;
			data[31559] <= 8'h10 ;
			data[31560] <= 8'h10 ;
			data[31561] <= 8'h10 ;
			data[31562] <= 8'h10 ;
			data[31563] <= 8'h10 ;
			data[31564] <= 8'h10 ;
			data[31565] <= 8'h10 ;
			data[31566] <= 8'h10 ;
			data[31567] <= 8'h10 ;
			data[31568] <= 8'h10 ;
			data[31569] <= 8'h10 ;
			data[31570] <= 8'h10 ;
			data[31571] <= 8'h10 ;
			data[31572] <= 8'h10 ;
			data[31573] <= 8'h10 ;
			data[31574] <= 8'h10 ;
			data[31575] <= 8'h10 ;
			data[31576] <= 8'h10 ;
			data[31577] <= 8'h10 ;
			data[31578] <= 8'h10 ;
			data[31579] <= 8'h10 ;
			data[31580] <= 8'h10 ;
			data[31581] <= 8'h10 ;
			data[31582] <= 8'h10 ;
			data[31583] <= 8'h10 ;
			data[31584] <= 8'h10 ;
			data[31585] <= 8'h10 ;
			data[31586] <= 8'h10 ;
			data[31587] <= 8'h10 ;
			data[31588] <= 8'h10 ;
			data[31589] <= 8'h10 ;
			data[31590] <= 8'h10 ;
			data[31591] <= 8'h10 ;
			data[31592] <= 8'h10 ;
			data[31593] <= 8'h10 ;
			data[31594] <= 8'h10 ;
			data[31595] <= 8'h10 ;
			data[31596] <= 8'h10 ;
			data[31597] <= 8'h10 ;
			data[31598] <= 8'h10 ;
			data[31599] <= 8'h10 ;
			data[31600] <= 8'h10 ;
			data[31601] <= 8'h10 ;
			data[31602] <= 8'h10 ;
			data[31603] <= 8'h10 ;
			data[31604] <= 8'h10 ;
			data[31605] <= 8'h10 ;
			data[31606] <= 8'h10 ;
			data[31607] <= 8'h10 ;
			data[31608] <= 8'h10 ;
			data[31609] <= 8'h10 ;
			data[31610] <= 8'h10 ;
			data[31611] <= 8'h10 ;
			data[31612] <= 8'h10 ;
			data[31613] <= 8'h10 ;
			data[31614] <= 8'h10 ;
			data[31615] <= 8'h10 ;
			data[31616] <= 8'h10 ;
			data[31617] <= 8'h10 ;
			data[31618] <= 8'h10 ;
			data[31619] <= 8'h10 ;
			data[31620] <= 8'h10 ;
			data[31621] <= 8'h10 ;
			data[31622] <= 8'h10 ;
			data[31623] <= 8'h10 ;
			data[31624] <= 8'h10 ;
			data[31625] <= 8'h10 ;
			data[31626] <= 8'h10 ;
			data[31627] <= 8'h10 ;
			data[31628] <= 8'h10 ;
			data[31629] <= 8'h10 ;
			data[31630] <= 8'h10 ;
			data[31631] <= 8'h10 ;
			data[31632] <= 8'h10 ;
			data[31633] <= 8'h10 ;
			data[31634] <= 8'h10 ;
			data[31635] <= 8'h10 ;
			data[31636] <= 8'h10 ;
			data[31637] <= 8'h10 ;
			data[31638] <= 8'h10 ;
			data[31639] <= 8'h10 ;
			data[31640] <= 8'h10 ;
			data[31641] <= 8'h10 ;
			data[31642] <= 8'h10 ;
			data[31643] <= 8'h10 ;
			data[31644] <= 8'h10 ;
			data[31645] <= 8'h10 ;
			data[31646] <= 8'h10 ;
			data[31647] <= 8'h10 ;
			data[31648] <= 8'h10 ;
			data[31649] <= 8'h10 ;
			data[31650] <= 8'h10 ;
			data[31651] <= 8'h10 ;
			data[31652] <= 8'h10 ;
			data[31653] <= 8'h10 ;
			data[31654] <= 8'h10 ;
			data[31655] <= 8'h10 ;
			data[31656] <= 8'h10 ;
			data[31657] <= 8'h10 ;
			data[31658] <= 8'h10 ;
			data[31659] <= 8'h10 ;
			data[31660] <= 8'h10 ;
			data[31661] <= 8'h10 ;
			data[31662] <= 8'h10 ;
			data[31663] <= 8'h10 ;
			data[31664] <= 8'h10 ;
			data[31665] <= 8'h10 ;
			data[31666] <= 8'h10 ;
			data[31667] <= 8'h10 ;
			data[31668] <= 8'h10 ;
			data[31669] <= 8'h10 ;
			data[31670] <= 8'h10 ;
			data[31671] <= 8'h10 ;
			data[31672] <= 8'h10 ;
			data[31673] <= 8'h10 ;
			data[31674] <= 8'h10 ;
			data[31675] <= 8'h10 ;
			data[31676] <= 8'h10 ;
			data[31677] <= 8'h10 ;
			data[31678] <= 8'h10 ;
			data[31679] <= 8'h10 ;
			data[31680] <= 8'h10 ;
			data[31681] <= 8'h10 ;
			data[31682] <= 8'h10 ;
			data[31683] <= 8'h10 ;
			data[31684] <= 8'h10 ;
			data[31685] <= 8'h10 ;
			data[31686] <= 8'h10 ;
			data[31687] <= 8'h10 ;
			data[31688] <= 8'h10 ;
			data[31689] <= 8'h10 ;
			data[31690] <= 8'h10 ;
			data[31691] <= 8'h10 ;
			data[31692] <= 8'h10 ;
			data[31693] <= 8'h10 ;
			data[31694] <= 8'h10 ;
			data[31695] <= 8'h10 ;
			data[31696] <= 8'h10 ;
			data[31697] <= 8'h10 ;
			data[31698] <= 8'h10 ;
			data[31699] <= 8'h10 ;
			data[31700] <= 8'h10 ;
			data[31701] <= 8'h10 ;
			data[31702] <= 8'h10 ;
			data[31703] <= 8'h10 ;
			data[31704] <= 8'h10 ;
			data[31705] <= 8'h10 ;
			data[31706] <= 8'h10 ;
			data[31707] <= 8'h10 ;
			data[31708] <= 8'h10 ;
			data[31709] <= 8'h10 ;
			data[31710] <= 8'h10 ;
			data[31711] <= 8'h10 ;
			data[31712] <= 8'h10 ;
			data[31713] <= 8'h10 ;
			data[31714] <= 8'h10 ;
			data[31715] <= 8'h10 ;
			data[31716] <= 8'h10 ;
			data[31717] <= 8'h10 ;
			data[31718] <= 8'h10 ;
			data[31719] <= 8'h10 ;
			data[31720] <= 8'h10 ;
			data[31721] <= 8'h10 ;
			data[31722] <= 8'h10 ;
			data[31723] <= 8'h10 ;
			data[31724] <= 8'h10 ;
			data[31725] <= 8'h10 ;
			data[31726] <= 8'h10 ;
			data[31727] <= 8'h10 ;
			data[31728] <= 8'h10 ;
			data[31729] <= 8'h10 ;
			data[31730] <= 8'h10 ;
			data[31731] <= 8'h10 ;
			data[31732] <= 8'h10 ;
			data[31733] <= 8'h10 ;
			data[31734] <= 8'h10 ;
			data[31735] <= 8'h10 ;
			data[31736] <= 8'h10 ;
			data[31737] <= 8'h10 ;
			data[31738] <= 8'h10 ;
			data[31739] <= 8'h10 ;
			data[31740] <= 8'h10 ;
			data[31741] <= 8'h10 ;
			data[31742] <= 8'h10 ;
			data[31743] <= 8'h10 ;
			data[31744] <= 8'h10 ;
			data[31745] <= 8'h10 ;
			data[31746] <= 8'h10 ;
			data[31747] <= 8'h10 ;
			data[31748] <= 8'h10 ;
			data[31749] <= 8'h10 ;
			data[31750] <= 8'h10 ;
			data[31751] <= 8'h10 ;
			data[31752] <= 8'h10 ;
			data[31753] <= 8'h10 ;
			data[31754] <= 8'h10 ;
			data[31755] <= 8'h10 ;
			data[31756] <= 8'h10 ;
			data[31757] <= 8'h10 ;
			data[31758] <= 8'h10 ;
			data[31759] <= 8'h10 ;
			data[31760] <= 8'h10 ;
			data[31761] <= 8'h10 ;
			data[31762] <= 8'h10 ;
			data[31763] <= 8'h10 ;
			data[31764] <= 8'h10 ;
			data[31765] <= 8'h10 ;
			data[31766] <= 8'h10 ;
			data[31767] <= 8'h10 ;
			data[31768] <= 8'h10 ;
			data[31769] <= 8'h10 ;
			data[31770] <= 8'h10 ;
			data[31771] <= 8'h10 ;
			data[31772] <= 8'h10 ;
			data[31773] <= 8'h10 ;
			data[31774] <= 8'h10 ;
			data[31775] <= 8'h10 ;
			data[31776] <= 8'h10 ;
			data[31777] <= 8'h10 ;
			data[31778] <= 8'h10 ;
			data[31779] <= 8'h10 ;
			data[31780] <= 8'h10 ;
			data[31781] <= 8'h10 ;
			data[31782] <= 8'h10 ;
			data[31783] <= 8'h10 ;
			data[31784] <= 8'h10 ;
			data[31785] <= 8'h10 ;
			data[31786] <= 8'h10 ;
			data[31787] <= 8'h10 ;
			data[31788] <= 8'h10 ;
			data[31789] <= 8'h10 ;
			data[31790] <= 8'h10 ;
			data[31791] <= 8'h10 ;
			data[31792] <= 8'h10 ;
			data[31793] <= 8'h10 ;
			data[31794] <= 8'h10 ;
			data[31795] <= 8'h10 ;
			data[31796] <= 8'h10 ;
			data[31797] <= 8'h10 ;
			data[31798] <= 8'h10 ;
			data[31799] <= 8'h10 ;
			data[31800] <= 8'h10 ;
			data[31801] <= 8'h10 ;
			data[31802] <= 8'h10 ;
			data[31803] <= 8'h10 ;
			data[31804] <= 8'h10 ;
			data[31805] <= 8'h10 ;
			data[31806] <= 8'h10 ;
			data[31807] <= 8'h10 ;
			data[31808] <= 8'h10 ;
			data[31809] <= 8'h10 ;
			data[31810] <= 8'h10 ;
			data[31811] <= 8'h10 ;
			data[31812] <= 8'h10 ;
			data[31813] <= 8'h10 ;
			data[31814] <= 8'h10 ;
			data[31815] <= 8'h10 ;
			data[31816] <= 8'h10 ;
			data[31817] <= 8'h10 ;
			data[31818] <= 8'h10 ;
			data[31819] <= 8'h10 ;
			data[31820] <= 8'h10 ;
			data[31821] <= 8'h10 ;
			data[31822] <= 8'h10 ;
			data[31823] <= 8'h10 ;
			data[31824] <= 8'h10 ;
			data[31825] <= 8'h10 ;
			data[31826] <= 8'h10 ;
			data[31827] <= 8'h10 ;
			data[31828] <= 8'h10 ;
			data[31829] <= 8'h10 ;
			data[31830] <= 8'h10 ;
			data[31831] <= 8'h10 ;
			data[31832] <= 8'h10 ;
			data[31833] <= 8'h10 ;
			data[31834] <= 8'h10 ;
			data[31835] <= 8'h10 ;
			data[31836] <= 8'h10 ;
			data[31837] <= 8'h10 ;
			data[31838] <= 8'h10 ;
			data[31839] <= 8'h10 ;
			data[31840] <= 8'h10 ;
			data[31841] <= 8'h10 ;
			data[31842] <= 8'h10 ;
			data[31843] <= 8'h10 ;
			data[31844] <= 8'h10 ;
			data[31845] <= 8'h10 ;
			data[31846] <= 8'h10 ;
			data[31847] <= 8'h10 ;
			data[31848] <= 8'h10 ;
			data[31849] <= 8'h10 ;
			data[31850] <= 8'h10 ;
			data[31851] <= 8'h10 ;
			data[31852] <= 8'h10 ;
			data[31853] <= 8'h10 ;
			data[31854] <= 8'h10 ;
			data[31855] <= 8'h10 ;
			data[31856] <= 8'h10 ;
			data[31857] <= 8'h10 ;
			data[31858] <= 8'h10 ;
			data[31859] <= 8'h10 ;
			data[31860] <= 8'h10 ;
			data[31861] <= 8'h10 ;
			data[31862] <= 8'h10 ;
			data[31863] <= 8'h10 ;
			data[31864] <= 8'h10 ;
			data[31865] <= 8'h10 ;
			data[31866] <= 8'h10 ;
			data[31867] <= 8'h10 ;
			data[31868] <= 8'h10 ;
			data[31869] <= 8'h10 ;
			data[31870] <= 8'h10 ;
			data[31871] <= 8'h10 ;
			data[31872] <= 8'h10 ;
			data[31873] <= 8'h10 ;
			data[31874] <= 8'h10 ;
			data[31875] <= 8'h10 ;
			data[31876] <= 8'h10 ;
			data[31877] <= 8'h10 ;
			data[31878] <= 8'h10 ;
			data[31879] <= 8'h10 ;
			data[31880] <= 8'h10 ;
			data[31881] <= 8'h10 ;
			data[31882] <= 8'h10 ;
			data[31883] <= 8'h10 ;
			data[31884] <= 8'h10 ;
			data[31885] <= 8'h10 ;
			data[31886] <= 8'h10 ;
			data[31887] <= 8'h10 ;
			data[31888] <= 8'h10 ;
			data[31889] <= 8'h10 ;
			data[31890] <= 8'h10 ;
			data[31891] <= 8'h10 ;
			data[31892] <= 8'h10 ;
			data[31893] <= 8'h10 ;
			data[31894] <= 8'h10 ;
			data[31895] <= 8'h10 ;
			data[31896] <= 8'h10 ;
			data[31897] <= 8'h10 ;
			data[31898] <= 8'h10 ;
			data[31899] <= 8'h10 ;
			data[31900] <= 8'h10 ;
			data[31901] <= 8'h10 ;
			data[31902] <= 8'h10 ;
			data[31903] <= 8'h10 ;
			data[31904] <= 8'h10 ;
			data[31905] <= 8'h10 ;
			data[31906] <= 8'h10 ;
			data[31907] <= 8'h10 ;
			data[31908] <= 8'h10 ;
			data[31909] <= 8'h10 ;
			data[31910] <= 8'h10 ;
			data[31911] <= 8'h10 ;
			data[31912] <= 8'h10 ;
			data[31913] <= 8'h10 ;
			data[31914] <= 8'h10 ;
			data[31915] <= 8'h10 ;
			data[31916] <= 8'h10 ;
			data[31917] <= 8'h10 ;
			data[31918] <= 8'h10 ;
			data[31919] <= 8'h10 ;
			data[31920] <= 8'h10 ;
			data[31921] <= 8'h10 ;
			data[31922] <= 8'h10 ;
			data[31923] <= 8'h10 ;
			data[31924] <= 8'h10 ;
			data[31925] <= 8'h10 ;
			data[31926] <= 8'h10 ;
			data[31927] <= 8'h10 ;
			data[31928] <= 8'h10 ;
			data[31929] <= 8'h10 ;
			data[31930] <= 8'h10 ;
			data[31931] <= 8'h10 ;
			data[31932] <= 8'h10 ;
			data[31933] <= 8'h10 ;
			data[31934] <= 8'h10 ;
			data[31935] <= 8'h10 ;
			data[31936] <= 8'h10 ;
			data[31937] <= 8'h10 ;
			data[31938] <= 8'h10 ;
			data[31939] <= 8'h10 ;
			data[31940] <= 8'h10 ;
			data[31941] <= 8'h10 ;
			data[31942] <= 8'h10 ;
			data[31943] <= 8'h10 ;
			data[31944] <= 8'h10 ;
			data[31945] <= 8'h10 ;
			data[31946] <= 8'h10 ;
			data[31947] <= 8'h10 ;
			data[31948] <= 8'h10 ;
			data[31949] <= 8'h10 ;
			data[31950] <= 8'h10 ;
			data[31951] <= 8'h10 ;
			data[31952] <= 8'h10 ;
			data[31953] <= 8'h10 ;
			data[31954] <= 8'h10 ;
			data[31955] <= 8'h10 ;
			data[31956] <= 8'h10 ;
			data[31957] <= 8'h10 ;
			data[31958] <= 8'h10 ;
			data[31959] <= 8'h10 ;
			data[31960] <= 8'h10 ;
			data[31961] <= 8'h10 ;
			data[31962] <= 8'h10 ;
			data[31963] <= 8'h10 ;
			data[31964] <= 8'h10 ;
			data[31965] <= 8'h10 ;
			data[31966] <= 8'h10 ;
			data[31967] <= 8'h10 ;
			data[31968] <= 8'h10 ;
			data[31969] <= 8'h10 ;
			data[31970] <= 8'h10 ;
			data[31971] <= 8'h10 ;
			data[31972] <= 8'h10 ;
			data[31973] <= 8'h10 ;
			data[31974] <= 8'h10 ;
			data[31975] <= 8'h10 ;
			data[31976] <= 8'h10 ;
			data[31977] <= 8'h10 ;
			data[31978] <= 8'h10 ;
			data[31979] <= 8'h10 ;
			data[31980] <= 8'h10 ;
			data[31981] <= 8'h10 ;
			data[31982] <= 8'h10 ;
			data[31983] <= 8'h10 ;
			data[31984] <= 8'h10 ;
			data[31985] <= 8'h10 ;
			data[31986] <= 8'h10 ;
			data[31987] <= 8'h10 ;
			data[31988] <= 8'h10 ;
			data[31989] <= 8'h10 ;
			data[31990] <= 8'h10 ;
			data[31991] <= 8'h10 ;
			data[31992] <= 8'h10 ;
			data[31993] <= 8'h10 ;
			data[31994] <= 8'h10 ;
			data[31995] <= 8'h10 ;
			data[31996] <= 8'h10 ;
			data[31997] <= 8'h10 ;
			data[31998] <= 8'h10 ;
			data[31999] <= 8'h10 ;
			data[32000] <= 8'h10 ;
			data[32001] <= 8'h10 ;
			data[32002] <= 8'h10 ;
			data[32003] <= 8'h10 ;
			data[32004] <= 8'h10 ;
			data[32005] <= 8'h10 ;
			data[32006] <= 8'h10 ;
			data[32007] <= 8'h10 ;
			data[32008] <= 8'h10 ;
			data[32009] <= 8'h10 ;
			data[32010] <= 8'h10 ;
			data[32011] <= 8'h10 ;
			data[32012] <= 8'h10 ;
			data[32013] <= 8'h10 ;
			data[32014] <= 8'h10 ;
			data[32015] <= 8'h10 ;
			data[32016] <= 8'h10 ;
			data[32017] <= 8'h10 ;
			data[32018] <= 8'h10 ;
			data[32019] <= 8'h10 ;
			data[32020] <= 8'h10 ;
			data[32021] <= 8'h10 ;
			data[32022] <= 8'h10 ;
			data[32023] <= 8'h10 ;
			data[32024] <= 8'h10 ;
			data[32025] <= 8'h10 ;
			data[32026] <= 8'h10 ;
			data[32027] <= 8'h10 ;
			data[32028] <= 8'h10 ;
			data[32029] <= 8'h10 ;
			data[32030] <= 8'h10 ;
			data[32031] <= 8'h10 ;
			data[32032] <= 8'h10 ;
			data[32033] <= 8'h10 ;
			data[32034] <= 8'h10 ;
			data[32035] <= 8'h10 ;
			data[32036] <= 8'h10 ;
			data[32037] <= 8'h10 ;
			data[32038] <= 8'h10 ;
			data[32039] <= 8'h10 ;
			data[32040] <= 8'h10 ;
			data[32041] <= 8'h10 ;
			data[32042] <= 8'h10 ;
			data[32043] <= 8'h10 ;
			data[32044] <= 8'h10 ;
			data[32045] <= 8'h10 ;
			data[32046] <= 8'h10 ;
			data[32047] <= 8'h10 ;
			data[32048] <= 8'h10 ;
			data[32049] <= 8'h10 ;
			data[32050] <= 8'h10 ;
			data[32051] <= 8'h10 ;
			data[32052] <= 8'h10 ;
			data[32053] <= 8'h10 ;
			data[32054] <= 8'h10 ;
			data[32055] <= 8'h10 ;
			data[32056] <= 8'h10 ;
			data[32057] <= 8'h10 ;
			data[32058] <= 8'h10 ;
			data[32059] <= 8'h10 ;
			data[32060] <= 8'h10 ;
			data[32061] <= 8'h10 ;
			data[32062] <= 8'h10 ;
			data[32063] <= 8'h10 ;
			data[32064] <= 8'h10 ;
			data[32065] <= 8'h10 ;
			data[32066] <= 8'h10 ;
			data[32067] <= 8'h10 ;
			data[32068] <= 8'h10 ;
			data[32069] <= 8'h10 ;
			data[32070] <= 8'h10 ;
			data[32071] <= 8'h10 ;
			data[32072] <= 8'h10 ;
			data[32073] <= 8'h10 ;
			data[32074] <= 8'h10 ;
			data[32075] <= 8'h10 ;
			data[32076] <= 8'h10 ;
			data[32077] <= 8'h10 ;
			data[32078] <= 8'h10 ;
			data[32079] <= 8'h10 ;
			data[32080] <= 8'h10 ;
			data[32081] <= 8'h10 ;
			data[32082] <= 8'h10 ;
			data[32083] <= 8'h10 ;
			data[32084] <= 8'h10 ;
			data[32085] <= 8'h10 ;
			data[32086] <= 8'h10 ;
			data[32087] <= 8'h10 ;
			data[32088] <= 8'h10 ;
			data[32089] <= 8'h10 ;
			data[32090] <= 8'h10 ;
			data[32091] <= 8'h10 ;
			data[32092] <= 8'h10 ;
			data[32093] <= 8'h10 ;
			data[32094] <= 8'h10 ;
			data[32095] <= 8'h10 ;
			data[32096] <= 8'h10 ;
			data[32097] <= 8'h10 ;
			data[32098] <= 8'h10 ;
			data[32099] <= 8'h10 ;
			data[32100] <= 8'h10 ;
			data[32101] <= 8'h10 ;
			data[32102] <= 8'h10 ;
			data[32103] <= 8'h10 ;
			data[32104] <= 8'h10 ;
			data[32105] <= 8'h10 ;
			data[32106] <= 8'h10 ;
			data[32107] <= 8'h10 ;
			data[32108] <= 8'h10 ;
			data[32109] <= 8'h10 ;
			data[32110] <= 8'h10 ;
			data[32111] <= 8'h10 ;
			data[32112] <= 8'h10 ;
			data[32113] <= 8'h10 ;
			data[32114] <= 8'h10 ;
			data[32115] <= 8'h10 ;
			data[32116] <= 8'h10 ;
			data[32117] <= 8'h10 ;
			data[32118] <= 8'h10 ;
			data[32119] <= 8'h10 ;
			data[32120] <= 8'h10 ;
			data[32121] <= 8'h10 ;
			data[32122] <= 8'h10 ;
			data[32123] <= 8'h10 ;
			data[32124] <= 8'h10 ;
			data[32125] <= 8'h10 ;
			data[32126] <= 8'h10 ;
			data[32127] <= 8'h10 ;
			data[32128] <= 8'h10 ;
			data[32129] <= 8'h10 ;
			data[32130] <= 8'h10 ;
			data[32131] <= 8'h10 ;
			data[32132] <= 8'h10 ;
			data[32133] <= 8'h10 ;
			data[32134] <= 8'h10 ;
			data[32135] <= 8'h10 ;
			data[32136] <= 8'h10 ;
			data[32137] <= 8'h10 ;
			data[32138] <= 8'h10 ;
			data[32139] <= 8'h10 ;
			data[32140] <= 8'h10 ;
			data[32141] <= 8'h10 ;
			data[32142] <= 8'h10 ;
			data[32143] <= 8'h10 ;
			data[32144] <= 8'h10 ;
			data[32145] <= 8'h10 ;
			data[32146] <= 8'h10 ;
			data[32147] <= 8'h10 ;
			data[32148] <= 8'h10 ;
			data[32149] <= 8'h10 ;
			data[32150] <= 8'h10 ;
			data[32151] <= 8'h10 ;
			data[32152] <= 8'h10 ;
			data[32153] <= 8'h10 ;
			data[32154] <= 8'h10 ;
			data[32155] <= 8'h10 ;
			data[32156] <= 8'h10 ;
			data[32157] <= 8'h10 ;
			data[32158] <= 8'h10 ;
			data[32159] <= 8'h10 ;
			data[32160] <= 8'h10 ;
			data[32161] <= 8'h10 ;
			data[32162] <= 8'h10 ;
			data[32163] <= 8'h10 ;
			data[32164] <= 8'h10 ;
			data[32165] <= 8'h10 ;
			data[32166] <= 8'h10 ;
			data[32167] <= 8'h10 ;
			data[32168] <= 8'h10 ;
			data[32169] <= 8'h10 ;
			data[32170] <= 8'h10 ;
			data[32171] <= 8'h10 ;
			data[32172] <= 8'h10 ;
			data[32173] <= 8'h10 ;
			data[32174] <= 8'h10 ;
			data[32175] <= 8'h10 ;
			data[32176] <= 8'h10 ;
			data[32177] <= 8'h10 ;
			data[32178] <= 8'h10 ;
			data[32179] <= 8'h10 ;
			data[32180] <= 8'h10 ;
			data[32181] <= 8'h10 ;
			data[32182] <= 8'h10 ;
			data[32183] <= 8'h10 ;
			data[32184] <= 8'h10 ;
			data[32185] <= 8'h10 ;
			data[32186] <= 8'h10 ;
			data[32187] <= 8'h10 ;
			data[32188] <= 8'h10 ;
			data[32189] <= 8'h10 ;
			data[32190] <= 8'h10 ;
			data[32191] <= 8'h10 ;
			data[32192] <= 8'h10 ;
			data[32193] <= 8'h10 ;
			data[32194] <= 8'h10 ;
			data[32195] <= 8'h10 ;
			data[32196] <= 8'h10 ;
			data[32197] <= 8'h10 ;
			data[32198] <= 8'h10 ;
			data[32199] <= 8'h10 ;
			data[32200] <= 8'h10 ;
			data[32201] <= 8'h10 ;
			data[32202] <= 8'h10 ;
			data[32203] <= 8'h10 ;
			data[32204] <= 8'h10 ;
			data[32205] <= 8'h10 ;
			data[32206] <= 8'h10 ;
			data[32207] <= 8'h10 ;
			data[32208] <= 8'h10 ;
			data[32209] <= 8'h10 ;
			data[32210] <= 8'h10 ;
			data[32211] <= 8'h10 ;
			data[32212] <= 8'h10 ;
			data[32213] <= 8'h10 ;
			data[32214] <= 8'h10 ;
			data[32215] <= 8'h10 ;
			data[32216] <= 8'h10 ;
			data[32217] <= 8'h10 ;
			data[32218] <= 8'h10 ;
			data[32219] <= 8'h10 ;
			data[32220] <= 8'h10 ;
			data[32221] <= 8'h10 ;
			data[32222] <= 8'h10 ;
			data[32223] <= 8'h10 ;
			data[32224] <= 8'h10 ;
			data[32225] <= 8'h10 ;
			data[32226] <= 8'h10 ;
			data[32227] <= 8'h10 ;
			data[32228] <= 8'h10 ;
			data[32229] <= 8'h10 ;
			data[32230] <= 8'h10 ;
			data[32231] <= 8'h10 ;
			data[32232] <= 8'h10 ;
			data[32233] <= 8'h10 ;
			data[32234] <= 8'h10 ;
			data[32235] <= 8'h10 ;
			data[32236] <= 8'h10 ;
			data[32237] <= 8'h10 ;
			data[32238] <= 8'h10 ;
			data[32239] <= 8'h10 ;
			data[32240] <= 8'h10 ;
			data[32241] <= 8'h10 ;
			data[32242] <= 8'h10 ;
			data[32243] <= 8'h10 ;
			data[32244] <= 8'h10 ;
			data[32245] <= 8'h10 ;
			data[32246] <= 8'h10 ;
			data[32247] <= 8'h10 ;
			data[32248] <= 8'h10 ;
			data[32249] <= 8'h10 ;
			data[32250] <= 8'h10 ;
			data[32251] <= 8'h10 ;
			data[32252] <= 8'h10 ;
			data[32253] <= 8'h10 ;
			data[32254] <= 8'h10 ;
			data[32255] <= 8'h10 ;
			data[32256] <= 8'h10 ;
			data[32257] <= 8'h10 ;
			data[32258] <= 8'h10 ;
			data[32259] <= 8'h10 ;
			data[32260] <= 8'h10 ;
			data[32261] <= 8'h10 ;
			data[32262] <= 8'h10 ;
			data[32263] <= 8'h10 ;
			data[32264] <= 8'h10 ;
			data[32265] <= 8'h10 ;
			data[32266] <= 8'h10 ;
			data[32267] <= 8'h10 ;
			data[32268] <= 8'h10 ;
			data[32269] <= 8'h10 ;
			data[32270] <= 8'h10 ;
			data[32271] <= 8'h10 ;
			data[32272] <= 8'h10 ;
			data[32273] <= 8'h10 ;
			data[32274] <= 8'h10 ;
			data[32275] <= 8'h10 ;
			data[32276] <= 8'h10 ;
			data[32277] <= 8'h10 ;
			data[32278] <= 8'h10 ;
			data[32279] <= 8'h10 ;
			data[32280] <= 8'h10 ;
			data[32281] <= 8'h10 ;
			data[32282] <= 8'h10 ;
			data[32283] <= 8'h10 ;
			data[32284] <= 8'h10 ;
			data[32285] <= 8'h10 ;
			data[32286] <= 8'h10 ;
			data[32287] <= 8'h10 ;
			data[32288] <= 8'h10 ;
			data[32289] <= 8'h10 ;
			data[32290] <= 8'h10 ;
			data[32291] <= 8'h10 ;
			data[32292] <= 8'h10 ;
			data[32293] <= 8'h10 ;
			data[32294] <= 8'h10 ;
			data[32295] <= 8'h10 ;
			data[32296] <= 8'h10 ;
			data[32297] <= 8'h10 ;
			data[32298] <= 8'h10 ;
			data[32299] <= 8'h10 ;
			data[32300] <= 8'h10 ;
			data[32301] <= 8'h10 ;
			data[32302] <= 8'h10 ;
			data[32303] <= 8'h10 ;
			data[32304] <= 8'h10 ;
			data[32305] <= 8'h10 ;
			data[32306] <= 8'h10 ;
			data[32307] <= 8'h10 ;
			data[32308] <= 8'h10 ;
			data[32309] <= 8'h10 ;
			data[32310] <= 8'h10 ;
			data[32311] <= 8'h10 ;
			data[32312] <= 8'h10 ;
			data[32313] <= 8'h10 ;
			data[32314] <= 8'h10 ;
			data[32315] <= 8'h10 ;
			data[32316] <= 8'h10 ;
			data[32317] <= 8'h10 ;
			data[32318] <= 8'h10 ;
			data[32319] <= 8'h10 ;
			data[32320] <= 8'h10 ;
			data[32321] <= 8'h10 ;
			data[32322] <= 8'h10 ;
			data[32323] <= 8'h10 ;
			data[32324] <= 8'h10 ;
			data[32325] <= 8'h10 ;
			data[32326] <= 8'h10 ;
			data[32327] <= 8'h10 ;
			data[32328] <= 8'h10 ;
			data[32329] <= 8'h10 ;
			data[32330] <= 8'h10 ;
			data[32331] <= 8'h10 ;
			data[32332] <= 8'h10 ;
			data[32333] <= 8'h10 ;
			data[32334] <= 8'h10 ;
			data[32335] <= 8'h10 ;
			data[32336] <= 8'h10 ;
			data[32337] <= 8'h10 ;
			data[32338] <= 8'h10 ;
			data[32339] <= 8'h10 ;
			data[32340] <= 8'h10 ;
			data[32341] <= 8'h10 ;
			data[32342] <= 8'h10 ;
			data[32343] <= 8'h10 ;
			data[32344] <= 8'h10 ;
			data[32345] <= 8'h10 ;
			data[32346] <= 8'h10 ;
			data[32347] <= 8'h10 ;
			data[32348] <= 8'h10 ;
			data[32349] <= 8'h10 ;
			data[32350] <= 8'h10 ;
			data[32351] <= 8'h10 ;
			data[32352] <= 8'h10 ;
			data[32353] <= 8'h10 ;
			data[32354] <= 8'h10 ;
			data[32355] <= 8'h10 ;
			data[32356] <= 8'h10 ;
			data[32357] <= 8'h10 ;
			data[32358] <= 8'h10 ;
			data[32359] <= 8'h10 ;
			data[32360] <= 8'h10 ;
			data[32361] <= 8'h10 ;
			data[32362] <= 8'h10 ;
			data[32363] <= 8'h10 ;
			data[32364] <= 8'h10 ;
			data[32365] <= 8'h10 ;
			data[32366] <= 8'h10 ;
			data[32367] <= 8'h10 ;
			data[32368] <= 8'h10 ;
			data[32369] <= 8'h10 ;
			data[32370] <= 8'h10 ;
			data[32371] <= 8'h10 ;
			data[32372] <= 8'h10 ;
			data[32373] <= 8'h10 ;
			data[32374] <= 8'h10 ;
			data[32375] <= 8'h10 ;
			data[32376] <= 8'h10 ;
			data[32377] <= 8'h10 ;
			data[32378] <= 8'h10 ;
			data[32379] <= 8'h10 ;
			data[32380] <= 8'h10 ;
			data[32381] <= 8'h10 ;
			data[32382] <= 8'h10 ;
			data[32383] <= 8'h10 ;
			data[32384] <= 8'h10 ;
			data[32385] <= 8'h10 ;
			data[32386] <= 8'h10 ;
			data[32387] <= 8'h10 ;
			data[32388] <= 8'h10 ;
			data[32389] <= 8'h10 ;
			data[32390] <= 8'h10 ;
			data[32391] <= 8'h10 ;
			data[32392] <= 8'h10 ;
			data[32393] <= 8'h10 ;
			data[32394] <= 8'h10 ;
			data[32395] <= 8'h10 ;
			data[32396] <= 8'h10 ;
			data[32397] <= 8'h10 ;
			data[32398] <= 8'h10 ;
			data[32399] <= 8'h10 ;
			data[32400] <= 8'h10 ;
			data[32401] <= 8'h10 ;
			data[32402] <= 8'h10 ;
			data[32403] <= 8'h10 ;
			data[32404] <= 8'h10 ;
			data[32405] <= 8'h10 ;
			data[32406] <= 8'h10 ;
			data[32407] <= 8'h10 ;
			data[32408] <= 8'h10 ;
			data[32409] <= 8'h10 ;
			data[32410] <= 8'h10 ;
			data[32411] <= 8'h10 ;
			data[32412] <= 8'h10 ;
			data[32413] <= 8'h10 ;
			data[32414] <= 8'h10 ;
			data[32415] <= 8'h10 ;
			data[32416] <= 8'h10 ;
			data[32417] <= 8'h10 ;
			data[32418] <= 8'h10 ;
			data[32419] <= 8'h10 ;
			data[32420] <= 8'h10 ;
			data[32421] <= 8'h10 ;
			data[32422] <= 8'h10 ;
			data[32423] <= 8'h10 ;
			data[32424] <= 8'h10 ;
			data[32425] <= 8'h10 ;
			data[32426] <= 8'h10 ;
			data[32427] <= 8'h10 ;
			data[32428] <= 8'h10 ;
			data[32429] <= 8'h10 ;
			data[32430] <= 8'h10 ;
			data[32431] <= 8'h10 ;
			data[32432] <= 8'h10 ;
			data[32433] <= 8'h10 ;
			data[32434] <= 8'h10 ;
			data[32435] <= 8'h10 ;
			data[32436] <= 8'h10 ;
			data[32437] <= 8'h10 ;
			data[32438] <= 8'h10 ;
			data[32439] <= 8'h10 ;
			data[32440] <= 8'h10 ;
			data[32441] <= 8'h10 ;
			data[32442] <= 8'h10 ;
			data[32443] <= 8'h10 ;
			data[32444] <= 8'h10 ;
			data[32445] <= 8'h10 ;
			data[32446] <= 8'h10 ;
			data[32447] <= 8'h10 ;
			data[32448] <= 8'h10 ;
			data[32449] <= 8'h10 ;
			data[32450] <= 8'h10 ;
			data[32451] <= 8'h10 ;
			data[32452] <= 8'h10 ;
			data[32453] <= 8'h10 ;
			data[32454] <= 8'h10 ;
			data[32455] <= 8'h10 ;
			data[32456] <= 8'h10 ;
			data[32457] <= 8'h10 ;
			data[32458] <= 8'h10 ;
			data[32459] <= 8'h10 ;
			data[32460] <= 8'h10 ;
			data[32461] <= 8'h10 ;
			data[32462] <= 8'h10 ;
			data[32463] <= 8'h10 ;
			data[32464] <= 8'h10 ;
			data[32465] <= 8'h10 ;
			data[32466] <= 8'h10 ;
			data[32467] <= 8'h10 ;
			data[32468] <= 8'h10 ;
			data[32469] <= 8'h10 ;
			data[32470] <= 8'h10 ;
			data[32471] <= 8'h10 ;
			data[32472] <= 8'h10 ;
			data[32473] <= 8'h10 ;
			data[32474] <= 8'h10 ;
			data[32475] <= 8'h10 ;
			data[32476] <= 8'h10 ;
			data[32477] <= 8'h10 ;
			data[32478] <= 8'h10 ;
			data[32479] <= 8'h10 ;
			data[32480] <= 8'h10 ;
			data[32481] <= 8'h10 ;
			data[32482] <= 8'h10 ;
			data[32483] <= 8'h10 ;
			data[32484] <= 8'h10 ;
			data[32485] <= 8'h10 ;
			data[32486] <= 8'h10 ;
			data[32487] <= 8'h10 ;
			data[32488] <= 8'h10 ;
			data[32489] <= 8'h10 ;
			data[32490] <= 8'h10 ;
			data[32491] <= 8'h10 ;
			data[32492] <= 8'h10 ;
			data[32493] <= 8'h10 ;
			data[32494] <= 8'h10 ;
			data[32495] <= 8'h10 ;
			data[32496] <= 8'h10 ;
			data[32497] <= 8'h10 ;
			data[32498] <= 8'h10 ;
			data[32499] <= 8'h10 ;
			data[32500] <= 8'h10 ;
			data[32501] <= 8'h10 ;
			data[32502] <= 8'h10 ;
			data[32503] <= 8'h10 ;
			data[32504] <= 8'h10 ;
			data[32505] <= 8'h10 ;
			data[32506] <= 8'h10 ;
			data[32507] <= 8'h10 ;
			data[32508] <= 8'h10 ;
			data[32509] <= 8'h10 ;
			data[32510] <= 8'h10 ;
			data[32511] <= 8'h10 ;
			data[32512] <= 8'h10 ;
			data[32513] <= 8'h10 ;
			data[32514] <= 8'h10 ;
			data[32515] <= 8'h10 ;
			data[32516] <= 8'h10 ;
			data[32517] <= 8'h10 ;
			data[32518] <= 8'h10 ;
			data[32519] <= 8'h10 ;
			data[32520] <= 8'h10 ;
			data[32521] <= 8'h10 ;
			data[32522] <= 8'h10 ;
			data[32523] <= 8'h10 ;
			data[32524] <= 8'h10 ;
			data[32525] <= 8'h10 ;
			data[32526] <= 8'h10 ;
			data[32527] <= 8'h10 ;
			data[32528] <= 8'h10 ;
			data[32529] <= 8'h10 ;
			data[32530] <= 8'h10 ;
			data[32531] <= 8'h10 ;
			data[32532] <= 8'h10 ;
			data[32533] <= 8'h10 ;
			data[32534] <= 8'h10 ;
			data[32535] <= 8'h10 ;
			data[32536] <= 8'h10 ;
			data[32537] <= 8'h10 ;
			data[32538] <= 8'h10 ;
			data[32539] <= 8'h10 ;
			data[32540] <= 8'h10 ;
			data[32541] <= 8'h10 ;
			data[32542] <= 8'h10 ;
			data[32543] <= 8'h10 ;
			data[32544] <= 8'h10 ;
			data[32545] <= 8'h10 ;
			data[32546] <= 8'h10 ;
			data[32547] <= 8'h10 ;
			data[32548] <= 8'h10 ;
			data[32549] <= 8'h10 ;
			data[32550] <= 8'h10 ;
			data[32551] <= 8'h10 ;
			data[32552] <= 8'h10 ;
			data[32553] <= 8'h10 ;
			data[32554] <= 8'h10 ;
			data[32555] <= 8'h10 ;
			data[32556] <= 8'h10 ;
			data[32557] <= 8'h10 ;
			data[32558] <= 8'h10 ;
			data[32559] <= 8'h10 ;
			data[32560] <= 8'h10 ;
			data[32561] <= 8'h10 ;
			data[32562] <= 8'h10 ;
			data[32563] <= 8'h10 ;
			data[32564] <= 8'h10 ;
			data[32565] <= 8'h10 ;
			data[32566] <= 8'h10 ;
			data[32567] <= 8'h10 ;
			data[32568] <= 8'h10 ;
			data[32569] <= 8'h10 ;
			data[32570] <= 8'h10 ;
			data[32571] <= 8'h10 ;
			data[32572] <= 8'h10 ;
			data[32573] <= 8'h10 ;
			data[32574] <= 8'h10 ;
			data[32575] <= 8'h10 ;
			data[32576] <= 8'h10 ;
			data[32577] <= 8'h10 ;
			data[32578] <= 8'h10 ;
			data[32579] <= 8'h10 ;
			data[32580] <= 8'h10 ;
			data[32581] <= 8'h10 ;
			data[32582] <= 8'h10 ;
			data[32583] <= 8'h10 ;
			data[32584] <= 8'h10 ;
			data[32585] <= 8'h10 ;
			data[32586] <= 8'h10 ;
			data[32587] <= 8'h10 ;
			data[32588] <= 8'h10 ;
			data[32589] <= 8'h10 ;
			data[32590] <= 8'h10 ;
			data[32591] <= 8'h10 ;
			data[32592] <= 8'h10 ;
			data[32593] <= 8'h10 ;
			data[32594] <= 8'h10 ;
			data[32595] <= 8'h10 ;
			data[32596] <= 8'h10 ;
			data[32597] <= 8'h10 ;
			data[32598] <= 8'h10 ;
			data[32599] <= 8'h10 ;
			data[32600] <= 8'h10 ;
			data[32601] <= 8'h10 ;
			data[32602] <= 8'h10 ;
			data[32603] <= 8'h10 ;
			data[32604] <= 8'h10 ;
			data[32605] <= 8'h10 ;
			data[32606] <= 8'h10 ;
			data[32607] <= 8'h10 ;
			data[32608] <= 8'h10 ;
			data[32609] <= 8'h10 ;
			data[32610] <= 8'h10 ;
			data[32611] <= 8'h10 ;
			data[32612] <= 8'h10 ;
			data[32613] <= 8'h10 ;
			data[32614] <= 8'h10 ;
			data[32615] <= 8'h10 ;
			data[32616] <= 8'h10 ;
			data[32617] <= 8'h10 ;
			data[32618] <= 8'h10 ;
			data[32619] <= 8'h10 ;
			data[32620] <= 8'h10 ;
			data[32621] <= 8'h10 ;
			data[32622] <= 8'h10 ;
			data[32623] <= 8'h10 ;
			data[32624] <= 8'h10 ;
			data[32625] <= 8'h10 ;
			data[32626] <= 8'h10 ;
			data[32627] <= 8'h10 ;
			data[32628] <= 8'h10 ;
			data[32629] <= 8'h10 ;
			data[32630] <= 8'h10 ;
			data[32631] <= 8'h10 ;
			data[32632] <= 8'h10 ;
			data[32633] <= 8'h10 ;
			data[32634] <= 8'h10 ;
			data[32635] <= 8'h10 ;
			data[32636] <= 8'h10 ;
			data[32637] <= 8'h10 ;
			data[32638] <= 8'h10 ;
			data[32639] <= 8'h10 ;
			data[32640] <= 8'h10 ;
			data[32641] <= 8'h10 ;
			data[32642] <= 8'h10 ;
			data[32643] <= 8'h10 ;
			data[32644] <= 8'h10 ;
			data[32645] <= 8'h10 ;
			data[32646] <= 8'h10 ;
			data[32647] <= 8'h10 ;
			data[32648] <= 8'h10 ;
			data[32649] <= 8'h10 ;
			data[32650] <= 8'h10 ;
			data[32651] <= 8'h10 ;
			data[32652] <= 8'h10 ;
			data[32653] <= 8'h10 ;
			data[32654] <= 8'h10 ;
			data[32655] <= 8'h10 ;
			data[32656] <= 8'h10 ;
			data[32657] <= 8'h10 ;
			data[32658] <= 8'h10 ;
			data[32659] <= 8'h10 ;
			data[32660] <= 8'h10 ;
			data[32661] <= 8'h10 ;
			data[32662] <= 8'h10 ;
			data[32663] <= 8'h10 ;
			data[32664] <= 8'h10 ;
			data[32665] <= 8'h10 ;
			data[32666] <= 8'h10 ;
			data[32667] <= 8'h10 ;
			data[32668] <= 8'h10 ;
			data[32669] <= 8'h10 ;
			data[32670] <= 8'h10 ;
			data[32671] <= 8'h10 ;
			data[32672] <= 8'h10 ;
			data[32673] <= 8'h10 ;
			data[32674] <= 8'h10 ;
			data[32675] <= 8'h10 ;
			data[32676] <= 8'h10 ;
			data[32677] <= 8'h10 ;
			data[32678] <= 8'h10 ;
			data[32679] <= 8'h10 ;
			data[32680] <= 8'h10 ;
			data[32681] <= 8'h10 ;
			data[32682] <= 8'h10 ;
			data[32683] <= 8'h10 ;
			data[32684] <= 8'h10 ;
			data[32685] <= 8'h10 ;
			data[32686] <= 8'h10 ;
			data[32687] <= 8'h10 ;
			data[32688] <= 8'h10 ;
			data[32689] <= 8'h10 ;
			data[32690] <= 8'h10 ;
			data[32691] <= 8'h10 ;
			data[32692] <= 8'h10 ;
			data[32693] <= 8'h10 ;
			data[32694] <= 8'h10 ;
			data[32695] <= 8'h10 ;
			data[32696] <= 8'h10 ;
			data[32697] <= 8'h10 ;
			data[32698] <= 8'h10 ;
			data[32699] <= 8'h10 ;
			data[32700] <= 8'h10 ;
			data[32701] <= 8'h10 ;
			data[32702] <= 8'h10 ;
			data[32703] <= 8'h10 ;
			data[32704] <= 8'h10 ;
			data[32705] <= 8'h10 ;
			data[32706] <= 8'h10 ;
			data[32707] <= 8'h10 ;
			data[32708] <= 8'h10 ;
			data[32709] <= 8'h10 ;
			data[32710] <= 8'h10 ;
			data[32711] <= 8'h10 ;
			data[32712] <= 8'h10 ;
			data[32713] <= 8'h10 ;
			data[32714] <= 8'h10 ;
			data[32715] <= 8'h10 ;
			data[32716] <= 8'h10 ;
			data[32717] <= 8'h10 ;
			data[32718] <= 8'h10 ;
			data[32719] <= 8'h10 ;
			data[32720] <= 8'h10 ;
			data[32721] <= 8'h10 ;
			data[32722] <= 8'h10 ;
			data[32723] <= 8'h10 ;
			data[32724] <= 8'h10 ;
			data[32725] <= 8'h10 ;
			data[32726] <= 8'h10 ;
			data[32727] <= 8'h10 ;
			data[32728] <= 8'h10 ;
			data[32729] <= 8'h10 ;
			data[32730] <= 8'h10 ;
			data[32731] <= 8'h10 ;
			data[32732] <= 8'h10 ;
			data[32733] <= 8'h10 ;
			data[32734] <= 8'h10 ;
			data[32735] <= 8'h10 ;
			data[32736] <= 8'h10 ;
			data[32737] <= 8'h10 ;
			data[32738] <= 8'h10 ;
			data[32739] <= 8'h10 ;
			data[32740] <= 8'h10 ;
			data[32741] <= 8'h10 ;
			data[32742] <= 8'h10 ;
			data[32743] <= 8'h10 ;
			data[32744] <= 8'h10 ;
			data[32745] <= 8'h10 ;
			data[32746] <= 8'h10 ;
			data[32747] <= 8'h10 ;
			data[32748] <= 8'h10 ;
			data[32749] <= 8'h10 ;
			data[32750] <= 8'h10 ;
			data[32751] <= 8'h10 ;
			data[32752] <= 8'h10 ;
			data[32753] <= 8'h10 ;
			data[32754] <= 8'h10 ;
			data[32755] <= 8'h10 ;
			data[32756] <= 8'h10 ;
			data[32757] <= 8'h10 ;
			data[32758] <= 8'h10 ;
			data[32759] <= 8'h10 ;
			data[32760] <= 8'h10 ;
			data[32761] <= 8'h10 ;
			data[32762] <= 8'h10 ;
			data[32763] <= 8'h10 ;
			data[32764] <= 8'h10 ;
			data[32765] <= 8'h10 ;
			data[32766] <= 8'h10 ;
			data[32767] <= 8'h10 ;
			data[32768] <= 8'h10 ;
			data[32769] <= 8'h10 ;
			data[32770] <= 8'h10 ;
			data[32771] <= 8'h10 ;
			data[32772] <= 8'h10 ;
			data[32773] <= 8'h10 ;
			data[32774] <= 8'h10 ;
			data[32775] <= 8'h10 ;
			data[32776] <= 8'h10 ;
			data[32777] <= 8'h10 ;
			data[32778] <= 8'h10 ;
			data[32779] <= 8'h10 ;
			data[32780] <= 8'h10 ;
			data[32781] <= 8'h10 ;
			data[32782] <= 8'h10 ;
			data[32783] <= 8'h10 ;
			data[32784] <= 8'h10 ;
			data[32785] <= 8'h10 ;
			data[32786] <= 8'h10 ;
			data[32787] <= 8'h10 ;
			data[32788] <= 8'h10 ;
			data[32789] <= 8'h10 ;
			data[32790] <= 8'h10 ;
			data[32791] <= 8'h10 ;
			data[32792] <= 8'h10 ;
			data[32793] <= 8'h10 ;
			data[32794] <= 8'h10 ;
			data[32795] <= 8'h10 ;
			data[32796] <= 8'h10 ;
			data[32797] <= 8'h10 ;
			data[32798] <= 8'h10 ;
			data[32799] <= 8'h10 ;
			data[32800] <= 8'h10 ;
			data[32801] <= 8'h10 ;
			data[32802] <= 8'h10 ;
			data[32803] <= 8'h10 ;
			data[32804] <= 8'h10 ;
			data[32805] <= 8'h10 ;
			data[32806] <= 8'h10 ;
			data[32807] <= 8'h10 ;
			data[32808] <= 8'h10 ;
			data[32809] <= 8'h10 ;
			data[32810] <= 8'h10 ;
			data[32811] <= 8'h10 ;
			data[32812] <= 8'h10 ;
			data[32813] <= 8'h10 ;
			data[32814] <= 8'h10 ;
			data[32815] <= 8'h10 ;
			data[32816] <= 8'h10 ;
			data[32817] <= 8'h10 ;
			data[32818] <= 8'h10 ;
			data[32819] <= 8'h10 ;
			data[32820] <= 8'h10 ;
			data[32821] <= 8'h10 ;
			data[32822] <= 8'h10 ;
			data[32823] <= 8'h10 ;
			data[32824] <= 8'h10 ;
			data[32825] <= 8'h10 ;
			data[32826] <= 8'h10 ;
			data[32827] <= 8'h10 ;
			data[32828] <= 8'h10 ;
			data[32829] <= 8'h10 ;
			data[32830] <= 8'h10 ;
			data[32831] <= 8'h10 ;
			data[32832] <= 8'h10 ;
			data[32833] <= 8'h10 ;
			data[32834] <= 8'h10 ;
			data[32835] <= 8'h10 ;
			data[32836] <= 8'h10 ;
			data[32837] <= 8'h10 ;
			data[32838] <= 8'h10 ;
			data[32839] <= 8'h10 ;
			data[32840] <= 8'h10 ;
			data[32841] <= 8'h10 ;
			data[32842] <= 8'h10 ;
			data[32843] <= 8'h10 ;
			data[32844] <= 8'h10 ;
			data[32845] <= 8'h10 ;
			data[32846] <= 8'h10 ;
			data[32847] <= 8'h10 ;
			data[32848] <= 8'h10 ;
			data[32849] <= 8'h10 ;
			data[32850] <= 8'h10 ;
			data[32851] <= 8'h10 ;
			data[32852] <= 8'h10 ;
			data[32853] <= 8'h10 ;
			data[32854] <= 8'h10 ;
			data[32855] <= 8'h10 ;
			data[32856] <= 8'h10 ;
			data[32857] <= 8'h10 ;
			data[32858] <= 8'h10 ;
			data[32859] <= 8'h10 ;
			data[32860] <= 8'h10 ;
			data[32861] <= 8'h10 ;
			data[32862] <= 8'h10 ;
			data[32863] <= 8'h10 ;
			data[32864] <= 8'h10 ;
			data[32865] <= 8'h10 ;
			data[32866] <= 8'h10 ;
			data[32867] <= 8'h10 ;
			data[32868] <= 8'h10 ;
			data[32869] <= 8'h10 ;
			data[32870] <= 8'h10 ;
			data[32871] <= 8'h10 ;
			data[32872] <= 8'h10 ;
			data[32873] <= 8'h10 ;
			data[32874] <= 8'h10 ;
			data[32875] <= 8'h10 ;
			data[32876] <= 8'h10 ;
			data[32877] <= 8'h10 ;
			data[32878] <= 8'h10 ;
			data[32879] <= 8'h10 ;
			data[32880] <= 8'h10 ;
			data[32881] <= 8'h10 ;
			data[32882] <= 8'h10 ;
			data[32883] <= 8'h10 ;
			data[32884] <= 8'h10 ;
			data[32885] <= 8'h10 ;
			data[32886] <= 8'h10 ;
			data[32887] <= 8'h10 ;
			data[32888] <= 8'h10 ;
			data[32889] <= 8'h10 ;
			data[32890] <= 8'h10 ;
			data[32891] <= 8'h10 ;
			data[32892] <= 8'h10 ;
			data[32893] <= 8'h10 ;
			data[32894] <= 8'h10 ;
			data[32895] <= 8'h10 ;
			data[32896] <= 8'h10 ;
			data[32897] <= 8'h10 ;
			data[32898] <= 8'h10 ;
			data[32899] <= 8'h10 ;
			data[32900] <= 8'h10 ;
			data[32901] <= 8'h10 ;
			data[32902] <= 8'h10 ;
			data[32903] <= 8'h10 ;
			data[32904] <= 8'h10 ;
			data[32905] <= 8'h10 ;
			data[32906] <= 8'h10 ;
			data[32907] <= 8'h10 ;
			data[32908] <= 8'h10 ;
			data[32909] <= 8'h10 ;
			data[32910] <= 8'h10 ;
			data[32911] <= 8'h10 ;
			data[32912] <= 8'h10 ;
			data[32913] <= 8'h10 ;
			data[32914] <= 8'h10 ;
			data[32915] <= 8'h10 ;
			data[32916] <= 8'h10 ;
			data[32917] <= 8'h10 ;
			data[32918] <= 8'h10 ;
			data[32919] <= 8'h10 ;
			data[32920] <= 8'h10 ;
			data[32921] <= 8'h10 ;
			data[32922] <= 8'h10 ;
			data[32923] <= 8'h10 ;
			data[32924] <= 8'h10 ;
			data[32925] <= 8'h10 ;
			data[32926] <= 8'h10 ;
			data[32927] <= 8'h10 ;
			data[32928] <= 8'h10 ;
			data[32929] <= 8'h10 ;
			data[32930] <= 8'h10 ;
			data[32931] <= 8'h10 ;
			data[32932] <= 8'h10 ;
			data[32933] <= 8'h10 ;
			data[32934] <= 8'h10 ;
			data[32935] <= 8'h10 ;
			data[32936] <= 8'h10 ;
			data[32937] <= 8'h10 ;
			data[32938] <= 8'h10 ;
			data[32939] <= 8'h10 ;
			data[32940] <= 8'h10 ;
			data[32941] <= 8'h10 ;
			data[32942] <= 8'h10 ;
			data[32943] <= 8'h10 ;
			data[32944] <= 8'h10 ;
			data[32945] <= 8'h10 ;
			data[32946] <= 8'h10 ;
			data[32947] <= 8'h10 ;
			data[32948] <= 8'h10 ;
			data[32949] <= 8'h10 ;
			data[32950] <= 8'h10 ;
			data[32951] <= 8'h10 ;
			data[32952] <= 8'h10 ;
			data[32953] <= 8'h10 ;
			data[32954] <= 8'h10 ;
			data[32955] <= 8'h10 ;
			data[32956] <= 8'h10 ;
			data[32957] <= 8'h10 ;
			data[32958] <= 8'h10 ;
			data[32959] <= 8'h10 ;
			data[32960] <= 8'h10 ;
			data[32961] <= 8'h10 ;
			data[32962] <= 8'h10 ;
			data[32963] <= 8'h10 ;
			data[32964] <= 8'h10 ;
			data[32965] <= 8'h10 ;
			data[32966] <= 8'h10 ;
			data[32967] <= 8'h10 ;
			data[32968] <= 8'h10 ;
			data[32969] <= 8'h10 ;
			data[32970] <= 8'h10 ;
			data[32971] <= 8'h10 ;
			data[32972] <= 8'h10 ;
			data[32973] <= 8'h10 ;
			data[32974] <= 8'h10 ;
			data[32975] <= 8'h10 ;
			data[32976] <= 8'h10 ;
			data[32977] <= 8'h10 ;
			data[32978] <= 8'h10 ;
			data[32979] <= 8'h10 ;
			data[32980] <= 8'h10 ;
			data[32981] <= 8'h10 ;
			data[32982] <= 8'h10 ;
			data[32983] <= 8'h10 ;
			data[32984] <= 8'h10 ;
			data[32985] <= 8'h10 ;
			data[32986] <= 8'h10 ;
			data[32987] <= 8'h10 ;
			data[32988] <= 8'h10 ;
			data[32989] <= 8'h10 ;
			data[32990] <= 8'h10 ;
			data[32991] <= 8'h10 ;
			data[32992] <= 8'h10 ;
			data[32993] <= 8'h10 ;
			data[32994] <= 8'h10 ;
			data[32995] <= 8'h10 ;
			data[32996] <= 8'h10 ;
			data[32997] <= 8'h10 ;
			data[32998] <= 8'h10 ;
			data[32999] <= 8'h10 ;
			data[33000] <= 8'h10 ;
			data[33001] <= 8'h10 ;
			data[33002] <= 8'h10 ;
			data[33003] <= 8'h10 ;
			data[33004] <= 8'h10 ;
			data[33005] <= 8'h10 ;
			data[33006] <= 8'h10 ;
			data[33007] <= 8'h10 ;
			data[33008] <= 8'h10 ;
			data[33009] <= 8'h10 ;
			data[33010] <= 8'h10 ;
			data[33011] <= 8'h10 ;
			data[33012] <= 8'h10 ;
			data[33013] <= 8'h10 ;
			data[33014] <= 8'h10 ;
			data[33015] <= 8'h10 ;
			data[33016] <= 8'h10 ;
			data[33017] <= 8'h10 ;
			data[33018] <= 8'h10 ;
			data[33019] <= 8'h10 ;
			data[33020] <= 8'h10 ;
			data[33021] <= 8'h10 ;
			data[33022] <= 8'h10 ;
			data[33023] <= 8'h10 ;
			data[33024] <= 8'h10 ;
			data[33025] <= 8'h10 ;
			data[33026] <= 8'h10 ;
			data[33027] <= 8'h10 ;
			data[33028] <= 8'h10 ;
			data[33029] <= 8'h10 ;
			data[33030] <= 8'h10 ;
			data[33031] <= 8'h10 ;
			data[33032] <= 8'h10 ;
			data[33033] <= 8'h10 ;
			data[33034] <= 8'h10 ;
			data[33035] <= 8'h10 ;
			data[33036] <= 8'h10 ;
			data[33037] <= 8'h10 ;
			data[33038] <= 8'h10 ;
			data[33039] <= 8'h10 ;
			data[33040] <= 8'h10 ;
			data[33041] <= 8'h10 ;
			data[33042] <= 8'h10 ;
			data[33043] <= 8'h10 ;
			data[33044] <= 8'h10 ;
			data[33045] <= 8'h10 ;
			data[33046] <= 8'h10 ;
			data[33047] <= 8'h10 ;
			data[33048] <= 8'h10 ;
			data[33049] <= 8'h10 ;
			data[33050] <= 8'h10 ;
			data[33051] <= 8'h10 ;
			data[33052] <= 8'h10 ;
			data[33053] <= 8'h10 ;
			data[33054] <= 8'h10 ;
			data[33055] <= 8'h10 ;
			data[33056] <= 8'h10 ;
			data[33057] <= 8'h10 ;
			data[33058] <= 8'h10 ;
			data[33059] <= 8'h10 ;
			data[33060] <= 8'h10 ;
			data[33061] <= 8'h10 ;
			data[33062] <= 8'h10 ;
			data[33063] <= 8'h10 ;
			data[33064] <= 8'h10 ;
			data[33065] <= 8'h10 ;
			data[33066] <= 8'h10 ;
			data[33067] <= 8'h10 ;
			data[33068] <= 8'h10 ;
			data[33069] <= 8'h10 ;
			data[33070] <= 8'h10 ;
			data[33071] <= 8'h10 ;
			data[33072] <= 8'h10 ;
			data[33073] <= 8'h10 ;
			data[33074] <= 8'h10 ;
			data[33075] <= 8'h10 ;
			data[33076] <= 8'h10 ;
			data[33077] <= 8'h10 ;
			data[33078] <= 8'h10 ;
			data[33079] <= 8'h10 ;
			data[33080] <= 8'h10 ;
			data[33081] <= 8'h10 ;
			data[33082] <= 8'h10 ;
			data[33083] <= 8'h10 ;
			data[33084] <= 8'h10 ;
			data[33085] <= 8'h10 ;
			data[33086] <= 8'h10 ;
			data[33087] <= 8'h10 ;
			data[33088] <= 8'h10 ;
			data[33089] <= 8'h10 ;
			data[33090] <= 8'h10 ;
			data[33091] <= 8'h10 ;
			data[33092] <= 8'h10 ;
			data[33093] <= 8'h10 ;
			data[33094] <= 8'h10 ;
			data[33095] <= 8'h10 ;
			data[33096] <= 8'h10 ;
			data[33097] <= 8'h10 ;
			data[33098] <= 8'h10 ;
			data[33099] <= 8'h10 ;
			data[33100] <= 8'h10 ;
			data[33101] <= 8'h10 ;
			data[33102] <= 8'h10 ;
			data[33103] <= 8'h10 ;
			data[33104] <= 8'h10 ;
			data[33105] <= 8'h10 ;
			data[33106] <= 8'h10 ;
			data[33107] <= 8'h10 ;
			data[33108] <= 8'h10 ;
			data[33109] <= 8'h10 ;
			data[33110] <= 8'h10 ;
			data[33111] <= 8'h10 ;
			data[33112] <= 8'h10 ;
			data[33113] <= 8'h10 ;
			data[33114] <= 8'h10 ;
			data[33115] <= 8'h10 ;
			data[33116] <= 8'h10 ;
			data[33117] <= 8'h10 ;
			data[33118] <= 8'h10 ;
			data[33119] <= 8'h10 ;
			data[33120] <= 8'h10 ;
			data[33121] <= 8'h10 ;
			data[33122] <= 8'h10 ;
			data[33123] <= 8'h10 ;
			data[33124] <= 8'h10 ;
			data[33125] <= 8'h10 ;
			data[33126] <= 8'h10 ;
			data[33127] <= 8'h10 ;
			data[33128] <= 8'h10 ;
			data[33129] <= 8'h10 ;
			data[33130] <= 8'h10 ;
			data[33131] <= 8'h10 ;
			data[33132] <= 8'h10 ;
			data[33133] <= 8'h10 ;
			data[33134] <= 8'h10 ;
			data[33135] <= 8'h10 ;
			data[33136] <= 8'h10 ;
			data[33137] <= 8'h10 ;
			data[33138] <= 8'h10 ;
			data[33139] <= 8'h10 ;
			data[33140] <= 8'h10 ;
			data[33141] <= 8'h10 ;
			data[33142] <= 8'h10 ;
			data[33143] <= 8'h10 ;
			data[33144] <= 8'h10 ;
			data[33145] <= 8'h10 ;
			data[33146] <= 8'h10 ;
			data[33147] <= 8'h10 ;
			data[33148] <= 8'h10 ;
			data[33149] <= 8'h10 ;
			data[33150] <= 8'h10 ;
			data[33151] <= 8'h10 ;
			data[33152] <= 8'h10 ;
			data[33153] <= 8'h10 ;
			data[33154] <= 8'h10 ;
			data[33155] <= 8'h10 ;
			data[33156] <= 8'h10 ;
			data[33157] <= 8'h10 ;
			data[33158] <= 8'h10 ;
			data[33159] <= 8'h10 ;
			data[33160] <= 8'h10 ;
			data[33161] <= 8'h10 ;
			data[33162] <= 8'h10 ;
			data[33163] <= 8'h10 ;
			data[33164] <= 8'h10 ;
			data[33165] <= 8'h10 ;
			data[33166] <= 8'h10 ;
			data[33167] <= 8'h10 ;
			data[33168] <= 8'h10 ;
			data[33169] <= 8'h10 ;
			data[33170] <= 8'h10 ;
			data[33171] <= 8'h10 ;
			data[33172] <= 8'h10 ;
			data[33173] <= 8'h10 ;
			data[33174] <= 8'h10 ;
			data[33175] <= 8'h10 ;
			data[33176] <= 8'h10 ;
			data[33177] <= 8'h10 ;
			data[33178] <= 8'h10 ;
			data[33179] <= 8'h10 ;
			data[33180] <= 8'h10 ;
			data[33181] <= 8'h10 ;
			data[33182] <= 8'h10 ;
			data[33183] <= 8'h10 ;
			data[33184] <= 8'h10 ;
			data[33185] <= 8'h10 ;
			data[33186] <= 8'h10 ;
			data[33187] <= 8'h10 ;
			data[33188] <= 8'h10 ;
			data[33189] <= 8'h10 ;
			data[33190] <= 8'h10 ;
			data[33191] <= 8'h10 ;
			data[33192] <= 8'h10 ;
			data[33193] <= 8'h10 ;
			data[33194] <= 8'h10 ;
			data[33195] <= 8'h10 ;
			data[33196] <= 8'h10 ;
			data[33197] <= 8'h10 ;
			data[33198] <= 8'h10 ;
			data[33199] <= 8'h10 ;
			data[33200] <= 8'h10 ;
			data[33201] <= 8'h10 ;
			data[33202] <= 8'h10 ;
			data[33203] <= 8'h10 ;
			data[33204] <= 8'h10 ;
			data[33205] <= 8'h10 ;
			data[33206] <= 8'h10 ;
			data[33207] <= 8'h10 ;
			data[33208] <= 8'h10 ;
			data[33209] <= 8'h10 ;
			data[33210] <= 8'h10 ;
			data[33211] <= 8'h10 ;
			data[33212] <= 8'h10 ;
			data[33213] <= 8'h10 ;
			data[33214] <= 8'h10 ;
			data[33215] <= 8'h10 ;
			data[33216] <= 8'h10 ;
			data[33217] <= 8'h10 ;
			data[33218] <= 8'h10 ;
			data[33219] <= 8'h10 ;
			data[33220] <= 8'h10 ;
			data[33221] <= 8'h10 ;
			data[33222] <= 8'h10 ;
			data[33223] <= 8'h10 ;
			data[33224] <= 8'h10 ;
			data[33225] <= 8'h10 ;
			data[33226] <= 8'h10 ;
			data[33227] <= 8'h10 ;
			data[33228] <= 8'h10 ;
			data[33229] <= 8'h10 ;
			data[33230] <= 8'h10 ;
			data[33231] <= 8'h10 ;
			data[33232] <= 8'h10 ;
			data[33233] <= 8'h10 ;
			data[33234] <= 8'h10 ;
			data[33235] <= 8'h10 ;
			data[33236] <= 8'h10 ;
			data[33237] <= 8'h10 ;
			data[33238] <= 8'h10 ;
			data[33239] <= 8'h10 ;
			data[33240] <= 8'h10 ;
			data[33241] <= 8'h10 ;
			data[33242] <= 8'h10 ;
			data[33243] <= 8'h10 ;
			data[33244] <= 8'h10 ;
			data[33245] <= 8'h10 ;
			data[33246] <= 8'h10 ;
			data[33247] <= 8'h10 ;
			data[33248] <= 8'h10 ;
			data[33249] <= 8'h10 ;
			data[33250] <= 8'h10 ;
			data[33251] <= 8'h10 ;
			data[33252] <= 8'h10 ;
			data[33253] <= 8'h10 ;
			data[33254] <= 8'h10 ;
			data[33255] <= 8'h10 ;
			data[33256] <= 8'h10 ;
			data[33257] <= 8'h10 ;
			data[33258] <= 8'h10 ;
			data[33259] <= 8'h10 ;
			data[33260] <= 8'h10 ;
			data[33261] <= 8'h10 ;
			data[33262] <= 8'h10 ;
			data[33263] <= 8'h10 ;
			data[33264] <= 8'h10 ;
			data[33265] <= 8'h10 ;
			data[33266] <= 8'h10 ;
			data[33267] <= 8'h10 ;
			data[33268] <= 8'h10 ;
			data[33269] <= 8'h10 ;
			data[33270] <= 8'h10 ;
			data[33271] <= 8'h10 ;
			data[33272] <= 8'h10 ;
			data[33273] <= 8'h10 ;
			data[33274] <= 8'h10 ;
			data[33275] <= 8'h10 ;
			data[33276] <= 8'h10 ;
			data[33277] <= 8'h10 ;
			data[33278] <= 8'h10 ;
			data[33279] <= 8'h10 ;
			data[33280] <= 8'h10 ;
			data[33281] <= 8'h10 ;
			data[33282] <= 8'h10 ;
			data[33283] <= 8'h10 ;
			data[33284] <= 8'h10 ;
			data[33285] <= 8'h10 ;
			data[33286] <= 8'h10 ;
			data[33287] <= 8'h10 ;
			data[33288] <= 8'h10 ;
			data[33289] <= 8'h10 ;
			data[33290] <= 8'h10 ;
			data[33291] <= 8'h10 ;
			data[33292] <= 8'h10 ;
			data[33293] <= 8'h10 ;
			data[33294] <= 8'h10 ;
			data[33295] <= 8'h10 ;
			data[33296] <= 8'h10 ;
			data[33297] <= 8'h10 ;
			data[33298] <= 8'h10 ;
			data[33299] <= 8'h10 ;
			data[33300] <= 8'h10 ;
			data[33301] <= 8'h10 ;
			data[33302] <= 8'h10 ;
			data[33303] <= 8'h10 ;
			data[33304] <= 8'h10 ;
			data[33305] <= 8'h10 ;
			data[33306] <= 8'h10 ;
			data[33307] <= 8'h10 ;
			data[33308] <= 8'h10 ;
			data[33309] <= 8'h10 ;
			data[33310] <= 8'h10 ;
			data[33311] <= 8'h10 ;
			data[33312] <= 8'h10 ;
			data[33313] <= 8'h10 ;
			data[33314] <= 8'h10 ;
			data[33315] <= 8'h10 ;
			data[33316] <= 8'h10 ;
			data[33317] <= 8'h10 ;
			data[33318] <= 8'h10 ;
			data[33319] <= 8'h10 ;
			data[33320] <= 8'h10 ;
			data[33321] <= 8'h10 ;
			data[33322] <= 8'h10 ;
			data[33323] <= 8'h10 ;
			data[33324] <= 8'h10 ;
			data[33325] <= 8'h10 ;
			data[33326] <= 8'h10 ;
			data[33327] <= 8'h10 ;
			data[33328] <= 8'h10 ;
			data[33329] <= 8'h10 ;
			data[33330] <= 8'h10 ;
			data[33331] <= 8'h10 ;
			data[33332] <= 8'h10 ;
			data[33333] <= 8'h10 ;
			data[33334] <= 8'h10 ;
			data[33335] <= 8'h10 ;
			data[33336] <= 8'h10 ;
			data[33337] <= 8'h10 ;
			data[33338] <= 8'h10 ;
			data[33339] <= 8'h10 ;
			data[33340] <= 8'h10 ;
			data[33341] <= 8'h10 ;
			data[33342] <= 8'h10 ;
			data[33343] <= 8'h10 ;
			data[33344] <= 8'h10 ;
			data[33345] <= 8'h10 ;
			data[33346] <= 8'h10 ;
			data[33347] <= 8'h10 ;
			data[33348] <= 8'h10 ;
			data[33349] <= 8'h10 ;
			data[33350] <= 8'h10 ;
			data[33351] <= 8'h10 ;
			data[33352] <= 8'h10 ;
			data[33353] <= 8'h10 ;
			data[33354] <= 8'h10 ;
			data[33355] <= 8'h10 ;
			data[33356] <= 8'h10 ;
			data[33357] <= 8'h10 ;
			data[33358] <= 8'h10 ;
			data[33359] <= 8'h10 ;
			data[33360] <= 8'h10 ;
			data[33361] <= 8'h10 ;
			data[33362] <= 8'h10 ;
			data[33363] <= 8'h10 ;
			data[33364] <= 8'h10 ;
			data[33365] <= 8'h10 ;
			data[33366] <= 8'h10 ;
			data[33367] <= 8'h10 ;
			data[33368] <= 8'h10 ;
			data[33369] <= 8'h10 ;
			data[33370] <= 8'h10 ;
			data[33371] <= 8'h10 ;
			data[33372] <= 8'h10 ;
			data[33373] <= 8'h10 ;
			data[33374] <= 8'h10 ;
			data[33375] <= 8'h10 ;
			data[33376] <= 8'h10 ;
			data[33377] <= 8'h10 ;
			data[33378] <= 8'h10 ;
			data[33379] <= 8'h10 ;
			data[33380] <= 8'h10 ;
			data[33381] <= 8'h10 ;
			data[33382] <= 8'h10 ;
			data[33383] <= 8'h10 ;
			data[33384] <= 8'h10 ;
			data[33385] <= 8'h10 ;
			data[33386] <= 8'h10 ;
			data[33387] <= 8'h10 ;
			data[33388] <= 8'h10 ;
			data[33389] <= 8'h10 ;
			data[33390] <= 8'h10 ;
			data[33391] <= 8'h10 ;
			data[33392] <= 8'h10 ;
			data[33393] <= 8'h10 ;
			data[33394] <= 8'h10 ;
			data[33395] <= 8'h10 ;
			data[33396] <= 8'h10 ;
			data[33397] <= 8'h10 ;
			data[33398] <= 8'h10 ;
			data[33399] <= 8'h10 ;
			data[33400] <= 8'h10 ;
			data[33401] <= 8'h10 ;
			data[33402] <= 8'h10 ;
			data[33403] <= 8'h10 ;
			data[33404] <= 8'h10 ;
			data[33405] <= 8'h10 ;
			data[33406] <= 8'h10 ;
			data[33407] <= 8'h10 ;
			data[33408] <= 8'h10 ;
			data[33409] <= 8'h10 ;
			data[33410] <= 8'h10 ;
			data[33411] <= 8'h10 ;
			data[33412] <= 8'h10 ;
			data[33413] <= 8'h10 ;
			data[33414] <= 8'h10 ;
			data[33415] <= 8'h10 ;
			data[33416] <= 8'h10 ;
			data[33417] <= 8'h10 ;
			data[33418] <= 8'h10 ;
			data[33419] <= 8'h10 ;
			data[33420] <= 8'h10 ;
			data[33421] <= 8'h10 ;
			data[33422] <= 8'h10 ;
			data[33423] <= 8'h10 ;
			data[33424] <= 8'h10 ;
			data[33425] <= 8'h10 ;
			data[33426] <= 8'h10 ;
			data[33427] <= 8'h10 ;
			data[33428] <= 8'h10 ;
			data[33429] <= 8'h10 ;
			data[33430] <= 8'h10 ;
			data[33431] <= 8'h10 ;
			data[33432] <= 8'h10 ;
			data[33433] <= 8'h10 ;
			data[33434] <= 8'h10 ;
			data[33435] <= 8'h10 ;
			data[33436] <= 8'h10 ;
			data[33437] <= 8'h10 ;
			data[33438] <= 8'h10 ;
			data[33439] <= 8'h10 ;
			data[33440] <= 8'h10 ;
			data[33441] <= 8'h10 ;
			data[33442] <= 8'h10 ;
			data[33443] <= 8'h10 ;
			data[33444] <= 8'h10 ;
			data[33445] <= 8'h10 ;
			data[33446] <= 8'h10 ;
			data[33447] <= 8'h10 ;
			data[33448] <= 8'h10 ;
			data[33449] <= 8'h10 ;
			data[33450] <= 8'h10 ;
			data[33451] <= 8'h10 ;
			data[33452] <= 8'h10 ;
			data[33453] <= 8'h10 ;
			data[33454] <= 8'h10 ;
			data[33455] <= 8'h10 ;
			data[33456] <= 8'h10 ;
			data[33457] <= 8'h10 ;
			data[33458] <= 8'h10 ;
			data[33459] <= 8'h10 ;
			data[33460] <= 8'h10 ;
			data[33461] <= 8'h10 ;
			data[33462] <= 8'h10 ;
			data[33463] <= 8'h10 ;
			data[33464] <= 8'h10 ;
			data[33465] <= 8'h10 ;
			data[33466] <= 8'h10 ;
			data[33467] <= 8'h10 ;
			data[33468] <= 8'h10 ;
			data[33469] <= 8'h10 ;
			data[33470] <= 8'h10 ;
			data[33471] <= 8'h10 ;
			data[33472] <= 8'h10 ;
			data[33473] <= 8'h10 ;
			data[33474] <= 8'h10 ;
			data[33475] <= 8'h10 ;
			data[33476] <= 8'h10 ;
			data[33477] <= 8'h10 ;
			data[33478] <= 8'h10 ;
			data[33479] <= 8'h10 ;
			data[33480] <= 8'h10 ;
			data[33481] <= 8'h10 ;
			data[33482] <= 8'h10 ;
			data[33483] <= 8'h10 ;
			data[33484] <= 8'h10 ;
			data[33485] <= 8'h10 ;
			data[33486] <= 8'h10 ;
			data[33487] <= 8'h10 ;
			data[33488] <= 8'h10 ;
			data[33489] <= 8'h10 ;
			data[33490] <= 8'h10 ;
			data[33491] <= 8'h10 ;
			data[33492] <= 8'h10 ;
			data[33493] <= 8'h10 ;
			data[33494] <= 8'h10 ;
			data[33495] <= 8'h10 ;
			data[33496] <= 8'h10 ;
			data[33497] <= 8'h10 ;
			data[33498] <= 8'h10 ;
			data[33499] <= 8'h10 ;
			data[33500] <= 8'h10 ;
			data[33501] <= 8'h10 ;
			data[33502] <= 8'h10 ;
			data[33503] <= 8'h10 ;
			data[33504] <= 8'h10 ;
			data[33505] <= 8'h10 ;
			data[33506] <= 8'h10 ;
			data[33507] <= 8'h10 ;
			data[33508] <= 8'h10 ;
			data[33509] <= 8'h10 ;
			data[33510] <= 8'h10 ;
			data[33511] <= 8'h10 ;
			data[33512] <= 8'h10 ;
			data[33513] <= 8'h10 ;
			data[33514] <= 8'h10 ;
			data[33515] <= 8'h10 ;
			data[33516] <= 8'h10 ;
			data[33517] <= 8'h10 ;
			data[33518] <= 8'h10 ;
			data[33519] <= 8'h10 ;
			data[33520] <= 8'h10 ;
			data[33521] <= 8'h10 ;
			data[33522] <= 8'h10 ;
			data[33523] <= 8'h10 ;
			data[33524] <= 8'h10 ;
			data[33525] <= 8'h10 ;
			data[33526] <= 8'h10 ;
			data[33527] <= 8'h10 ;
			data[33528] <= 8'h10 ;
			data[33529] <= 8'h10 ;
			data[33530] <= 8'h10 ;
			data[33531] <= 8'h10 ;
			data[33532] <= 8'h10 ;
			data[33533] <= 8'h10 ;
			data[33534] <= 8'h10 ;
			data[33535] <= 8'h10 ;
			data[33536] <= 8'h10 ;
			data[33537] <= 8'h10 ;
			data[33538] <= 8'h10 ;
			data[33539] <= 8'h10 ;
			data[33540] <= 8'h10 ;
			data[33541] <= 8'h10 ;
			data[33542] <= 8'h10 ;
			data[33543] <= 8'h10 ;
			data[33544] <= 8'h10 ;
			data[33545] <= 8'h10 ;
			data[33546] <= 8'h10 ;
			data[33547] <= 8'h10 ;
			data[33548] <= 8'h10 ;
			data[33549] <= 8'h10 ;
			data[33550] <= 8'h10 ;
			data[33551] <= 8'h10 ;
			data[33552] <= 8'h10 ;
			data[33553] <= 8'h10 ;
			data[33554] <= 8'h10 ;
			data[33555] <= 8'h10 ;
			data[33556] <= 8'h10 ;
			data[33557] <= 8'h10 ;
			data[33558] <= 8'h10 ;
			data[33559] <= 8'h10 ;
			data[33560] <= 8'h10 ;
			data[33561] <= 8'h10 ;
			data[33562] <= 8'h10 ;
			data[33563] <= 8'h10 ;
			data[33564] <= 8'h10 ;
			data[33565] <= 8'h10 ;
			data[33566] <= 8'h10 ;
			data[33567] <= 8'h10 ;
			data[33568] <= 8'h10 ;
			data[33569] <= 8'h10 ;
			data[33570] <= 8'h10 ;
			data[33571] <= 8'h10 ;
			data[33572] <= 8'h10 ;
			data[33573] <= 8'h10 ;
			data[33574] <= 8'h10 ;
			data[33575] <= 8'h10 ;
			data[33576] <= 8'h10 ;
			data[33577] <= 8'h10 ;
			data[33578] <= 8'h10 ;
			data[33579] <= 8'h10 ;
			data[33580] <= 8'h10 ;
			data[33581] <= 8'h10 ;
			data[33582] <= 8'h10 ;
			data[33583] <= 8'h10 ;
			data[33584] <= 8'h10 ;
			data[33585] <= 8'h10 ;
			data[33586] <= 8'h10 ;
			data[33587] <= 8'h10 ;
			data[33588] <= 8'h10 ;
			data[33589] <= 8'h10 ;
			data[33590] <= 8'h10 ;
			data[33591] <= 8'h10 ;
			data[33592] <= 8'h10 ;
			data[33593] <= 8'h10 ;
			data[33594] <= 8'h10 ;
			data[33595] <= 8'h10 ;
			data[33596] <= 8'h10 ;
			data[33597] <= 8'h10 ;
			data[33598] <= 8'h10 ;
			data[33599] <= 8'h10 ;
			data[33600] <= 8'h10 ;
			data[33601] <= 8'h10 ;
			data[33602] <= 8'h10 ;
			data[33603] <= 8'h10 ;
			data[33604] <= 8'h10 ;
			data[33605] <= 8'h10 ;
			data[33606] <= 8'h10 ;
			data[33607] <= 8'h10 ;
			data[33608] <= 8'h10 ;
			data[33609] <= 8'h10 ;
			data[33610] <= 8'h10 ;
			data[33611] <= 8'h10 ;
			data[33612] <= 8'h10 ;
			data[33613] <= 8'h10 ;
			data[33614] <= 8'h10 ;
			data[33615] <= 8'h10 ;
			data[33616] <= 8'h10 ;
			data[33617] <= 8'h10 ;
			data[33618] <= 8'h10 ;
			data[33619] <= 8'h10 ;
			data[33620] <= 8'h10 ;
			data[33621] <= 8'h10 ;
			data[33622] <= 8'h10 ;
			data[33623] <= 8'h10 ;
			data[33624] <= 8'h10 ;
			data[33625] <= 8'h10 ;
			data[33626] <= 8'h10 ;
			data[33627] <= 8'h10 ;
			data[33628] <= 8'h10 ;
			data[33629] <= 8'h10 ;
			data[33630] <= 8'h10 ;
			data[33631] <= 8'h10 ;
			data[33632] <= 8'h10 ;
			data[33633] <= 8'h10 ;
			data[33634] <= 8'h10 ;
			data[33635] <= 8'h10 ;
			data[33636] <= 8'h10 ;
			data[33637] <= 8'h10 ;
			data[33638] <= 8'h10 ;
			data[33639] <= 8'h10 ;
			data[33640] <= 8'h10 ;
			data[33641] <= 8'h10 ;
			data[33642] <= 8'h10 ;
			data[33643] <= 8'h10 ;
			data[33644] <= 8'h10 ;
			data[33645] <= 8'h10 ;
			data[33646] <= 8'h10 ;
			data[33647] <= 8'h10 ;
			data[33648] <= 8'h10 ;
			data[33649] <= 8'h10 ;
			data[33650] <= 8'h10 ;
			data[33651] <= 8'h10 ;
			data[33652] <= 8'h10 ;
			data[33653] <= 8'h10 ;
			data[33654] <= 8'h10 ;
			data[33655] <= 8'h10 ;
			data[33656] <= 8'h10 ;
			data[33657] <= 8'h10 ;
			data[33658] <= 8'h10 ;
			data[33659] <= 8'h10 ;
			data[33660] <= 8'h10 ;
			data[33661] <= 8'h10 ;
			data[33662] <= 8'h10 ;
			data[33663] <= 8'h10 ;
			data[33664] <= 8'h10 ;
			data[33665] <= 8'h10 ;
			data[33666] <= 8'h10 ;
			data[33667] <= 8'h10 ;
			data[33668] <= 8'h10 ;
			data[33669] <= 8'h10 ;
			data[33670] <= 8'h10 ;
			data[33671] <= 8'h10 ;
			data[33672] <= 8'h10 ;
			data[33673] <= 8'h10 ;
			data[33674] <= 8'h10 ;
			data[33675] <= 8'h10 ;
			data[33676] <= 8'h10 ;
			data[33677] <= 8'h10 ;
			data[33678] <= 8'h10 ;
			data[33679] <= 8'h10 ;
			data[33680] <= 8'h10 ;
			data[33681] <= 8'h10 ;
			data[33682] <= 8'h10 ;
			data[33683] <= 8'h10 ;
			data[33684] <= 8'h10 ;
			data[33685] <= 8'h10 ;
			data[33686] <= 8'h10 ;
			data[33687] <= 8'h10 ;
			data[33688] <= 8'h10 ;
			data[33689] <= 8'h10 ;
			data[33690] <= 8'h10 ;
			data[33691] <= 8'h10 ;
			data[33692] <= 8'h10 ;
			data[33693] <= 8'h10 ;
			data[33694] <= 8'h10 ;
			data[33695] <= 8'h10 ;
			data[33696] <= 8'h10 ;
			data[33697] <= 8'h10 ;
			data[33698] <= 8'h10 ;
			data[33699] <= 8'h10 ;
			data[33700] <= 8'h10 ;
			data[33701] <= 8'h10 ;
			data[33702] <= 8'h10 ;
			data[33703] <= 8'h10 ;
			data[33704] <= 8'h10 ;
			data[33705] <= 8'h10 ;
			data[33706] <= 8'h10 ;
			data[33707] <= 8'h10 ;
			data[33708] <= 8'h10 ;
			data[33709] <= 8'h10 ;
			data[33710] <= 8'h10 ;
			data[33711] <= 8'h10 ;
			data[33712] <= 8'h10 ;
			data[33713] <= 8'h10 ;
			data[33714] <= 8'h10 ;
			data[33715] <= 8'h10 ;
			data[33716] <= 8'h10 ;
			data[33717] <= 8'h10 ;
			data[33718] <= 8'h10 ;
			data[33719] <= 8'h10 ;
			data[33720] <= 8'h10 ;
			data[33721] <= 8'h10 ;
			data[33722] <= 8'h10 ;
			data[33723] <= 8'h10 ;
			data[33724] <= 8'h10 ;
			data[33725] <= 8'h10 ;
			data[33726] <= 8'h10 ;
			data[33727] <= 8'h10 ;
			data[33728] <= 8'h10 ;
			data[33729] <= 8'h10 ;
			data[33730] <= 8'h10 ;
			data[33731] <= 8'h10 ;
			data[33732] <= 8'h10 ;
			data[33733] <= 8'h10 ;
			data[33734] <= 8'h10 ;
			data[33735] <= 8'h10 ;
			data[33736] <= 8'h10 ;
			data[33737] <= 8'h10 ;
			data[33738] <= 8'h10 ;
			data[33739] <= 8'h10 ;
			data[33740] <= 8'h10 ;
			data[33741] <= 8'h10 ;
			data[33742] <= 8'h10 ;
			data[33743] <= 8'h10 ;
			data[33744] <= 8'h10 ;
			data[33745] <= 8'h10 ;
			data[33746] <= 8'h10 ;
			data[33747] <= 8'h10 ;
			data[33748] <= 8'h10 ;
			data[33749] <= 8'h10 ;
			data[33750] <= 8'h10 ;
			data[33751] <= 8'h10 ;
			data[33752] <= 8'h10 ;
			data[33753] <= 8'h10 ;
			data[33754] <= 8'h10 ;
			data[33755] <= 8'h10 ;
			data[33756] <= 8'h10 ;
			data[33757] <= 8'h10 ;
			data[33758] <= 8'h10 ;
			data[33759] <= 8'h10 ;
			data[33760] <= 8'h10 ;
			data[33761] <= 8'h10 ;
			data[33762] <= 8'h10 ;
			data[33763] <= 8'h10 ;
			data[33764] <= 8'h10 ;
			data[33765] <= 8'h10 ;
			data[33766] <= 8'h10 ;
			data[33767] <= 8'h10 ;
			data[33768] <= 8'h10 ;
			data[33769] <= 8'h10 ;
			data[33770] <= 8'h10 ;
			data[33771] <= 8'h10 ;
			data[33772] <= 8'h10 ;
			data[33773] <= 8'h10 ;
			data[33774] <= 8'h10 ;
			data[33775] <= 8'h10 ;
			data[33776] <= 8'h10 ;
			data[33777] <= 8'h10 ;
			data[33778] <= 8'h10 ;
			data[33779] <= 8'h10 ;
			data[33780] <= 8'h10 ;
			data[33781] <= 8'h10 ;
			data[33782] <= 8'h10 ;
			data[33783] <= 8'h10 ;
			data[33784] <= 8'h10 ;
			data[33785] <= 8'h10 ;
			data[33786] <= 8'h10 ;
			data[33787] <= 8'h10 ;
			data[33788] <= 8'h10 ;
			data[33789] <= 8'h10 ;
			data[33790] <= 8'h10 ;
			data[33791] <= 8'h10 ;
			data[33792] <= 8'h10 ;
			data[33793] <= 8'h10 ;
			data[33794] <= 8'h10 ;
			data[33795] <= 8'h10 ;
			data[33796] <= 8'h10 ;
			data[33797] <= 8'h10 ;
			data[33798] <= 8'h10 ;
			data[33799] <= 8'h10 ;
			data[33800] <= 8'h10 ;
			data[33801] <= 8'h10 ;
			data[33802] <= 8'h10 ;
			data[33803] <= 8'h10 ;
			data[33804] <= 8'h10 ;
			data[33805] <= 8'h10 ;
			data[33806] <= 8'h10 ;
			data[33807] <= 8'h10 ;
			data[33808] <= 8'h10 ;
			data[33809] <= 8'h10 ;
			data[33810] <= 8'h10 ;
			data[33811] <= 8'h10 ;
			data[33812] <= 8'h10 ;
			data[33813] <= 8'h10 ;
			data[33814] <= 8'h10 ;
			data[33815] <= 8'h10 ;
			data[33816] <= 8'h10 ;
			data[33817] <= 8'h10 ;
			data[33818] <= 8'h10 ;
			data[33819] <= 8'h10 ;
			data[33820] <= 8'h10 ;
			data[33821] <= 8'h10 ;
			data[33822] <= 8'h10 ;
			data[33823] <= 8'h10 ;
			data[33824] <= 8'h10 ;
			data[33825] <= 8'h10 ;
			data[33826] <= 8'h10 ;
			data[33827] <= 8'h10 ;
			data[33828] <= 8'h10 ;
			data[33829] <= 8'h10 ;
			data[33830] <= 8'h10 ;
			data[33831] <= 8'h10 ;
			data[33832] <= 8'h10 ;
			data[33833] <= 8'h10 ;
			data[33834] <= 8'h10 ;
			data[33835] <= 8'h10 ;
			data[33836] <= 8'h10 ;
			data[33837] <= 8'h10 ;
			data[33838] <= 8'h10 ;
			data[33839] <= 8'h10 ;
			data[33840] <= 8'h10 ;
			data[33841] <= 8'h10 ;
			data[33842] <= 8'h10 ;
			data[33843] <= 8'h10 ;
			data[33844] <= 8'h10 ;
			data[33845] <= 8'h10 ;
			data[33846] <= 8'h10 ;
			data[33847] <= 8'h10 ;
			data[33848] <= 8'h10 ;
			data[33849] <= 8'h10 ;
			data[33850] <= 8'h10 ;
			data[33851] <= 8'h10 ;
			data[33852] <= 8'h10 ;
			data[33853] <= 8'h10 ;
			data[33854] <= 8'h10 ;
			data[33855] <= 8'h10 ;
			data[33856] <= 8'h10 ;
			data[33857] <= 8'h10 ;
			data[33858] <= 8'h10 ;
			data[33859] <= 8'h10 ;
			data[33860] <= 8'h10 ;
			data[33861] <= 8'h10 ;
			data[33862] <= 8'h10 ;
			data[33863] <= 8'h10 ;
			data[33864] <= 8'h10 ;
			data[33865] <= 8'h10 ;
			data[33866] <= 8'h10 ;
			data[33867] <= 8'h10 ;
			data[33868] <= 8'h10 ;
			data[33869] <= 8'h10 ;
			data[33870] <= 8'h10 ;
			data[33871] <= 8'h10 ;
			data[33872] <= 8'h10 ;
			data[33873] <= 8'h10 ;
			data[33874] <= 8'h10 ;
			data[33875] <= 8'h10 ;
			data[33876] <= 8'h10 ;
			data[33877] <= 8'h10 ;
			data[33878] <= 8'h10 ;
			data[33879] <= 8'h10 ;
			data[33880] <= 8'h10 ;
			data[33881] <= 8'h10 ;
			data[33882] <= 8'h10 ;
			data[33883] <= 8'h10 ;
			data[33884] <= 8'h10 ;
			data[33885] <= 8'h10 ;
			data[33886] <= 8'h10 ;
			data[33887] <= 8'h10 ;
			data[33888] <= 8'h10 ;
			data[33889] <= 8'h10 ;
			data[33890] <= 8'h10 ;
			data[33891] <= 8'h10 ;
			data[33892] <= 8'h10 ;
			data[33893] <= 8'h10 ;
			data[33894] <= 8'h10 ;
			data[33895] <= 8'h10 ;
			data[33896] <= 8'h10 ;
			data[33897] <= 8'h10 ;
			data[33898] <= 8'h10 ;
			data[33899] <= 8'h10 ;
			data[33900] <= 8'h10 ;
			data[33901] <= 8'h10 ;
			data[33902] <= 8'h10 ;
			data[33903] <= 8'h10 ;
			data[33904] <= 8'h10 ;
			data[33905] <= 8'h10 ;
			data[33906] <= 8'h10 ;
			data[33907] <= 8'h10 ;
			data[33908] <= 8'h10 ;
			data[33909] <= 8'h10 ;
			data[33910] <= 8'h10 ;
			data[33911] <= 8'h10 ;
			data[33912] <= 8'h10 ;
			data[33913] <= 8'h10 ;
			data[33914] <= 8'h10 ;
			data[33915] <= 8'h10 ;
			data[33916] <= 8'h10 ;
			data[33917] <= 8'h10 ;
			data[33918] <= 8'h10 ;
			data[33919] <= 8'h10 ;
			data[33920] <= 8'h10 ;
			data[33921] <= 8'h10 ;
			data[33922] <= 8'h10 ;
			data[33923] <= 8'h10 ;
			data[33924] <= 8'h10 ;
			data[33925] <= 8'h10 ;
			data[33926] <= 8'h10 ;
			data[33927] <= 8'h10 ;
			data[33928] <= 8'h10 ;
			data[33929] <= 8'h10 ;
			data[33930] <= 8'h10 ;
			data[33931] <= 8'h10 ;
			data[33932] <= 8'h10 ;
			data[33933] <= 8'h10 ;
			data[33934] <= 8'h10 ;
			data[33935] <= 8'h10 ;
			data[33936] <= 8'h10 ;
			data[33937] <= 8'h10 ;
			data[33938] <= 8'h10 ;
			data[33939] <= 8'h10 ;
			data[33940] <= 8'h10 ;
			data[33941] <= 8'h10 ;
			data[33942] <= 8'h10 ;
			data[33943] <= 8'h10 ;
			data[33944] <= 8'h10 ;
			data[33945] <= 8'h10 ;
			data[33946] <= 8'h10 ;
			data[33947] <= 8'h10 ;
			data[33948] <= 8'h10 ;
			data[33949] <= 8'h10 ;
			data[33950] <= 8'h10 ;
			data[33951] <= 8'h10 ;
			data[33952] <= 8'h10 ;
			data[33953] <= 8'h10 ;
			data[33954] <= 8'h10 ;
			data[33955] <= 8'h10 ;
			data[33956] <= 8'h10 ;
			data[33957] <= 8'h10 ;
			data[33958] <= 8'h10 ;
			data[33959] <= 8'h10 ;
			data[33960] <= 8'h10 ;
			data[33961] <= 8'h10 ;
			data[33962] <= 8'h10 ;
			data[33963] <= 8'h10 ;
			data[33964] <= 8'h10 ;
			data[33965] <= 8'h10 ;
			data[33966] <= 8'h10 ;
			data[33967] <= 8'h10 ;
			data[33968] <= 8'h10 ;
			data[33969] <= 8'h10 ;
			data[33970] <= 8'h10 ;
			data[33971] <= 8'h10 ;
			data[33972] <= 8'h10 ;
			data[33973] <= 8'h10 ;
			data[33974] <= 8'h10 ;
			data[33975] <= 8'h10 ;
			data[33976] <= 8'h10 ;
			data[33977] <= 8'h10 ;
			data[33978] <= 8'h10 ;
			data[33979] <= 8'h10 ;
			data[33980] <= 8'h10 ;
			data[33981] <= 8'h10 ;
			data[33982] <= 8'h10 ;
			data[33983] <= 8'h10 ;
			data[33984] <= 8'h10 ;
			data[33985] <= 8'h10 ;
			data[33986] <= 8'h10 ;
			data[33987] <= 8'h10 ;
			data[33988] <= 8'h10 ;
			data[33989] <= 8'h10 ;
			data[33990] <= 8'h10 ;
			data[33991] <= 8'h10 ;
			data[33992] <= 8'h10 ;
			data[33993] <= 8'h10 ;
			data[33994] <= 8'h10 ;
			data[33995] <= 8'h10 ;
			data[33996] <= 8'h10 ;
			data[33997] <= 8'h10 ;
			data[33998] <= 8'h10 ;
			data[33999] <= 8'h10 ;
			data[34000] <= 8'h10 ;
			data[34001] <= 8'h10 ;
			data[34002] <= 8'h10 ;
			data[34003] <= 8'h10 ;
			data[34004] <= 8'h10 ;
			data[34005] <= 8'h10 ;
			data[34006] <= 8'h10 ;
			data[34007] <= 8'h10 ;
			data[34008] <= 8'h10 ;
			data[34009] <= 8'h10 ;
			data[34010] <= 8'h10 ;
			data[34011] <= 8'h10 ;
			data[34012] <= 8'h10 ;
			data[34013] <= 8'h10 ;
			data[34014] <= 8'h10 ;
			data[34015] <= 8'h10 ;
			data[34016] <= 8'h10 ;
			data[34017] <= 8'h10 ;
			data[34018] <= 8'h10 ;
			data[34019] <= 8'h10 ;
			data[34020] <= 8'h10 ;
			data[34021] <= 8'h10 ;
			data[34022] <= 8'h10 ;
			data[34023] <= 8'h10 ;
			data[34024] <= 8'h10 ;
			data[34025] <= 8'h10 ;
			data[34026] <= 8'h10 ;
			data[34027] <= 8'h10 ;
			data[34028] <= 8'h10 ;
			data[34029] <= 8'h10 ;
			data[34030] <= 8'h10 ;
			data[34031] <= 8'h10 ;
			data[34032] <= 8'h10 ;
			data[34033] <= 8'h10 ;
			data[34034] <= 8'h10 ;
			data[34035] <= 8'h10 ;
			data[34036] <= 8'h10 ;
			data[34037] <= 8'h10 ;
			data[34038] <= 8'h10 ;
			data[34039] <= 8'h10 ;
			data[34040] <= 8'h10 ;
			data[34041] <= 8'h10 ;
			data[34042] <= 8'h10 ;
			data[34043] <= 8'h10 ;
			data[34044] <= 8'h10 ;
			data[34045] <= 8'h10 ;
			data[34046] <= 8'h10 ;
			data[34047] <= 8'h10 ;
			data[34048] <= 8'h10 ;
			data[34049] <= 8'h10 ;
			data[34050] <= 8'h10 ;
			data[34051] <= 8'h10 ;
			data[34052] <= 8'h10 ;
			data[34053] <= 8'h10 ;
			data[34054] <= 8'h10 ;
			data[34055] <= 8'h10 ;
			data[34056] <= 8'h10 ;
			data[34057] <= 8'h10 ;
			data[34058] <= 8'h10 ;
			data[34059] <= 8'h10 ;
			data[34060] <= 8'h10 ;
			data[34061] <= 8'h10 ;
			data[34062] <= 8'h10 ;
			data[34063] <= 8'h10 ;
			data[34064] <= 8'h10 ;
			data[34065] <= 8'h10 ;
			data[34066] <= 8'h10 ;
			data[34067] <= 8'h10 ;
			data[34068] <= 8'h10 ;
			data[34069] <= 8'h10 ;
			data[34070] <= 8'h10 ;
			data[34071] <= 8'h10 ;
			data[34072] <= 8'h10 ;
			data[34073] <= 8'h10 ;
			data[34074] <= 8'h10 ;
			data[34075] <= 8'h10 ;
			data[34076] <= 8'h10 ;
			data[34077] <= 8'h10 ;
			data[34078] <= 8'h10 ;
			data[34079] <= 8'h10 ;
			data[34080] <= 8'h10 ;
			data[34081] <= 8'h10 ;
			data[34082] <= 8'h10 ;
			data[34083] <= 8'h10 ;
			data[34084] <= 8'h10 ;
			data[34085] <= 8'h10 ;
			data[34086] <= 8'h10 ;
			data[34087] <= 8'h10 ;
			data[34088] <= 8'h10 ;
			data[34089] <= 8'h10 ;
			data[34090] <= 8'h10 ;
			data[34091] <= 8'h10 ;
			data[34092] <= 8'h10 ;
			data[34093] <= 8'h10 ;
			data[34094] <= 8'h10 ;
			data[34095] <= 8'h10 ;
			data[34096] <= 8'h10 ;
			data[34097] <= 8'h10 ;
			data[34098] <= 8'h10 ;
			data[34099] <= 8'h10 ;
			data[34100] <= 8'h10 ;
			data[34101] <= 8'h10 ;
			data[34102] <= 8'h10 ;
			data[34103] <= 8'h10 ;
			data[34104] <= 8'h10 ;
			data[34105] <= 8'h10 ;
			data[34106] <= 8'h10 ;
			data[34107] <= 8'h10 ;
			data[34108] <= 8'h10 ;
			data[34109] <= 8'h10 ;
			data[34110] <= 8'h10 ;
			data[34111] <= 8'h10 ;
			data[34112] <= 8'h10 ;
			data[34113] <= 8'h10 ;
			data[34114] <= 8'h10 ;
			data[34115] <= 8'h10 ;
			data[34116] <= 8'h10 ;
			data[34117] <= 8'h10 ;
			data[34118] <= 8'h10 ;
			data[34119] <= 8'h10 ;
			data[34120] <= 8'h10 ;
			data[34121] <= 8'h10 ;
			data[34122] <= 8'h10 ;
			data[34123] <= 8'h10 ;
			data[34124] <= 8'h10 ;
			data[34125] <= 8'h10 ;
			data[34126] <= 8'h10 ;
			data[34127] <= 8'h10 ;
			data[34128] <= 8'h10 ;
			data[34129] <= 8'h10 ;
			data[34130] <= 8'h10 ;
			data[34131] <= 8'h10 ;
			data[34132] <= 8'h10 ;
			data[34133] <= 8'h10 ;
			data[34134] <= 8'h10 ;
			data[34135] <= 8'h10 ;
			data[34136] <= 8'h10 ;
			data[34137] <= 8'h10 ;
			data[34138] <= 8'h10 ;
			data[34139] <= 8'h10 ;
			data[34140] <= 8'h10 ;
			data[34141] <= 8'h10 ;
			data[34142] <= 8'h10 ;
			data[34143] <= 8'h10 ;
			data[34144] <= 8'h10 ;
			data[34145] <= 8'h10 ;
			data[34146] <= 8'h10 ;
			data[34147] <= 8'h10 ;
			data[34148] <= 8'h10 ;
			data[34149] <= 8'h10 ;
			data[34150] <= 8'h10 ;
			data[34151] <= 8'h10 ;
			data[34152] <= 8'h10 ;
			data[34153] <= 8'h10 ;
			data[34154] <= 8'h10 ;
			data[34155] <= 8'h10 ;
			data[34156] <= 8'h10 ;
			data[34157] <= 8'h10 ;
			data[34158] <= 8'h10 ;
			data[34159] <= 8'h10 ;
			data[34160] <= 8'h10 ;
			data[34161] <= 8'h10 ;
			data[34162] <= 8'h10 ;
			data[34163] <= 8'h10 ;
			data[34164] <= 8'h10 ;
			data[34165] <= 8'h10 ;
			data[34166] <= 8'h10 ;
			data[34167] <= 8'h10 ;
			data[34168] <= 8'h10 ;
			data[34169] <= 8'h10 ;
			data[34170] <= 8'h10 ;
			data[34171] <= 8'h10 ;
			data[34172] <= 8'h10 ;
			data[34173] <= 8'h10 ;
			data[34174] <= 8'h10 ;
			data[34175] <= 8'h10 ;
			data[34176] <= 8'h10 ;
			data[34177] <= 8'h10 ;
			data[34178] <= 8'h10 ;
			data[34179] <= 8'h10 ;
			data[34180] <= 8'h10 ;
			data[34181] <= 8'h10 ;
			data[34182] <= 8'h10 ;
			data[34183] <= 8'h10 ;
			data[34184] <= 8'h10 ;
			data[34185] <= 8'h10 ;
			data[34186] <= 8'h10 ;
			data[34187] <= 8'h10 ;
			data[34188] <= 8'h10 ;
			data[34189] <= 8'h10 ;
			data[34190] <= 8'h10 ;
			data[34191] <= 8'h10 ;
			data[34192] <= 8'h10 ;
			data[34193] <= 8'h10 ;
			data[34194] <= 8'h10 ;
			data[34195] <= 8'h10 ;
			data[34196] <= 8'h10 ;
			data[34197] <= 8'h10 ;
			data[34198] <= 8'h10 ;
			data[34199] <= 8'h10 ;
			data[34200] <= 8'h10 ;
			data[34201] <= 8'h10 ;
			data[34202] <= 8'h10 ;
			data[34203] <= 8'h10 ;
			data[34204] <= 8'h10 ;
			data[34205] <= 8'h10 ;
			data[34206] <= 8'h10 ;
			data[34207] <= 8'h10 ;
			data[34208] <= 8'h10 ;
			data[34209] <= 8'h10 ;
			data[34210] <= 8'h10 ;
			data[34211] <= 8'h10 ;
			data[34212] <= 8'h10 ;
			data[34213] <= 8'h10 ;
			data[34214] <= 8'h10 ;
			data[34215] <= 8'h10 ;
			data[34216] <= 8'h10 ;
			data[34217] <= 8'h10 ;
			data[34218] <= 8'h10 ;
			data[34219] <= 8'h10 ;
			data[34220] <= 8'h10 ;
			data[34221] <= 8'h10 ;
			data[34222] <= 8'h10 ;
			data[34223] <= 8'h10 ;
			data[34224] <= 8'h10 ;
			data[34225] <= 8'h10 ;
			data[34226] <= 8'h10 ;
			data[34227] <= 8'h10 ;
			data[34228] <= 8'h10 ;
			data[34229] <= 8'h10 ;
			data[34230] <= 8'h10 ;
			data[34231] <= 8'h10 ;
			data[34232] <= 8'h10 ;
			data[34233] <= 8'h10 ;
			data[34234] <= 8'h10 ;
			data[34235] <= 8'h10 ;
			data[34236] <= 8'h10 ;
			data[34237] <= 8'h10 ;
			data[34238] <= 8'h10 ;
			data[34239] <= 8'h10 ;
			data[34240] <= 8'h10 ;
			data[34241] <= 8'h10 ;
			data[34242] <= 8'h10 ;
			data[34243] <= 8'h10 ;
			data[34244] <= 8'h10 ;
			data[34245] <= 8'h10 ;
			data[34246] <= 8'h10 ;
			data[34247] <= 8'h10 ;
			data[34248] <= 8'h10 ;
			data[34249] <= 8'h10 ;
			data[34250] <= 8'h10 ;
			data[34251] <= 8'h10 ;
			data[34252] <= 8'h10 ;
			data[34253] <= 8'h10 ;
			data[34254] <= 8'h10 ;
			data[34255] <= 8'h10 ;
			data[34256] <= 8'h10 ;
			data[34257] <= 8'h10 ;
			data[34258] <= 8'h10 ;
			data[34259] <= 8'h10 ;
			data[34260] <= 8'h10 ;
			data[34261] <= 8'h10 ;
			data[34262] <= 8'h10 ;
			data[34263] <= 8'h10 ;
			data[34264] <= 8'h10 ;
			data[34265] <= 8'h10 ;
			data[34266] <= 8'h10 ;
			data[34267] <= 8'h10 ;
			data[34268] <= 8'h10 ;
			data[34269] <= 8'h10 ;
			data[34270] <= 8'h10 ;
			data[34271] <= 8'h10 ;
			data[34272] <= 8'h10 ;
			data[34273] <= 8'h10 ;
			data[34274] <= 8'h10 ;
			data[34275] <= 8'h10 ;
			data[34276] <= 8'h10 ;
			data[34277] <= 8'h10 ;
			data[34278] <= 8'h10 ;
			data[34279] <= 8'h10 ;
			data[34280] <= 8'h10 ;
			data[34281] <= 8'h10 ;
			data[34282] <= 8'h10 ;
			data[34283] <= 8'h10 ;
			data[34284] <= 8'h10 ;
			data[34285] <= 8'h10 ;
			data[34286] <= 8'h10 ;
			data[34287] <= 8'h10 ;
			data[34288] <= 8'h10 ;
			data[34289] <= 8'h10 ;
			data[34290] <= 8'h10 ;
			data[34291] <= 8'h10 ;
			data[34292] <= 8'h10 ;
			data[34293] <= 8'h10 ;
			data[34294] <= 8'h10 ;
			data[34295] <= 8'h10 ;
			data[34296] <= 8'h10 ;
			data[34297] <= 8'h10 ;
			data[34298] <= 8'h10 ;
			data[34299] <= 8'h10 ;
			data[34300] <= 8'h10 ;
			data[34301] <= 8'h10 ;
			data[34302] <= 8'h10 ;
			data[34303] <= 8'h10 ;
			data[34304] <= 8'h10 ;
			data[34305] <= 8'h10 ;
			data[34306] <= 8'h10 ;
			data[34307] <= 8'h10 ;
			data[34308] <= 8'h10 ;
			data[34309] <= 8'h10 ;
			data[34310] <= 8'h10 ;
			data[34311] <= 8'h10 ;
			data[34312] <= 8'h10 ;
			data[34313] <= 8'h10 ;
			data[34314] <= 8'h10 ;
			data[34315] <= 8'h10 ;
			data[34316] <= 8'h10 ;
			data[34317] <= 8'h10 ;
			data[34318] <= 8'h10 ;
			data[34319] <= 8'h10 ;
			data[34320] <= 8'h10 ;
			data[34321] <= 8'h10 ;
			data[34322] <= 8'h10 ;
			data[34323] <= 8'h10 ;
			data[34324] <= 8'h10 ;
			data[34325] <= 8'h10 ;
			data[34326] <= 8'h10 ;
			data[34327] <= 8'h10 ;
			data[34328] <= 8'h10 ;
			data[34329] <= 8'h10 ;
			data[34330] <= 8'h10 ;
			data[34331] <= 8'h10 ;
			data[34332] <= 8'h10 ;
			data[34333] <= 8'h10 ;
			data[34334] <= 8'h10 ;
			data[34335] <= 8'h10 ;
			data[34336] <= 8'h10 ;
			data[34337] <= 8'h10 ;
			data[34338] <= 8'h10 ;
			data[34339] <= 8'h10 ;
			data[34340] <= 8'h10 ;
			data[34341] <= 8'h10 ;
			data[34342] <= 8'h10 ;
			data[34343] <= 8'h10 ;
			data[34344] <= 8'h10 ;
			data[34345] <= 8'h10 ;
			data[34346] <= 8'h10 ;
			data[34347] <= 8'h10 ;
			data[34348] <= 8'h10 ;
			data[34349] <= 8'h10 ;
			data[34350] <= 8'h10 ;
			data[34351] <= 8'h10 ;
			data[34352] <= 8'h10 ;
			data[34353] <= 8'h10 ;
			data[34354] <= 8'h10 ;
			data[34355] <= 8'h10 ;
			data[34356] <= 8'h10 ;
			data[34357] <= 8'h10 ;
			data[34358] <= 8'h10 ;
			data[34359] <= 8'h10 ;
			data[34360] <= 8'h10 ;
			data[34361] <= 8'h10 ;
			data[34362] <= 8'h10 ;
			data[34363] <= 8'h10 ;
			data[34364] <= 8'h10 ;
			data[34365] <= 8'h10 ;
			data[34366] <= 8'h10 ;
			data[34367] <= 8'h10 ;
			data[34368] <= 8'h10 ;
			data[34369] <= 8'h10 ;
			data[34370] <= 8'h10 ;
			data[34371] <= 8'h10 ;
			data[34372] <= 8'h10 ;
			data[34373] <= 8'h10 ;
			data[34374] <= 8'h10 ;
			data[34375] <= 8'h10 ;
			data[34376] <= 8'h10 ;
			data[34377] <= 8'h10 ;
			data[34378] <= 8'h10 ;
			data[34379] <= 8'h10 ;
			data[34380] <= 8'h10 ;
			data[34381] <= 8'h10 ;
			data[34382] <= 8'h10 ;
			data[34383] <= 8'h10 ;
			data[34384] <= 8'h10 ;
			data[34385] <= 8'h10 ;
			data[34386] <= 8'h10 ;
			data[34387] <= 8'h10 ;
			data[34388] <= 8'h10 ;
			data[34389] <= 8'h10 ;
			data[34390] <= 8'h10 ;
			data[34391] <= 8'h10 ;
			data[34392] <= 8'h10 ;
			data[34393] <= 8'h10 ;
			data[34394] <= 8'h10 ;
			data[34395] <= 8'h10 ;
			data[34396] <= 8'h10 ;
			data[34397] <= 8'h10 ;
			data[34398] <= 8'h10 ;
			data[34399] <= 8'h10 ;
			data[34400] <= 8'h10 ;
			data[34401] <= 8'h10 ;
			data[34402] <= 8'h10 ;
			data[34403] <= 8'h10 ;
			data[34404] <= 8'h10 ;
			data[34405] <= 8'h10 ;
			data[34406] <= 8'h10 ;
			data[34407] <= 8'h10 ;
			data[34408] <= 8'h10 ;
			data[34409] <= 8'h10 ;
			data[34410] <= 8'h10 ;
			data[34411] <= 8'h10 ;
			data[34412] <= 8'h10 ;
			data[34413] <= 8'h10 ;
			data[34414] <= 8'h10 ;
			data[34415] <= 8'h10 ;
			data[34416] <= 8'h10 ;
			data[34417] <= 8'h10 ;
			data[34418] <= 8'h10 ;
			data[34419] <= 8'h10 ;
			data[34420] <= 8'h10 ;
			data[34421] <= 8'h10 ;
			data[34422] <= 8'h10 ;
			data[34423] <= 8'h10 ;
			data[34424] <= 8'h10 ;
			data[34425] <= 8'h10 ;
			data[34426] <= 8'h10 ;
			data[34427] <= 8'h10 ;
			data[34428] <= 8'h10 ;
			data[34429] <= 8'h10 ;
			data[34430] <= 8'h10 ;
			data[34431] <= 8'h10 ;
			data[34432] <= 8'h10 ;
			data[34433] <= 8'h10 ;
			data[34434] <= 8'h10 ;
			data[34435] <= 8'h10 ;
			data[34436] <= 8'h10 ;
			data[34437] <= 8'h10 ;
			data[34438] <= 8'h10 ;
			data[34439] <= 8'h10 ;
			data[34440] <= 8'h10 ;
			data[34441] <= 8'h10 ;
			data[34442] <= 8'h10 ;
			data[34443] <= 8'h10 ;
			data[34444] <= 8'h10 ;
			data[34445] <= 8'h10 ;
			data[34446] <= 8'h10 ;
			data[34447] <= 8'h10 ;
			data[34448] <= 8'h10 ;
			data[34449] <= 8'h10 ;
			data[34450] <= 8'h10 ;
			data[34451] <= 8'h10 ;
			data[34452] <= 8'h10 ;
			data[34453] <= 8'h10 ;
			data[34454] <= 8'h10 ;
			data[34455] <= 8'h10 ;
			data[34456] <= 8'h10 ;
			data[34457] <= 8'h10 ;
			data[34458] <= 8'h10 ;
			data[34459] <= 8'h10 ;
			data[34460] <= 8'h10 ;
			data[34461] <= 8'h10 ;
			data[34462] <= 8'h10 ;
			data[34463] <= 8'h10 ;
			data[34464] <= 8'h10 ;
			data[34465] <= 8'h10 ;
			data[34466] <= 8'h10 ;
			data[34467] <= 8'h10 ;
			data[34468] <= 8'h10 ;
			data[34469] <= 8'h10 ;
			data[34470] <= 8'h10 ;
			data[34471] <= 8'h10 ;
			data[34472] <= 8'h10 ;
			data[34473] <= 8'h10 ;
			data[34474] <= 8'h10 ;
			data[34475] <= 8'h10 ;
			data[34476] <= 8'h10 ;
			data[34477] <= 8'h10 ;
			data[34478] <= 8'h10 ;
			data[34479] <= 8'h10 ;
			data[34480] <= 8'h10 ;
			data[34481] <= 8'h10 ;
			data[34482] <= 8'h10 ;
			data[34483] <= 8'h10 ;
			data[34484] <= 8'h10 ;
			data[34485] <= 8'h10 ;
			data[34486] <= 8'h10 ;
			data[34487] <= 8'h10 ;
			data[34488] <= 8'h10 ;
			data[34489] <= 8'h10 ;
			data[34490] <= 8'h10 ;
			data[34491] <= 8'h10 ;
			data[34492] <= 8'h10 ;
			data[34493] <= 8'h10 ;
			data[34494] <= 8'h10 ;
			data[34495] <= 8'h10 ;
			data[34496] <= 8'h10 ;
			data[34497] <= 8'h10 ;
			data[34498] <= 8'h10 ;
			data[34499] <= 8'h10 ;
			data[34500] <= 8'h10 ;
			data[34501] <= 8'h10 ;
			data[34502] <= 8'h10 ;
			data[34503] <= 8'h10 ;
			data[34504] <= 8'h10 ;
			data[34505] <= 8'h10 ;
			data[34506] <= 8'h10 ;
			data[34507] <= 8'h10 ;
			data[34508] <= 8'h10 ;
			data[34509] <= 8'h10 ;
			data[34510] <= 8'h10 ;
			data[34511] <= 8'h10 ;
			data[34512] <= 8'h10 ;
			data[34513] <= 8'h10 ;
			data[34514] <= 8'h10 ;
			data[34515] <= 8'h10 ;
			data[34516] <= 8'h10 ;
			data[34517] <= 8'h10 ;
			data[34518] <= 8'h10 ;
			data[34519] <= 8'h10 ;
			data[34520] <= 8'h10 ;
			data[34521] <= 8'h10 ;
			data[34522] <= 8'h10 ;
			data[34523] <= 8'h10 ;
			data[34524] <= 8'h10 ;
			data[34525] <= 8'h10 ;
			data[34526] <= 8'h10 ;
			data[34527] <= 8'h10 ;
			data[34528] <= 8'h10 ;
			data[34529] <= 8'h10 ;
			data[34530] <= 8'h10 ;
			data[34531] <= 8'h10 ;
			data[34532] <= 8'h10 ;
			data[34533] <= 8'h10 ;
			data[34534] <= 8'h10 ;
			data[34535] <= 8'h10 ;
			data[34536] <= 8'h10 ;
			data[34537] <= 8'h10 ;
			data[34538] <= 8'h10 ;
			data[34539] <= 8'h10 ;
			data[34540] <= 8'h10 ;
			data[34541] <= 8'h10 ;
			data[34542] <= 8'h10 ;
			data[34543] <= 8'h10 ;
			data[34544] <= 8'h10 ;
			data[34545] <= 8'h10 ;
			data[34546] <= 8'h10 ;
			data[34547] <= 8'h10 ;
			data[34548] <= 8'h10 ;
			data[34549] <= 8'h10 ;
			data[34550] <= 8'h10 ;
			data[34551] <= 8'h10 ;
			data[34552] <= 8'h10 ;
			data[34553] <= 8'h10 ;
			data[34554] <= 8'h10 ;
			data[34555] <= 8'h10 ;
			data[34556] <= 8'h10 ;
			data[34557] <= 8'h10 ;
			data[34558] <= 8'h10 ;
			data[34559] <= 8'h10 ;
			data[34560] <= 8'h10 ;
			data[34561] <= 8'h10 ;
			data[34562] <= 8'h10 ;
			data[34563] <= 8'h10 ;
			data[34564] <= 8'h10 ;
			data[34565] <= 8'h10 ;
			data[34566] <= 8'h10 ;
			data[34567] <= 8'h10 ;
			data[34568] <= 8'h10 ;
			data[34569] <= 8'h10 ;
			data[34570] <= 8'h10 ;
			data[34571] <= 8'h10 ;
			data[34572] <= 8'h10 ;
			data[34573] <= 8'h10 ;
			data[34574] <= 8'h10 ;
			data[34575] <= 8'h10 ;
			data[34576] <= 8'h10 ;
			data[34577] <= 8'h10 ;
			data[34578] <= 8'h10 ;
			data[34579] <= 8'h10 ;
			data[34580] <= 8'h10 ;
			data[34581] <= 8'h10 ;
			data[34582] <= 8'h10 ;
			data[34583] <= 8'h10 ;
			data[34584] <= 8'h10 ;
			data[34585] <= 8'h10 ;
			data[34586] <= 8'h10 ;
			data[34587] <= 8'h10 ;
			data[34588] <= 8'h10 ;
			data[34589] <= 8'h10 ;
			data[34590] <= 8'h10 ;
			data[34591] <= 8'h10 ;
			data[34592] <= 8'h10 ;
			data[34593] <= 8'h10 ;
			data[34594] <= 8'h10 ;
			data[34595] <= 8'h10 ;
			data[34596] <= 8'h10 ;
			data[34597] <= 8'h10 ;
			data[34598] <= 8'h10 ;
			data[34599] <= 8'h10 ;
			data[34600] <= 8'h10 ;
			data[34601] <= 8'h10 ;
			data[34602] <= 8'h10 ;
			data[34603] <= 8'h10 ;
			data[34604] <= 8'h10 ;
			data[34605] <= 8'h10 ;
			data[34606] <= 8'h10 ;
			data[34607] <= 8'h10 ;
			data[34608] <= 8'h10 ;
			data[34609] <= 8'h10 ;
			data[34610] <= 8'h10 ;
			data[34611] <= 8'h10 ;
			data[34612] <= 8'h10 ;
			data[34613] <= 8'h10 ;
			data[34614] <= 8'h10 ;
			data[34615] <= 8'h10 ;
			data[34616] <= 8'h10 ;
			data[34617] <= 8'h10 ;
			data[34618] <= 8'h10 ;
			data[34619] <= 8'h10 ;
			data[34620] <= 8'h10 ;
			data[34621] <= 8'h10 ;
			data[34622] <= 8'h10 ;
			data[34623] <= 8'h10 ;
			data[34624] <= 8'h10 ;
			data[34625] <= 8'h10 ;
			data[34626] <= 8'h10 ;
			data[34627] <= 8'h10 ;
			data[34628] <= 8'h10 ;
			data[34629] <= 8'h10 ;
			data[34630] <= 8'h10 ;
			data[34631] <= 8'h10 ;
			data[34632] <= 8'h10 ;
			data[34633] <= 8'h10 ;
			data[34634] <= 8'h10 ;
			data[34635] <= 8'h10 ;
			data[34636] <= 8'h10 ;
			data[34637] <= 8'h10 ;
			data[34638] <= 8'h10 ;
			data[34639] <= 8'h10 ;
			data[34640] <= 8'h10 ;
			data[34641] <= 8'h10 ;
			data[34642] <= 8'h10 ;
			data[34643] <= 8'h10 ;
			data[34644] <= 8'h10 ;
			data[34645] <= 8'h10 ;
			data[34646] <= 8'h10 ;
			data[34647] <= 8'h10 ;
			data[34648] <= 8'h10 ;
			data[34649] <= 8'h10 ;
			data[34650] <= 8'h10 ;
			data[34651] <= 8'h10 ;
			data[34652] <= 8'h10 ;
			data[34653] <= 8'h10 ;
			data[34654] <= 8'h10 ;
			data[34655] <= 8'h10 ;
			data[34656] <= 8'h10 ;
			data[34657] <= 8'h10 ;
			data[34658] <= 8'h10 ;
			data[34659] <= 8'h10 ;
			data[34660] <= 8'h10 ;
			data[34661] <= 8'h10 ;
			data[34662] <= 8'h10 ;
			data[34663] <= 8'h10 ;
			data[34664] <= 8'h10 ;
			data[34665] <= 8'h10 ;
			data[34666] <= 8'h10 ;
			data[34667] <= 8'h10 ;
			data[34668] <= 8'h10 ;
			data[34669] <= 8'h10 ;
			data[34670] <= 8'h10 ;
			data[34671] <= 8'h10 ;
			data[34672] <= 8'h10 ;
			data[34673] <= 8'h10 ;
			data[34674] <= 8'h10 ;
			data[34675] <= 8'h10 ;
			data[34676] <= 8'h10 ;
			data[34677] <= 8'h10 ;
			data[34678] <= 8'h10 ;
			data[34679] <= 8'h10 ;
			data[34680] <= 8'h10 ;
			data[34681] <= 8'h10 ;
			data[34682] <= 8'h10 ;
			data[34683] <= 8'h10 ;
			data[34684] <= 8'h10 ;
			data[34685] <= 8'h10 ;
			data[34686] <= 8'h10 ;
			data[34687] <= 8'h10 ;
			data[34688] <= 8'h10 ;
			data[34689] <= 8'h10 ;
			data[34690] <= 8'h10 ;
			data[34691] <= 8'h10 ;
			data[34692] <= 8'h10 ;
			data[34693] <= 8'h10 ;
			data[34694] <= 8'h10 ;
			data[34695] <= 8'h10 ;
			data[34696] <= 8'h10 ;
			data[34697] <= 8'h10 ;
			data[34698] <= 8'h10 ;
			data[34699] <= 8'h10 ;
			data[34700] <= 8'h10 ;
			data[34701] <= 8'h10 ;
			data[34702] <= 8'h10 ;
			data[34703] <= 8'h10 ;
			data[34704] <= 8'h10 ;
			data[34705] <= 8'h10 ;
			data[34706] <= 8'h10 ;
			data[34707] <= 8'h10 ;
			data[34708] <= 8'h10 ;
			data[34709] <= 8'h10 ;
			data[34710] <= 8'h10 ;
			data[34711] <= 8'h10 ;
			data[34712] <= 8'h10 ;
			data[34713] <= 8'h10 ;
			data[34714] <= 8'h10 ;
			data[34715] <= 8'h10 ;
			data[34716] <= 8'h10 ;
			data[34717] <= 8'h10 ;
			data[34718] <= 8'h10 ;
			data[34719] <= 8'h10 ;
			data[34720] <= 8'h10 ;
			data[34721] <= 8'h10 ;
			data[34722] <= 8'h10 ;
			data[34723] <= 8'h10 ;
			data[34724] <= 8'h10 ;
			data[34725] <= 8'h10 ;
			data[34726] <= 8'h10 ;
			data[34727] <= 8'h10 ;
			data[34728] <= 8'h10 ;
			data[34729] <= 8'h10 ;
			data[34730] <= 8'h10 ;
			data[34731] <= 8'h10 ;
			data[34732] <= 8'h10 ;
			data[34733] <= 8'h10 ;
			data[34734] <= 8'h10 ;
			data[34735] <= 8'h10 ;
			data[34736] <= 8'h10 ;
			data[34737] <= 8'h10 ;
			data[34738] <= 8'h10 ;
			data[34739] <= 8'h10 ;
			data[34740] <= 8'h10 ;
			data[34741] <= 8'h10 ;
			data[34742] <= 8'h10 ;
			data[34743] <= 8'h10 ;
			data[34744] <= 8'h10 ;
			data[34745] <= 8'h10 ;
			data[34746] <= 8'h10 ;
			data[34747] <= 8'h10 ;
			data[34748] <= 8'h10 ;
			data[34749] <= 8'h10 ;
			data[34750] <= 8'h10 ;
			data[34751] <= 8'h10 ;
			data[34752] <= 8'h10 ;
			data[34753] <= 8'h10 ;
			data[34754] <= 8'h10 ;
			data[34755] <= 8'h10 ;
			data[34756] <= 8'h10 ;
			data[34757] <= 8'h10 ;
			data[34758] <= 8'h10 ;
			data[34759] <= 8'h10 ;
			data[34760] <= 8'h10 ;
			data[34761] <= 8'h10 ;
			data[34762] <= 8'h10 ;
			data[34763] <= 8'h10 ;
			data[34764] <= 8'h10 ;
			data[34765] <= 8'h10 ;
			data[34766] <= 8'h10 ;
			data[34767] <= 8'h10 ;
			data[34768] <= 8'h10 ;
			data[34769] <= 8'h10 ;
			data[34770] <= 8'h10 ;
			data[34771] <= 8'h10 ;
			data[34772] <= 8'h10 ;
			data[34773] <= 8'h10 ;
			data[34774] <= 8'h10 ;
			data[34775] <= 8'h10 ;
			data[34776] <= 8'h10 ;
			data[34777] <= 8'h10 ;
			data[34778] <= 8'h10 ;
			data[34779] <= 8'h10 ;
			data[34780] <= 8'h10 ;
			data[34781] <= 8'h10 ;
			data[34782] <= 8'h10 ;
			data[34783] <= 8'h10 ;
			data[34784] <= 8'h10 ;
			data[34785] <= 8'h10 ;
			data[34786] <= 8'h10 ;
			data[34787] <= 8'h10 ;
			data[34788] <= 8'h10 ;
			data[34789] <= 8'h10 ;
			data[34790] <= 8'h10 ;
			data[34791] <= 8'h10 ;
			data[34792] <= 8'h10 ;
			data[34793] <= 8'h10 ;
			data[34794] <= 8'h10 ;
			data[34795] <= 8'h10 ;
			data[34796] <= 8'h10 ;
			data[34797] <= 8'h10 ;
			data[34798] <= 8'h10 ;
			data[34799] <= 8'h10 ;
			data[34800] <= 8'h10 ;
			data[34801] <= 8'h10 ;
			data[34802] <= 8'h10 ;
			data[34803] <= 8'h10 ;
			data[34804] <= 8'h10 ;
			data[34805] <= 8'h10 ;
			data[34806] <= 8'h10 ;
			data[34807] <= 8'h10 ;
			data[34808] <= 8'h10 ;
			data[34809] <= 8'h10 ;
			data[34810] <= 8'h10 ;
			data[34811] <= 8'h10 ;
			data[34812] <= 8'h10 ;
			data[34813] <= 8'h10 ;
			data[34814] <= 8'h10 ;
			data[34815] <= 8'h10 ;
			data[34816] <= 8'h10 ;
			data[34817] <= 8'h10 ;
			data[34818] <= 8'h10 ;
			data[34819] <= 8'h10 ;
			data[34820] <= 8'h10 ;
			data[34821] <= 8'h10 ;
			data[34822] <= 8'h10 ;
			data[34823] <= 8'h10 ;
			data[34824] <= 8'h10 ;
			data[34825] <= 8'h10 ;
			data[34826] <= 8'h10 ;
			data[34827] <= 8'h10 ;
			data[34828] <= 8'h10 ;
			data[34829] <= 8'h10 ;
			data[34830] <= 8'h10 ;
			data[34831] <= 8'h10 ;
			data[34832] <= 8'h10 ;
			data[34833] <= 8'h10 ;
			data[34834] <= 8'h10 ;
			data[34835] <= 8'h10 ;
			data[34836] <= 8'h10 ;
			data[34837] <= 8'h10 ;
			data[34838] <= 8'h10 ;
			data[34839] <= 8'h10 ;
			data[34840] <= 8'h10 ;
			data[34841] <= 8'h10 ;
			data[34842] <= 8'h10 ;
			data[34843] <= 8'h10 ;
			data[34844] <= 8'h10 ;
			data[34845] <= 8'h10 ;
			data[34846] <= 8'h10 ;
			data[34847] <= 8'h10 ;
			data[34848] <= 8'h10 ;
			data[34849] <= 8'h10 ;
			data[34850] <= 8'h10 ;
			data[34851] <= 8'h10 ;
			data[34852] <= 8'h10 ;
			data[34853] <= 8'h10 ;
			data[34854] <= 8'h10 ;
			data[34855] <= 8'h10 ;
			data[34856] <= 8'h10 ;
			data[34857] <= 8'h10 ;
			data[34858] <= 8'h10 ;
			data[34859] <= 8'h10 ;
			data[34860] <= 8'h10 ;
			data[34861] <= 8'h10 ;
			data[34862] <= 8'h10 ;
			data[34863] <= 8'h10 ;
			data[34864] <= 8'h10 ;
			data[34865] <= 8'h10 ;
			data[34866] <= 8'h10 ;
			data[34867] <= 8'h10 ;
			data[34868] <= 8'h10 ;
			data[34869] <= 8'h10 ;
			data[34870] <= 8'h10 ;
			data[34871] <= 8'h10 ;
			data[34872] <= 8'h10 ;
			data[34873] <= 8'h10 ;
			data[34874] <= 8'h10 ;
			data[34875] <= 8'h10 ;
			data[34876] <= 8'h10 ;
			data[34877] <= 8'h10 ;
			data[34878] <= 8'h10 ;
			data[34879] <= 8'h10 ;
			data[34880] <= 8'h10 ;
			data[34881] <= 8'h10 ;
			data[34882] <= 8'h10 ;
			data[34883] <= 8'h10 ;
			data[34884] <= 8'h10 ;
			data[34885] <= 8'h10 ;
			data[34886] <= 8'h10 ;
			data[34887] <= 8'h10 ;
			data[34888] <= 8'h10 ;
			data[34889] <= 8'h10 ;
			data[34890] <= 8'h10 ;
			data[34891] <= 8'h10 ;
			data[34892] <= 8'h10 ;
			data[34893] <= 8'h10 ;
			data[34894] <= 8'h10 ;
			data[34895] <= 8'h10 ;
			data[34896] <= 8'h10 ;
			data[34897] <= 8'h10 ;
			data[34898] <= 8'h10 ;
			data[34899] <= 8'h10 ;
			data[34900] <= 8'h10 ;
			data[34901] <= 8'h10 ;
			data[34902] <= 8'h10 ;
			data[34903] <= 8'h10 ;
			data[34904] <= 8'h10 ;
			data[34905] <= 8'h10 ;
			data[34906] <= 8'h10 ;
			data[34907] <= 8'h10 ;
			data[34908] <= 8'h10 ;
			data[34909] <= 8'h10 ;
			data[34910] <= 8'h10 ;
			data[34911] <= 8'h10 ;
			data[34912] <= 8'h10 ;
			data[34913] <= 8'h10 ;
			data[34914] <= 8'h10 ;
			data[34915] <= 8'h10 ;
			data[34916] <= 8'h10 ;
			data[34917] <= 8'h10 ;
			data[34918] <= 8'h10 ;
			data[34919] <= 8'h10 ;
			data[34920] <= 8'h10 ;
			data[34921] <= 8'h10 ;
			data[34922] <= 8'h10 ;
			data[34923] <= 8'h10 ;
			data[34924] <= 8'h10 ;
			data[34925] <= 8'h10 ;
			data[34926] <= 8'h10 ;
			data[34927] <= 8'h10 ;
			data[34928] <= 8'h10 ;
			data[34929] <= 8'h10 ;
			data[34930] <= 8'h10 ;
			data[34931] <= 8'h10 ;
			data[34932] <= 8'h10 ;
			data[34933] <= 8'h10 ;
			data[34934] <= 8'h10 ;
			data[34935] <= 8'h10 ;
			data[34936] <= 8'h10 ;
			data[34937] <= 8'h10 ;
			data[34938] <= 8'h10 ;
			data[34939] <= 8'h10 ;
			data[34940] <= 8'h10 ;
			data[34941] <= 8'h10 ;
			data[34942] <= 8'h10 ;
			data[34943] <= 8'h10 ;
			data[34944] <= 8'h10 ;
			data[34945] <= 8'h10 ;
			data[34946] <= 8'h10 ;
			data[34947] <= 8'h10 ;
			data[34948] <= 8'h10 ;
			data[34949] <= 8'h10 ;
			data[34950] <= 8'h10 ;
			data[34951] <= 8'h10 ;
			data[34952] <= 8'h10 ;
			data[34953] <= 8'h10 ;
			data[34954] <= 8'h10 ;
			data[34955] <= 8'h10 ;
			data[34956] <= 8'h10 ;
			data[34957] <= 8'h10 ;
			data[34958] <= 8'h10 ;
			data[34959] <= 8'h10 ;
			data[34960] <= 8'h10 ;
			data[34961] <= 8'h10 ;
			data[34962] <= 8'h10 ;
			data[34963] <= 8'h10 ;
			data[34964] <= 8'h10 ;
			data[34965] <= 8'h10 ;
			data[34966] <= 8'h10 ;
			data[34967] <= 8'h10 ;
			data[34968] <= 8'h10 ;
			data[34969] <= 8'h10 ;
			data[34970] <= 8'h10 ;
			data[34971] <= 8'h10 ;
			data[34972] <= 8'h10 ;
			data[34973] <= 8'h10 ;
			data[34974] <= 8'h10 ;
			data[34975] <= 8'h10 ;
			data[34976] <= 8'h10 ;
			data[34977] <= 8'h10 ;
			data[34978] <= 8'h10 ;
			data[34979] <= 8'h10 ;
			data[34980] <= 8'h10 ;
			data[34981] <= 8'h10 ;
			data[34982] <= 8'h10 ;
			data[34983] <= 8'h10 ;
			data[34984] <= 8'h10 ;
			data[34985] <= 8'h10 ;
			data[34986] <= 8'h10 ;
			data[34987] <= 8'h10 ;
			data[34988] <= 8'h10 ;
			data[34989] <= 8'h10 ;
			data[34990] <= 8'h10 ;
			data[34991] <= 8'h10 ;
			data[34992] <= 8'h10 ;
			data[34993] <= 8'h10 ;
			data[34994] <= 8'h10 ;
			data[34995] <= 8'h10 ;
			data[34996] <= 8'h10 ;
			data[34997] <= 8'h10 ;
			data[34998] <= 8'h10 ;
			data[34999] <= 8'h10 ;
			data[35000] <= 8'h10 ;
			data[35001] <= 8'h10 ;
			data[35002] <= 8'h10 ;
			data[35003] <= 8'h10 ;
			data[35004] <= 8'h10 ;
			data[35005] <= 8'h10 ;
			data[35006] <= 8'h10 ;
			data[35007] <= 8'h10 ;
			data[35008] <= 8'h10 ;
			data[35009] <= 8'h10 ;
			data[35010] <= 8'h10 ;
			data[35011] <= 8'h10 ;
			data[35012] <= 8'h10 ;
			data[35013] <= 8'h10 ;
			data[35014] <= 8'h10 ;
			data[35015] <= 8'h10 ;
			data[35016] <= 8'h10 ;
			data[35017] <= 8'h10 ;
			data[35018] <= 8'h10 ;
			data[35019] <= 8'h10 ;
			data[35020] <= 8'h10 ;
			data[35021] <= 8'h10 ;
			data[35022] <= 8'h10 ;
			data[35023] <= 8'h10 ;
			data[35024] <= 8'h10 ;
			data[35025] <= 8'h10 ;
			data[35026] <= 8'h10 ;
			data[35027] <= 8'h10 ;
			data[35028] <= 8'h10 ;
			data[35029] <= 8'h10 ;
			data[35030] <= 8'h10 ;
			data[35031] <= 8'h10 ;
			data[35032] <= 8'h10 ;
			data[35033] <= 8'h10 ;
			data[35034] <= 8'h10 ;
			data[35035] <= 8'h10 ;
			data[35036] <= 8'h10 ;
			data[35037] <= 8'h10 ;
			data[35038] <= 8'h10 ;
			data[35039] <= 8'h10 ;
			data[35040] <= 8'h10 ;
			data[35041] <= 8'h10 ;
			data[35042] <= 8'h10 ;
			data[35043] <= 8'h10 ;
			data[35044] <= 8'h10 ;
			data[35045] <= 8'h10 ;
			data[35046] <= 8'h10 ;
			data[35047] <= 8'h10 ;
			data[35048] <= 8'h10 ;
			data[35049] <= 8'h10 ;
			data[35050] <= 8'h10 ;
			data[35051] <= 8'h10 ;
			data[35052] <= 8'h10 ;
			data[35053] <= 8'h10 ;
			data[35054] <= 8'h10 ;
			data[35055] <= 8'h10 ;
			data[35056] <= 8'h10 ;
			data[35057] <= 8'h10 ;
			data[35058] <= 8'h10 ;
			data[35059] <= 8'h10 ;
			data[35060] <= 8'h10 ;
			data[35061] <= 8'h10 ;
			data[35062] <= 8'h10 ;
			data[35063] <= 8'h10 ;
			data[35064] <= 8'h10 ;
			data[35065] <= 8'h10 ;
			data[35066] <= 8'h10 ;
			data[35067] <= 8'h10 ;
			data[35068] <= 8'h10 ;
			data[35069] <= 8'h10 ;
			data[35070] <= 8'h10 ;
			data[35071] <= 8'h10 ;
			data[35072] <= 8'h10 ;
			data[35073] <= 8'h10 ;
			data[35074] <= 8'h10 ;
			data[35075] <= 8'h10 ;
			data[35076] <= 8'h10 ;
			data[35077] <= 8'h10 ;
			data[35078] <= 8'h10 ;
			data[35079] <= 8'h10 ;
			data[35080] <= 8'h10 ;
			data[35081] <= 8'h10 ;
			data[35082] <= 8'h10 ;
			data[35083] <= 8'h10 ;
			data[35084] <= 8'h10 ;
			data[35085] <= 8'h10 ;
			data[35086] <= 8'h10 ;
			data[35087] <= 8'h10 ;
			data[35088] <= 8'h10 ;
			data[35089] <= 8'h10 ;
			data[35090] <= 8'h10 ;
			data[35091] <= 8'h10 ;
			data[35092] <= 8'h10 ;
			data[35093] <= 8'h10 ;
			data[35094] <= 8'h10 ;
			data[35095] <= 8'h10 ;
			data[35096] <= 8'h10 ;
			data[35097] <= 8'h10 ;
			data[35098] <= 8'h10 ;
			data[35099] <= 8'h10 ;
			data[35100] <= 8'h10 ;
			data[35101] <= 8'h10 ;
			data[35102] <= 8'h10 ;
			data[35103] <= 8'h10 ;
			data[35104] <= 8'h10 ;
			data[35105] <= 8'h10 ;
			data[35106] <= 8'h10 ;
			data[35107] <= 8'h10 ;
			data[35108] <= 8'h10 ;
			data[35109] <= 8'h10 ;
			data[35110] <= 8'h10 ;
			data[35111] <= 8'h10 ;
			data[35112] <= 8'h10 ;
			data[35113] <= 8'h10 ;
			data[35114] <= 8'h10 ;
			data[35115] <= 8'h10 ;
			data[35116] <= 8'h10 ;
			data[35117] <= 8'h10 ;
			data[35118] <= 8'h10 ;
			data[35119] <= 8'h10 ;
			data[35120] <= 8'h10 ;
			data[35121] <= 8'h10 ;
			data[35122] <= 8'h10 ;
			data[35123] <= 8'h10 ;
			data[35124] <= 8'h10 ;
			data[35125] <= 8'h10 ;
			data[35126] <= 8'h10 ;
			data[35127] <= 8'h10 ;
			data[35128] <= 8'h10 ;
			data[35129] <= 8'h10 ;
			data[35130] <= 8'h10 ;
			data[35131] <= 8'h10 ;
			data[35132] <= 8'h10 ;
			data[35133] <= 8'h10 ;
			data[35134] <= 8'h10 ;
			data[35135] <= 8'h10 ;
			data[35136] <= 8'h10 ;
			data[35137] <= 8'h10 ;
			data[35138] <= 8'h10 ;
			data[35139] <= 8'h10 ;
			data[35140] <= 8'h10 ;
			data[35141] <= 8'h10 ;
			data[35142] <= 8'h10 ;
			data[35143] <= 8'h10 ;
			data[35144] <= 8'h10 ;
			data[35145] <= 8'h10 ;
			data[35146] <= 8'h10 ;
			data[35147] <= 8'h10 ;
			data[35148] <= 8'h10 ;
			data[35149] <= 8'h10 ;
			data[35150] <= 8'h10 ;
			data[35151] <= 8'h10 ;
			data[35152] <= 8'h10 ;
			data[35153] <= 8'h10 ;
			data[35154] <= 8'h10 ;
			data[35155] <= 8'h10 ;
			data[35156] <= 8'h10 ;
			data[35157] <= 8'h10 ;
			data[35158] <= 8'h10 ;
			data[35159] <= 8'h10 ;
			data[35160] <= 8'h10 ;
			data[35161] <= 8'h10 ;
			data[35162] <= 8'h10 ;
			data[35163] <= 8'h10 ;
			data[35164] <= 8'h10 ;
			data[35165] <= 8'h10 ;
			data[35166] <= 8'h10 ;
			data[35167] <= 8'h10 ;
			data[35168] <= 8'h10 ;
			data[35169] <= 8'h10 ;
			data[35170] <= 8'h10 ;
			data[35171] <= 8'h10 ;
			data[35172] <= 8'h10 ;
			data[35173] <= 8'h10 ;
			data[35174] <= 8'h10 ;
			data[35175] <= 8'h10 ;
			data[35176] <= 8'h10 ;
			data[35177] <= 8'h10 ;
			data[35178] <= 8'h10 ;
			data[35179] <= 8'h10 ;
			data[35180] <= 8'h10 ;
			data[35181] <= 8'h10 ;
			data[35182] <= 8'h10 ;
			data[35183] <= 8'h10 ;
			data[35184] <= 8'h10 ;
			data[35185] <= 8'h10 ;
			data[35186] <= 8'h10 ;
			data[35187] <= 8'h10 ;
			data[35188] <= 8'h10 ;
			data[35189] <= 8'h10 ;
			data[35190] <= 8'h10 ;
			data[35191] <= 8'h10 ;
			data[35192] <= 8'h10 ;
			data[35193] <= 8'h10 ;
			data[35194] <= 8'h10 ;
			data[35195] <= 8'h10 ;
			data[35196] <= 8'h10 ;
			data[35197] <= 8'h10 ;
			data[35198] <= 8'h10 ;
			data[35199] <= 8'h10 ;
			data[35200] <= 8'h10 ;
			data[35201] <= 8'h10 ;
			data[35202] <= 8'h10 ;
			data[35203] <= 8'h10 ;
			data[35204] <= 8'h10 ;
			data[35205] <= 8'h10 ;
			data[35206] <= 8'h10 ;
			data[35207] <= 8'h10 ;
			data[35208] <= 8'h10 ;
			data[35209] <= 8'h10 ;
			data[35210] <= 8'h10 ;
			data[35211] <= 8'h10 ;
			data[35212] <= 8'h10 ;
			data[35213] <= 8'h10 ;
			data[35214] <= 8'h10 ;
			data[35215] <= 8'h10 ;
			data[35216] <= 8'h10 ;
			data[35217] <= 8'h10 ;
			data[35218] <= 8'h10 ;
			data[35219] <= 8'h10 ;
			data[35220] <= 8'h10 ;
			data[35221] <= 8'h10 ;
			data[35222] <= 8'h10 ;
			data[35223] <= 8'h10 ;
			data[35224] <= 8'h10 ;
			data[35225] <= 8'h10 ;
			data[35226] <= 8'h10 ;
			data[35227] <= 8'h10 ;
			data[35228] <= 8'h10 ;
			data[35229] <= 8'h10 ;
			data[35230] <= 8'h10 ;
			data[35231] <= 8'h10 ;
			data[35232] <= 8'h10 ;
			data[35233] <= 8'h10 ;
			data[35234] <= 8'h10 ;
			data[35235] <= 8'h10 ;
			data[35236] <= 8'h10 ;
			data[35237] <= 8'h10 ;
			data[35238] <= 8'h10 ;
			data[35239] <= 8'h10 ;
			data[35240] <= 8'h10 ;
			data[35241] <= 8'h10 ;
			data[35242] <= 8'h10 ;
			data[35243] <= 8'h10 ;
			data[35244] <= 8'h10 ;
			data[35245] <= 8'h10 ;
			data[35246] <= 8'h10 ;
			data[35247] <= 8'h10 ;
			data[35248] <= 8'h10 ;
			data[35249] <= 8'h10 ;
			data[35250] <= 8'h10 ;
			data[35251] <= 8'h10 ;
			data[35252] <= 8'h10 ;
			data[35253] <= 8'h10 ;
			data[35254] <= 8'h10 ;
			data[35255] <= 8'h10 ;
			data[35256] <= 8'h10 ;
			data[35257] <= 8'h10 ;
			data[35258] <= 8'h10 ;
			data[35259] <= 8'h10 ;
			data[35260] <= 8'h10 ;
			data[35261] <= 8'h10 ;
			data[35262] <= 8'h10 ;
			data[35263] <= 8'h10 ;
			data[35264] <= 8'h10 ;
			data[35265] <= 8'h10 ;
			data[35266] <= 8'h10 ;
			data[35267] <= 8'h10 ;
			data[35268] <= 8'h10 ;
			data[35269] <= 8'h10 ;
			data[35270] <= 8'h10 ;
			data[35271] <= 8'h10 ;
			data[35272] <= 8'h10 ;
			data[35273] <= 8'h10 ;
			data[35274] <= 8'h10 ;
			data[35275] <= 8'h10 ;
			data[35276] <= 8'h10 ;
			data[35277] <= 8'h10 ;
			data[35278] <= 8'h10 ;
			data[35279] <= 8'h10 ;
			data[35280] <= 8'h10 ;
			data[35281] <= 8'h10 ;
			data[35282] <= 8'h10 ;
			data[35283] <= 8'h10 ;
			data[35284] <= 8'h10 ;
			data[35285] <= 8'h10 ;
			data[35286] <= 8'h10 ;
			data[35287] <= 8'h10 ;
			data[35288] <= 8'h10 ;
			data[35289] <= 8'h10 ;
			data[35290] <= 8'h10 ;
			data[35291] <= 8'h10 ;
			data[35292] <= 8'h10 ;
			data[35293] <= 8'h10 ;
			data[35294] <= 8'h10 ;
			data[35295] <= 8'h10 ;
			data[35296] <= 8'h10 ;
			data[35297] <= 8'h10 ;
			data[35298] <= 8'h10 ;
			data[35299] <= 8'h10 ;
			data[35300] <= 8'h10 ;
			data[35301] <= 8'h10 ;
			data[35302] <= 8'h10 ;
			data[35303] <= 8'h10 ;
			data[35304] <= 8'h10 ;
			data[35305] <= 8'h10 ;
			data[35306] <= 8'h10 ;
			data[35307] <= 8'h10 ;
			data[35308] <= 8'h10 ;
			data[35309] <= 8'h10 ;
			data[35310] <= 8'h10 ;
			data[35311] <= 8'h10 ;
			data[35312] <= 8'h10 ;
			data[35313] <= 8'h10 ;
			data[35314] <= 8'h10 ;
			data[35315] <= 8'h10 ;
			data[35316] <= 8'h10 ;
			data[35317] <= 8'h10 ;
			data[35318] <= 8'h10 ;
			data[35319] <= 8'h10 ;
			data[35320] <= 8'h10 ;
			data[35321] <= 8'h10 ;
			data[35322] <= 8'h10 ;
			data[35323] <= 8'h10 ;
			data[35324] <= 8'h10 ;
			data[35325] <= 8'h10 ;
			data[35326] <= 8'h10 ;
			data[35327] <= 8'h10 ;
			data[35328] <= 8'h10 ;
			data[35329] <= 8'h10 ;
			data[35330] <= 8'h10 ;
			data[35331] <= 8'h10 ;
			data[35332] <= 8'h10 ;
			data[35333] <= 8'h10 ;
			data[35334] <= 8'h10 ;
			data[35335] <= 8'h10 ;
			data[35336] <= 8'h10 ;
			data[35337] <= 8'h10 ;
			data[35338] <= 8'h10 ;
			data[35339] <= 8'h10 ;
			data[35340] <= 8'h10 ;
			data[35341] <= 8'h10 ;
			data[35342] <= 8'h10 ;
			data[35343] <= 8'h10 ;
			data[35344] <= 8'h10 ;
			data[35345] <= 8'h10 ;
			data[35346] <= 8'h10 ;
			data[35347] <= 8'h10 ;
			data[35348] <= 8'h10 ;
			data[35349] <= 8'h10 ;
			data[35350] <= 8'h10 ;
			data[35351] <= 8'h10 ;
			data[35352] <= 8'h10 ;
			data[35353] <= 8'h10 ;
			data[35354] <= 8'h10 ;
			data[35355] <= 8'h10 ;
			data[35356] <= 8'h10 ;
			data[35357] <= 8'h10 ;
			data[35358] <= 8'h10 ;
			data[35359] <= 8'h10 ;
			data[35360] <= 8'h10 ;
			data[35361] <= 8'h10 ;
			data[35362] <= 8'h10 ;
			data[35363] <= 8'h10 ;
			data[35364] <= 8'h10 ;
			data[35365] <= 8'h10 ;
			data[35366] <= 8'h10 ;
			data[35367] <= 8'h10 ;
			data[35368] <= 8'h10 ;
			data[35369] <= 8'h10 ;
			data[35370] <= 8'h10 ;
			data[35371] <= 8'h10 ;
			data[35372] <= 8'h10 ;
			data[35373] <= 8'h10 ;
			data[35374] <= 8'h10 ;
			data[35375] <= 8'h10 ;
			data[35376] <= 8'h10 ;
			data[35377] <= 8'h10 ;
			data[35378] <= 8'h10 ;
			data[35379] <= 8'h10 ;
			data[35380] <= 8'h10 ;
			data[35381] <= 8'h10 ;
			data[35382] <= 8'h10 ;
			data[35383] <= 8'h10 ;
			data[35384] <= 8'h10 ;
			data[35385] <= 8'h10 ;
			data[35386] <= 8'h10 ;
			data[35387] <= 8'h10 ;
			data[35388] <= 8'h10 ;
			data[35389] <= 8'h10 ;
			data[35390] <= 8'h10 ;
			data[35391] <= 8'h10 ;
			data[35392] <= 8'h10 ;
			data[35393] <= 8'h10 ;
			data[35394] <= 8'h10 ;
			data[35395] <= 8'h10 ;
			data[35396] <= 8'h10 ;
			data[35397] <= 8'h10 ;
			data[35398] <= 8'h10 ;
			data[35399] <= 8'h10 ;
			data[35400] <= 8'h10 ;
			data[35401] <= 8'h10 ;
			data[35402] <= 8'h10 ;
			data[35403] <= 8'h10 ;
			data[35404] <= 8'h10 ;
			data[35405] <= 8'h10 ;
			data[35406] <= 8'h10 ;
			data[35407] <= 8'h10 ;
			data[35408] <= 8'h10 ;
			data[35409] <= 8'h10 ;
			data[35410] <= 8'h10 ;
			data[35411] <= 8'h10 ;
			data[35412] <= 8'h10 ;
			data[35413] <= 8'h10 ;
			data[35414] <= 8'h10 ;
			data[35415] <= 8'h10 ;
			data[35416] <= 8'h10 ;
			data[35417] <= 8'h10 ;
			data[35418] <= 8'h10 ;
			data[35419] <= 8'h10 ;
			data[35420] <= 8'h10 ;
			data[35421] <= 8'h10 ;
			data[35422] <= 8'h10 ;
			data[35423] <= 8'h10 ;
			data[35424] <= 8'h10 ;
			data[35425] <= 8'h10 ;
			data[35426] <= 8'h10 ;
			data[35427] <= 8'h10 ;
			data[35428] <= 8'h10 ;
			data[35429] <= 8'h10 ;
			data[35430] <= 8'h10 ;
			data[35431] <= 8'h10 ;
			data[35432] <= 8'h10 ;
			data[35433] <= 8'h10 ;
			data[35434] <= 8'h10 ;
			data[35435] <= 8'h10 ;
			data[35436] <= 8'h10 ;
			data[35437] <= 8'h10 ;
			data[35438] <= 8'h10 ;
			data[35439] <= 8'h10 ;
			data[35440] <= 8'h10 ;
			data[35441] <= 8'h10 ;
			data[35442] <= 8'h10 ;
			data[35443] <= 8'h10 ;
			data[35444] <= 8'h10 ;
			data[35445] <= 8'h10 ;
			data[35446] <= 8'h10 ;
			data[35447] <= 8'h10 ;
			data[35448] <= 8'h10 ;
			data[35449] <= 8'h10 ;
			data[35450] <= 8'h10 ;
			data[35451] <= 8'h10 ;
			data[35452] <= 8'h10 ;
			data[35453] <= 8'h10 ;
			data[35454] <= 8'h10 ;
			data[35455] <= 8'h10 ;
			data[35456] <= 8'h10 ;
			data[35457] <= 8'h10 ;
			data[35458] <= 8'h10 ;
			data[35459] <= 8'h10 ;
			data[35460] <= 8'h10 ;
			data[35461] <= 8'h10 ;
			data[35462] <= 8'h10 ;
			data[35463] <= 8'h10 ;
			data[35464] <= 8'h10 ;
			data[35465] <= 8'h10 ;
			data[35466] <= 8'h10 ;
			data[35467] <= 8'h10 ;
			data[35468] <= 8'h10 ;
			data[35469] <= 8'h10 ;
			data[35470] <= 8'h10 ;
			data[35471] <= 8'h10 ;
			data[35472] <= 8'h10 ;
			data[35473] <= 8'h10 ;
			data[35474] <= 8'h10 ;
			data[35475] <= 8'h10 ;
			data[35476] <= 8'h10 ;
			data[35477] <= 8'h10 ;
			data[35478] <= 8'h10 ;
			data[35479] <= 8'h10 ;
			data[35480] <= 8'h10 ;
			data[35481] <= 8'h10 ;
			data[35482] <= 8'h10 ;
			data[35483] <= 8'h10 ;
			data[35484] <= 8'h10 ;
			data[35485] <= 8'h10 ;
			data[35486] <= 8'h10 ;
			data[35487] <= 8'h10 ;
			data[35488] <= 8'h10 ;
			data[35489] <= 8'h10 ;
			data[35490] <= 8'h10 ;
			data[35491] <= 8'h10 ;
			data[35492] <= 8'h10 ;
			data[35493] <= 8'h10 ;
			data[35494] <= 8'h10 ;
			data[35495] <= 8'h10 ;
			data[35496] <= 8'h10 ;
			data[35497] <= 8'h10 ;
			data[35498] <= 8'h10 ;
			data[35499] <= 8'h10 ;
			data[35500] <= 8'h10 ;
			data[35501] <= 8'h10 ;
			data[35502] <= 8'h10 ;
			data[35503] <= 8'h10 ;
			data[35504] <= 8'h10 ;
			data[35505] <= 8'h10 ;
			data[35506] <= 8'h10 ;
			data[35507] <= 8'h10 ;
			data[35508] <= 8'h10 ;
			data[35509] <= 8'h10 ;
			data[35510] <= 8'h10 ;
			data[35511] <= 8'h10 ;
			data[35512] <= 8'h10 ;
			data[35513] <= 8'h10 ;
			data[35514] <= 8'h10 ;
			data[35515] <= 8'h10 ;
			data[35516] <= 8'h10 ;
			data[35517] <= 8'h10 ;
			data[35518] <= 8'h10 ;
			data[35519] <= 8'h10 ;
			data[35520] <= 8'h10 ;
			data[35521] <= 8'h10 ;
			data[35522] <= 8'h10 ;
			data[35523] <= 8'h10 ;
			data[35524] <= 8'h10 ;
			data[35525] <= 8'h10 ;
			data[35526] <= 8'h10 ;
			data[35527] <= 8'h10 ;
			data[35528] <= 8'h10 ;
			data[35529] <= 8'h10 ;
			data[35530] <= 8'h10 ;
			data[35531] <= 8'h10 ;
			data[35532] <= 8'h10 ;
			data[35533] <= 8'h10 ;
			data[35534] <= 8'h10 ;
			data[35535] <= 8'h10 ;
			data[35536] <= 8'h10 ;
			data[35537] <= 8'h10 ;
			data[35538] <= 8'h10 ;
			data[35539] <= 8'h10 ;
			data[35540] <= 8'h10 ;
			data[35541] <= 8'h10 ;
			data[35542] <= 8'h10 ;
			data[35543] <= 8'h10 ;
			data[35544] <= 8'h10 ;
			data[35545] <= 8'h10 ;
			data[35546] <= 8'h10 ;
			data[35547] <= 8'h10 ;
			data[35548] <= 8'h10 ;
			data[35549] <= 8'h10 ;
			data[35550] <= 8'h10 ;
			data[35551] <= 8'h10 ;
			data[35552] <= 8'h10 ;
			data[35553] <= 8'h10 ;
			data[35554] <= 8'h10 ;
			data[35555] <= 8'h10 ;
			data[35556] <= 8'h10 ;
			data[35557] <= 8'h10 ;
			data[35558] <= 8'h10 ;
			data[35559] <= 8'h10 ;
			data[35560] <= 8'h10 ;
			data[35561] <= 8'h10 ;
			data[35562] <= 8'h10 ;
			data[35563] <= 8'h10 ;
			data[35564] <= 8'h10 ;
			data[35565] <= 8'h10 ;
			data[35566] <= 8'h10 ;
			data[35567] <= 8'h10 ;
			data[35568] <= 8'h10 ;
			data[35569] <= 8'h10 ;
			data[35570] <= 8'h10 ;
			data[35571] <= 8'h10 ;
			data[35572] <= 8'h10 ;
			data[35573] <= 8'h10 ;
			data[35574] <= 8'h10 ;
			data[35575] <= 8'h10 ;
			data[35576] <= 8'h10 ;
			data[35577] <= 8'h10 ;
			data[35578] <= 8'h10 ;
			data[35579] <= 8'h10 ;
			data[35580] <= 8'h10 ;
			data[35581] <= 8'h10 ;
			data[35582] <= 8'h10 ;
			data[35583] <= 8'h10 ;
			data[35584] <= 8'h10 ;
			data[35585] <= 8'h10 ;
			data[35586] <= 8'h10 ;
			data[35587] <= 8'h10 ;
			data[35588] <= 8'h10 ;
			data[35589] <= 8'h10 ;
			data[35590] <= 8'h10 ;
			data[35591] <= 8'h10 ;
			data[35592] <= 8'h10 ;
			data[35593] <= 8'h10 ;
			data[35594] <= 8'h10 ;
			data[35595] <= 8'h10 ;
			data[35596] <= 8'h10 ;
			data[35597] <= 8'h10 ;
			data[35598] <= 8'h10 ;
			data[35599] <= 8'h10 ;
			data[35600] <= 8'h10 ;
			data[35601] <= 8'h10 ;
			data[35602] <= 8'h10 ;
			data[35603] <= 8'h10 ;
			data[35604] <= 8'h10 ;
			data[35605] <= 8'h10 ;
			data[35606] <= 8'h10 ;
			data[35607] <= 8'h10 ;
			data[35608] <= 8'h10 ;
			data[35609] <= 8'h10 ;
			data[35610] <= 8'h10 ;
			data[35611] <= 8'h10 ;
			data[35612] <= 8'h10 ;
			data[35613] <= 8'h10 ;
			data[35614] <= 8'h10 ;
			data[35615] <= 8'h10 ;
			data[35616] <= 8'h10 ;
			data[35617] <= 8'h10 ;
			data[35618] <= 8'h10 ;
			data[35619] <= 8'h10 ;
			data[35620] <= 8'h10 ;
			data[35621] <= 8'h10 ;
			data[35622] <= 8'h10 ;
			data[35623] <= 8'h10 ;
			data[35624] <= 8'h10 ;
			data[35625] <= 8'h10 ;
			data[35626] <= 8'h10 ;
			data[35627] <= 8'h10 ;
			data[35628] <= 8'h10 ;
			data[35629] <= 8'h10 ;
			data[35630] <= 8'h10 ;
			data[35631] <= 8'h10 ;
			data[35632] <= 8'h10 ;
			data[35633] <= 8'h10 ;
			data[35634] <= 8'h10 ;
			data[35635] <= 8'h10 ;
			data[35636] <= 8'h10 ;
			data[35637] <= 8'h10 ;
			data[35638] <= 8'h10 ;
			data[35639] <= 8'h10 ;
			data[35640] <= 8'h10 ;
			data[35641] <= 8'h10 ;
			data[35642] <= 8'h10 ;
			data[35643] <= 8'h10 ;
			data[35644] <= 8'h10 ;
			data[35645] <= 8'h10 ;
			data[35646] <= 8'h10 ;
			data[35647] <= 8'h10 ;
			data[35648] <= 8'h10 ;
			data[35649] <= 8'h10 ;
			data[35650] <= 8'h10 ;
			data[35651] <= 8'h10 ;
			data[35652] <= 8'h10 ;
			data[35653] <= 8'h10 ;
			data[35654] <= 8'h10 ;
			data[35655] <= 8'h10 ;
			data[35656] <= 8'h10 ;
			data[35657] <= 8'h10 ;
			data[35658] <= 8'h10 ;
			data[35659] <= 8'h10 ;
			data[35660] <= 8'h10 ;
			data[35661] <= 8'h10 ;
			data[35662] <= 8'h10 ;
			data[35663] <= 8'h10 ;
			data[35664] <= 8'h10 ;
			data[35665] <= 8'h10 ;
			data[35666] <= 8'h10 ;
			data[35667] <= 8'h10 ;
			data[35668] <= 8'h10 ;
			data[35669] <= 8'h10 ;
			data[35670] <= 8'h10 ;
			data[35671] <= 8'h10 ;
			data[35672] <= 8'h10 ;
			data[35673] <= 8'h10 ;
			data[35674] <= 8'h10 ;
			data[35675] <= 8'h10 ;
			data[35676] <= 8'h10 ;
			data[35677] <= 8'h10 ;
			data[35678] <= 8'h10 ;
			data[35679] <= 8'h10 ;
			data[35680] <= 8'h10 ;
			data[35681] <= 8'h10 ;
			data[35682] <= 8'h10 ;
			data[35683] <= 8'h10 ;
			data[35684] <= 8'h10 ;
			data[35685] <= 8'h10 ;
			data[35686] <= 8'h10 ;
			data[35687] <= 8'h10 ;
			data[35688] <= 8'h10 ;
			data[35689] <= 8'h10 ;
			data[35690] <= 8'h10 ;
			data[35691] <= 8'h10 ;
			data[35692] <= 8'h10 ;
			data[35693] <= 8'h10 ;
			data[35694] <= 8'h10 ;
			data[35695] <= 8'h10 ;
			data[35696] <= 8'h10 ;
			data[35697] <= 8'h10 ;
			data[35698] <= 8'h10 ;
			data[35699] <= 8'h10 ;
			data[35700] <= 8'h10 ;
			data[35701] <= 8'h10 ;
			data[35702] <= 8'h10 ;
			data[35703] <= 8'h10 ;
			data[35704] <= 8'h10 ;
			data[35705] <= 8'h10 ;
			data[35706] <= 8'h10 ;
			data[35707] <= 8'h10 ;
			data[35708] <= 8'h10 ;
			data[35709] <= 8'h10 ;
			data[35710] <= 8'h10 ;
			data[35711] <= 8'h10 ;
			data[35712] <= 8'h10 ;
			data[35713] <= 8'h10 ;
			data[35714] <= 8'h10 ;
			data[35715] <= 8'h10 ;
			data[35716] <= 8'h10 ;
			data[35717] <= 8'h10 ;
			data[35718] <= 8'h10 ;
			data[35719] <= 8'h10 ;
			data[35720] <= 8'h10 ;
			data[35721] <= 8'h10 ;
			data[35722] <= 8'h10 ;
			data[35723] <= 8'h10 ;
			data[35724] <= 8'h10 ;
			data[35725] <= 8'h10 ;
			data[35726] <= 8'h10 ;
			data[35727] <= 8'h10 ;
			data[35728] <= 8'h10 ;
			data[35729] <= 8'h10 ;
			data[35730] <= 8'h10 ;
			data[35731] <= 8'h10 ;
			data[35732] <= 8'h10 ;
			data[35733] <= 8'h10 ;
			data[35734] <= 8'h10 ;
			data[35735] <= 8'h10 ;
			data[35736] <= 8'h10 ;
			data[35737] <= 8'h10 ;
			data[35738] <= 8'h10 ;
			data[35739] <= 8'h10 ;
			data[35740] <= 8'h10 ;
			data[35741] <= 8'h10 ;
			data[35742] <= 8'h10 ;
			data[35743] <= 8'h10 ;
			data[35744] <= 8'h10 ;
			data[35745] <= 8'h10 ;
			data[35746] <= 8'h10 ;
			data[35747] <= 8'h10 ;
			data[35748] <= 8'h10 ;
			data[35749] <= 8'h10 ;
			data[35750] <= 8'h10 ;
			data[35751] <= 8'h10 ;
			data[35752] <= 8'h10 ;
			data[35753] <= 8'h10 ;
			data[35754] <= 8'h10 ;
			data[35755] <= 8'h10 ;
			data[35756] <= 8'h10 ;
			data[35757] <= 8'h10 ;
			data[35758] <= 8'h10 ;
			data[35759] <= 8'h10 ;
			data[35760] <= 8'h10 ;
			data[35761] <= 8'h10 ;
			data[35762] <= 8'h10 ;
			data[35763] <= 8'h10 ;
			data[35764] <= 8'h10 ;
			data[35765] <= 8'h10 ;
			data[35766] <= 8'h10 ;
			data[35767] <= 8'h10 ;
			data[35768] <= 8'h10 ;
			data[35769] <= 8'h10 ;
			data[35770] <= 8'h10 ;
			data[35771] <= 8'h10 ;
			data[35772] <= 8'h10 ;
			data[35773] <= 8'h10 ;
			data[35774] <= 8'h10 ;
			data[35775] <= 8'h10 ;
			data[35776] <= 8'h10 ;
			data[35777] <= 8'h10 ;
			data[35778] <= 8'h10 ;
			data[35779] <= 8'h10 ;
			data[35780] <= 8'h10 ;
			data[35781] <= 8'h10 ;
			data[35782] <= 8'h10 ;
			data[35783] <= 8'h10 ;
			data[35784] <= 8'h10 ;
			data[35785] <= 8'h10 ;
			data[35786] <= 8'h10 ;
			data[35787] <= 8'h10 ;
			data[35788] <= 8'h10 ;
			data[35789] <= 8'h10 ;
			data[35790] <= 8'h10 ;
			data[35791] <= 8'h10 ;
			data[35792] <= 8'h10 ;
			data[35793] <= 8'h10 ;
			data[35794] <= 8'h10 ;
			data[35795] <= 8'h10 ;
			data[35796] <= 8'h10 ;
			data[35797] <= 8'h10 ;
			data[35798] <= 8'h10 ;
			data[35799] <= 8'h10 ;
			data[35800] <= 8'h10 ;
			data[35801] <= 8'h10 ;
			data[35802] <= 8'h10 ;
			data[35803] <= 8'h10 ;
			data[35804] <= 8'h10 ;
			data[35805] <= 8'h10 ;
			data[35806] <= 8'h10 ;
			data[35807] <= 8'h10 ;
			data[35808] <= 8'h10 ;
			data[35809] <= 8'h10 ;
			data[35810] <= 8'h10 ;
			data[35811] <= 8'h10 ;
			data[35812] <= 8'h10 ;
			data[35813] <= 8'h10 ;
			data[35814] <= 8'h10 ;
			data[35815] <= 8'h10 ;
			data[35816] <= 8'h10 ;
			data[35817] <= 8'h10 ;
			data[35818] <= 8'h10 ;
			data[35819] <= 8'h10 ;
			data[35820] <= 8'h10 ;
			data[35821] <= 8'h10 ;
			data[35822] <= 8'h10 ;
			data[35823] <= 8'h10 ;
			data[35824] <= 8'h10 ;
			data[35825] <= 8'h10 ;
			data[35826] <= 8'h10 ;
			data[35827] <= 8'h10 ;
			data[35828] <= 8'h10 ;
			data[35829] <= 8'h10 ;
			data[35830] <= 8'h10 ;
			data[35831] <= 8'h10 ;
			data[35832] <= 8'h10 ;
			data[35833] <= 8'h10 ;
			data[35834] <= 8'h10 ;
			data[35835] <= 8'h10 ;
			data[35836] <= 8'h10 ;
			data[35837] <= 8'h10 ;
			data[35838] <= 8'h10 ;
			data[35839] <= 8'h10 ;
			data[35840] <= 8'h10 ;
			data[35841] <= 8'h10 ;
			data[35842] <= 8'h10 ;
			data[35843] <= 8'h10 ;
			data[35844] <= 8'h10 ;
			data[35845] <= 8'h10 ;
			data[35846] <= 8'h10 ;
			data[35847] <= 8'h10 ;
			data[35848] <= 8'h10 ;
			data[35849] <= 8'h10 ;
			data[35850] <= 8'h10 ;
			data[35851] <= 8'h10 ;
			data[35852] <= 8'h10 ;
			data[35853] <= 8'h10 ;
			data[35854] <= 8'h10 ;
			data[35855] <= 8'h10 ;
			data[35856] <= 8'h10 ;
			data[35857] <= 8'h10 ;
			data[35858] <= 8'h10 ;
			data[35859] <= 8'h10 ;
			data[35860] <= 8'h10 ;
			data[35861] <= 8'h10 ;
			data[35862] <= 8'h10 ;
			data[35863] <= 8'h10 ;
			data[35864] <= 8'h10 ;
			data[35865] <= 8'h10 ;
			data[35866] <= 8'h10 ;
			data[35867] <= 8'h10 ;
			data[35868] <= 8'h10 ;
			data[35869] <= 8'h10 ;
			data[35870] <= 8'h10 ;
			data[35871] <= 8'h10 ;
			data[35872] <= 8'h10 ;
			data[35873] <= 8'h10 ;
			data[35874] <= 8'h10 ;
			data[35875] <= 8'h10 ;
			data[35876] <= 8'h10 ;
			data[35877] <= 8'h10 ;
			data[35878] <= 8'h10 ;
			data[35879] <= 8'h10 ;
			data[35880] <= 8'h10 ;
			data[35881] <= 8'h10 ;
			data[35882] <= 8'h10 ;
			data[35883] <= 8'h10 ;
			data[35884] <= 8'h10 ;
			data[35885] <= 8'h10 ;
			data[35886] <= 8'h10 ;
			data[35887] <= 8'h10 ;
			data[35888] <= 8'h10 ;
			data[35889] <= 8'h10 ;
			data[35890] <= 8'h10 ;
			data[35891] <= 8'h10 ;
			data[35892] <= 8'h10 ;
			data[35893] <= 8'h10 ;
			data[35894] <= 8'h10 ;
			data[35895] <= 8'h10 ;
			data[35896] <= 8'h10 ;
			data[35897] <= 8'h10 ;
			data[35898] <= 8'h10 ;
			data[35899] <= 8'h10 ;
			data[35900] <= 8'h10 ;
			data[35901] <= 8'h10 ;
			data[35902] <= 8'h10 ;
			data[35903] <= 8'h10 ;
			data[35904] <= 8'h10 ;
			data[35905] <= 8'h10 ;
			data[35906] <= 8'h10 ;
			data[35907] <= 8'h10 ;
			data[35908] <= 8'h10 ;
			data[35909] <= 8'h10 ;
			data[35910] <= 8'h10 ;
			data[35911] <= 8'h10 ;
			data[35912] <= 8'h10 ;
			data[35913] <= 8'h10 ;
			data[35914] <= 8'h10 ;
			data[35915] <= 8'h10 ;
			data[35916] <= 8'h10 ;
			data[35917] <= 8'h10 ;
			data[35918] <= 8'h10 ;
			data[35919] <= 8'h10 ;
			data[35920] <= 8'h10 ;
			data[35921] <= 8'h10 ;
			data[35922] <= 8'h10 ;
			data[35923] <= 8'h10 ;
			data[35924] <= 8'h10 ;
			data[35925] <= 8'h10 ;
			data[35926] <= 8'h10 ;
			data[35927] <= 8'h10 ;
			data[35928] <= 8'h10 ;
			data[35929] <= 8'h10 ;
			data[35930] <= 8'h10 ;
			data[35931] <= 8'h10 ;
			data[35932] <= 8'h10 ;
			data[35933] <= 8'h10 ;
			data[35934] <= 8'h10 ;
			data[35935] <= 8'h10 ;
			data[35936] <= 8'h10 ;
			data[35937] <= 8'h10 ;
			data[35938] <= 8'h10 ;
			data[35939] <= 8'h10 ;
			data[35940] <= 8'h10 ;
			data[35941] <= 8'h10 ;
			data[35942] <= 8'h10 ;
			data[35943] <= 8'h10 ;
			data[35944] <= 8'h10 ;
			data[35945] <= 8'h10 ;
			data[35946] <= 8'h10 ;
			data[35947] <= 8'h10 ;
			data[35948] <= 8'h10 ;
			data[35949] <= 8'h10 ;
			data[35950] <= 8'h10 ;
			data[35951] <= 8'h10 ;
			data[35952] <= 8'h10 ;
			data[35953] <= 8'h10 ;
			data[35954] <= 8'h10 ;
			data[35955] <= 8'h10 ;
			data[35956] <= 8'h10 ;
			data[35957] <= 8'h10 ;
			data[35958] <= 8'h10 ;
			data[35959] <= 8'h10 ;
			data[35960] <= 8'h10 ;
			data[35961] <= 8'h10 ;
			data[35962] <= 8'h10 ;
			data[35963] <= 8'h10 ;
			data[35964] <= 8'h10 ;
			data[35965] <= 8'h10 ;
			data[35966] <= 8'h10 ;
			data[35967] <= 8'h10 ;
			data[35968] <= 8'h10 ;
			data[35969] <= 8'h10 ;
			data[35970] <= 8'h10 ;
			data[35971] <= 8'h10 ;
			data[35972] <= 8'h10 ;
			data[35973] <= 8'h10 ;
			data[35974] <= 8'h10 ;
			data[35975] <= 8'h10 ;
			data[35976] <= 8'h10 ;
			data[35977] <= 8'h10 ;
			data[35978] <= 8'h10 ;
			data[35979] <= 8'h10 ;
			data[35980] <= 8'h10 ;
			data[35981] <= 8'h10 ;
			data[35982] <= 8'h10 ;
			data[35983] <= 8'h10 ;
			data[35984] <= 8'h10 ;
			data[35985] <= 8'h10 ;
			data[35986] <= 8'h10 ;
			data[35987] <= 8'h10 ;
			data[35988] <= 8'h10 ;
			data[35989] <= 8'h10 ;
			data[35990] <= 8'h10 ;
			data[35991] <= 8'h10 ;
			data[35992] <= 8'h10 ;
			data[35993] <= 8'h10 ;
			data[35994] <= 8'h10 ;
			data[35995] <= 8'h10 ;
			data[35996] <= 8'h10 ;
			data[35997] <= 8'h10 ;
			data[35998] <= 8'h10 ;
			data[35999] <= 8'h10 ;
			data[36000] <= 8'h10 ;
			data[36001] <= 8'h10 ;
			data[36002] <= 8'h10 ;
			data[36003] <= 8'h10 ;
			data[36004] <= 8'h10 ;
			data[36005] <= 8'h10 ;
			data[36006] <= 8'h10 ;
			data[36007] <= 8'h10 ;
			data[36008] <= 8'h10 ;
			data[36009] <= 8'h10 ;
			data[36010] <= 8'h10 ;
			data[36011] <= 8'h10 ;
			data[36012] <= 8'h10 ;
			data[36013] <= 8'h10 ;
			data[36014] <= 8'h10 ;
			data[36015] <= 8'h10 ;
			data[36016] <= 8'h10 ;
			data[36017] <= 8'h10 ;
			data[36018] <= 8'h10 ;
			data[36019] <= 8'h10 ;
			data[36020] <= 8'h10 ;
			data[36021] <= 8'h10 ;
			data[36022] <= 8'h10 ;
			data[36023] <= 8'h10 ;
			data[36024] <= 8'h10 ;
			data[36025] <= 8'h10 ;
			data[36026] <= 8'h10 ;
			data[36027] <= 8'h10 ;
			data[36028] <= 8'h10 ;
			data[36029] <= 8'h10 ;
			data[36030] <= 8'h10 ;
			data[36031] <= 8'h10 ;
			data[36032] <= 8'h10 ;
			data[36033] <= 8'h10 ;
			data[36034] <= 8'h10 ;
			data[36035] <= 8'h10 ;
			data[36036] <= 8'h10 ;
			data[36037] <= 8'h10 ;
			data[36038] <= 8'h10 ;
			data[36039] <= 8'h10 ;
			data[36040] <= 8'h10 ;
			data[36041] <= 8'h10 ;
			data[36042] <= 8'h10 ;
			data[36043] <= 8'h10 ;
			data[36044] <= 8'h10 ;
			data[36045] <= 8'h10 ;
			data[36046] <= 8'h10 ;
			data[36047] <= 8'h10 ;
			data[36048] <= 8'h10 ;
			data[36049] <= 8'h10 ;
			data[36050] <= 8'h10 ;
			data[36051] <= 8'h10 ;
			data[36052] <= 8'h10 ;
			data[36053] <= 8'h10 ;
			data[36054] <= 8'h10 ;
			data[36055] <= 8'h10 ;
			data[36056] <= 8'h10 ;
			data[36057] <= 8'h10 ;
			data[36058] <= 8'h10 ;
			data[36059] <= 8'h10 ;
			data[36060] <= 8'h10 ;
			data[36061] <= 8'h10 ;
			data[36062] <= 8'h10 ;
			data[36063] <= 8'h10 ;
			data[36064] <= 8'h10 ;
			data[36065] <= 8'h10 ;
			data[36066] <= 8'h10 ;
			data[36067] <= 8'h10 ;
			data[36068] <= 8'h10 ;
			data[36069] <= 8'h10 ;
			data[36070] <= 8'h10 ;
			data[36071] <= 8'h10 ;
			data[36072] <= 8'h10 ;
			data[36073] <= 8'h10 ;
			data[36074] <= 8'h10 ;
			data[36075] <= 8'h10 ;
			data[36076] <= 8'h10 ;
			data[36077] <= 8'h10 ;
			data[36078] <= 8'h10 ;
			data[36079] <= 8'h10 ;
			data[36080] <= 8'h10 ;
			data[36081] <= 8'h10 ;
			data[36082] <= 8'h10 ;
			data[36083] <= 8'h10 ;
			data[36084] <= 8'h10 ;
			data[36085] <= 8'h10 ;
			data[36086] <= 8'h10 ;
			data[36087] <= 8'h10 ;
			data[36088] <= 8'h10 ;
			data[36089] <= 8'h10 ;
			data[36090] <= 8'h10 ;
			data[36091] <= 8'h10 ;
			data[36092] <= 8'h10 ;
			data[36093] <= 8'h10 ;
			data[36094] <= 8'h10 ;
			data[36095] <= 8'h10 ;
			data[36096] <= 8'h10 ;
			data[36097] <= 8'h10 ;
			data[36098] <= 8'h10 ;
			data[36099] <= 8'h10 ;
			data[36100] <= 8'h10 ;
			data[36101] <= 8'h10 ;
			data[36102] <= 8'h10 ;
			data[36103] <= 8'h10 ;
			data[36104] <= 8'h10 ;
			data[36105] <= 8'h10 ;
			data[36106] <= 8'h10 ;
			data[36107] <= 8'h10 ;
			data[36108] <= 8'h10 ;
			data[36109] <= 8'h10 ;
			data[36110] <= 8'h10 ;
			data[36111] <= 8'h10 ;
			data[36112] <= 8'h10 ;
			data[36113] <= 8'h10 ;
			data[36114] <= 8'h10 ;
			data[36115] <= 8'h10 ;
			data[36116] <= 8'h10 ;
			data[36117] <= 8'h10 ;
			data[36118] <= 8'h10 ;
			data[36119] <= 8'h10 ;
			data[36120] <= 8'h10 ;
			data[36121] <= 8'h10 ;
			data[36122] <= 8'h10 ;
			data[36123] <= 8'h10 ;
			data[36124] <= 8'h10 ;
			data[36125] <= 8'h10 ;
			data[36126] <= 8'h10 ;
			data[36127] <= 8'h10 ;
			data[36128] <= 8'h10 ;
			data[36129] <= 8'h10 ;
			data[36130] <= 8'h10 ;
			data[36131] <= 8'h10 ;
			data[36132] <= 8'h10 ;
			data[36133] <= 8'h10 ;
			data[36134] <= 8'h10 ;
			data[36135] <= 8'h10 ;
			data[36136] <= 8'h10 ;
			data[36137] <= 8'h10 ;
			data[36138] <= 8'h10 ;
			data[36139] <= 8'h10 ;
			data[36140] <= 8'h10 ;
			data[36141] <= 8'h10 ;
			data[36142] <= 8'h10 ;
			data[36143] <= 8'h10 ;
			data[36144] <= 8'h10 ;
			data[36145] <= 8'h10 ;
			data[36146] <= 8'h10 ;
			data[36147] <= 8'h10 ;
			data[36148] <= 8'h10 ;
			data[36149] <= 8'h10 ;
			data[36150] <= 8'h10 ;
			data[36151] <= 8'h10 ;
			data[36152] <= 8'h10 ;
			data[36153] <= 8'h10 ;
			data[36154] <= 8'h10 ;
			data[36155] <= 8'h10 ;
			data[36156] <= 8'h10 ;
			data[36157] <= 8'h10 ;
			data[36158] <= 8'h10 ;
			data[36159] <= 8'h10 ;
			data[36160] <= 8'h10 ;
			data[36161] <= 8'h10 ;
			data[36162] <= 8'h10 ;
			data[36163] <= 8'h10 ;
			data[36164] <= 8'h10 ;
			data[36165] <= 8'h10 ;
			data[36166] <= 8'h10 ;
			data[36167] <= 8'h10 ;
			data[36168] <= 8'h10 ;
			data[36169] <= 8'h10 ;
			data[36170] <= 8'h10 ;
			data[36171] <= 8'h10 ;
			data[36172] <= 8'h10 ;
			data[36173] <= 8'h10 ;
			data[36174] <= 8'h10 ;
			data[36175] <= 8'h10 ;
			data[36176] <= 8'h10 ;
			data[36177] <= 8'h10 ;
			data[36178] <= 8'h10 ;
			data[36179] <= 8'h10 ;
			data[36180] <= 8'h10 ;
			data[36181] <= 8'h10 ;
			data[36182] <= 8'h10 ;
			data[36183] <= 8'h10 ;
			data[36184] <= 8'h10 ;
			data[36185] <= 8'h10 ;
			data[36186] <= 8'h10 ;
			data[36187] <= 8'h10 ;
			data[36188] <= 8'h10 ;
			data[36189] <= 8'h10 ;
			data[36190] <= 8'h10 ;
			data[36191] <= 8'h10 ;
			data[36192] <= 8'h10 ;
			data[36193] <= 8'h10 ;
			data[36194] <= 8'h10 ;
			data[36195] <= 8'h10 ;
			data[36196] <= 8'h10 ;
			data[36197] <= 8'h10 ;
			data[36198] <= 8'h10 ;
			data[36199] <= 8'h10 ;
			data[36200] <= 8'h10 ;
			data[36201] <= 8'h10 ;
			data[36202] <= 8'h10 ;
			data[36203] <= 8'h10 ;
			data[36204] <= 8'h10 ;
			data[36205] <= 8'h10 ;
			data[36206] <= 8'h10 ;
			data[36207] <= 8'h10 ;
			data[36208] <= 8'h10 ;
			data[36209] <= 8'h10 ;
			data[36210] <= 8'h10 ;
			data[36211] <= 8'h10 ;
			data[36212] <= 8'h10 ;
			data[36213] <= 8'h10 ;
			data[36214] <= 8'h10 ;
			data[36215] <= 8'h10 ;
			data[36216] <= 8'h10 ;
			data[36217] <= 8'h10 ;
			data[36218] <= 8'h10 ;
			data[36219] <= 8'h10 ;
			data[36220] <= 8'h10 ;
			data[36221] <= 8'h10 ;
			data[36222] <= 8'h10 ;
			data[36223] <= 8'h10 ;
			data[36224] <= 8'h10 ;
			data[36225] <= 8'h10 ;
			data[36226] <= 8'h10 ;
			data[36227] <= 8'h10 ;
			data[36228] <= 8'h10 ;
			data[36229] <= 8'h10 ;
			data[36230] <= 8'h10 ;
			data[36231] <= 8'h10 ;
			data[36232] <= 8'h10 ;
			data[36233] <= 8'h10 ;
			data[36234] <= 8'h10 ;
			data[36235] <= 8'h10 ;
			data[36236] <= 8'h10 ;
			data[36237] <= 8'h10 ;
			data[36238] <= 8'h10 ;
			data[36239] <= 8'h10 ;
			data[36240] <= 8'h10 ;
			data[36241] <= 8'h10 ;
			data[36242] <= 8'h10 ;
			data[36243] <= 8'h10 ;
			data[36244] <= 8'h10 ;
			data[36245] <= 8'h10 ;
			data[36246] <= 8'h10 ;
			data[36247] <= 8'h10 ;
			data[36248] <= 8'h10 ;
			data[36249] <= 8'h10 ;
			data[36250] <= 8'h10 ;
			data[36251] <= 8'h10 ;
			data[36252] <= 8'h10 ;
			data[36253] <= 8'h10 ;
			data[36254] <= 8'h10 ;
			data[36255] <= 8'h10 ;
			data[36256] <= 8'h10 ;
			data[36257] <= 8'h10 ;
			data[36258] <= 8'h10 ;
			data[36259] <= 8'h10 ;
			data[36260] <= 8'h10 ;
			data[36261] <= 8'h10 ;
			data[36262] <= 8'h10 ;
			data[36263] <= 8'h10 ;
			data[36264] <= 8'h10 ;
			data[36265] <= 8'h10 ;
			data[36266] <= 8'h10 ;
			data[36267] <= 8'h10 ;
			data[36268] <= 8'h10 ;
			data[36269] <= 8'h10 ;
			data[36270] <= 8'h10 ;
			data[36271] <= 8'h10 ;
			data[36272] <= 8'h10 ;
			data[36273] <= 8'h10 ;
			data[36274] <= 8'h10 ;
			data[36275] <= 8'h10 ;
			data[36276] <= 8'h10 ;
			data[36277] <= 8'h10 ;
			data[36278] <= 8'h10 ;
			data[36279] <= 8'h10 ;
			data[36280] <= 8'h10 ;
			data[36281] <= 8'h10 ;
			data[36282] <= 8'h10 ;
			data[36283] <= 8'h10 ;
			data[36284] <= 8'h10 ;
			data[36285] <= 8'h10 ;
			data[36286] <= 8'h10 ;
			data[36287] <= 8'h10 ;
			data[36288] <= 8'h10 ;
			data[36289] <= 8'h10 ;
			data[36290] <= 8'h10 ;
			data[36291] <= 8'h10 ;
			data[36292] <= 8'h10 ;
			data[36293] <= 8'h10 ;
			data[36294] <= 8'h10 ;
			data[36295] <= 8'h10 ;
			data[36296] <= 8'h10 ;
			data[36297] <= 8'h10 ;
			data[36298] <= 8'h10 ;
			data[36299] <= 8'h10 ;
			data[36300] <= 8'h10 ;
			data[36301] <= 8'h10 ;
			data[36302] <= 8'h10 ;
			data[36303] <= 8'h10 ;
			data[36304] <= 8'h10 ;
			data[36305] <= 8'h10 ;
			data[36306] <= 8'h10 ;
			data[36307] <= 8'h10 ;
			data[36308] <= 8'h10 ;
			data[36309] <= 8'h10 ;
			data[36310] <= 8'h10 ;
			data[36311] <= 8'h10 ;
			data[36312] <= 8'h10 ;
			data[36313] <= 8'h10 ;
			data[36314] <= 8'h10 ;
			data[36315] <= 8'h10 ;
			data[36316] <= 8'h10 ;
			data[36317] <= 8'h10 ;
			data[36318] <= 8'h10 ;
			data[36319] <= 8'h10 ;
			data[36320] <= 8'h10 ;
			data[36321] <= 8'h10 ;
			data[36322] <= 8'h10 ;
			data[36323] <= 8'h10 ;
			data[36324] <= 8'h10 ;
			data[36325] <= 8'h10 ;
			data[36326] <= 8'h10 ;
			data[36327] <= 8'h10 ;
			data[36328] <= 8'h10 ;
			data[36329] <= 8'h10 ;
			data[36330] <= 8'h10 ;
			data[36331] <= 8'h10 ;
			data[36332] <= 8'h10 ;
			data[36333] <= 8'h10 ;
			data[36334] <= 8'h10 ;
			data[36335] <= 8'h10 ;
			data[36336] <= 8'h10 ;
			data[36337] <= 8'h10 ;
			data[36338] <= 8'h10 ;
			data[36339] <= 8'h10 ;
			data[36340] <= 8'h10 ;
			data[36341] <= 8'h10 ;
			data[36342] <= 8'h10 ;
			data[36343] <= 8'h10 ;
			data[36344] <= 8'h10 ;
			data[36345] <= 8'h10 ;
			data[36346] <= 8'h10 ;
			data[36347] <= 8'h10 ;
			data[36348] <= 8'h10 ;
			data[36349] <= 8'h10 ;
			data[36350] <= 8'h10 ;
			data[36351] <= 8'h10 ;
			data[36352] <= 8'h10 ;
			data[36353] <= 8'h10 ;
			data[36354] <= 8'h10 ;
			data[36355] <= 8'h10 ;
			data[36356] <= 8'h10 ;
			data[36357] <= 8'h10 ;
			data[36358] <= 8'h10 ;
			data[36359] <= 8'h10 ;
			data[36360] <= 8'h10 ;
			data[36361] <= 8'h10 ;
			data[36362] <= 8'h10 ;
			data[36363] <= 8'h10 ;
			data[36364] <= 8'h10 ;
			data[36365] <= 8'h10 ;
			data[36366] <= 8'h10 ;
			data[36367] <= 8'h10 ;
			data[36368] <= 8'h10 ;
			data[36369] <= 8'h10 ;
			data[36370] <= 8'h10 ;
			data[36371] <= 8'h10 ;
			data[36372] <= 8'h10 ;
			data[36373] <= 8'h10 ;
			data[36374] <= 8'h10 ;
			data[36375] <= 8'h10 ;
			data[36376] <= 8'h10 ;
			data[36377] <= 8'h10 ;
			data[36378] <= 8'h10 ;
			data[36379] <= 8'h10 ;
			data[36380] <= 8'h10 ;
			data[36381] <= 8'h10 ;
			data[36382] <= 8'h10 ;
			data[36383] <= 8'h10 ;
			data[36384] <= 8'h10 ;
			data[36385] <= 8'h10 ;
			data[36386] <= 8'h10 ;
			data[36387] <= 8'h10 ;
			data[36388] <= 8'h10 ;
			data[36389] <= 8'h10 ;
			data[36390] <= 8'h10 ;
			data[36391] <= 8'h10 ;
			data[36392] <= 8'h10 ;
			data[36393] <= 8'h10 ;
			data[36394] <= 8'h10 ;
			data[36395] <= 8'h10 ;
			data[36396] <= 8'h10 ;
			data[36397] <= 8'h10 ;
			data[36398] <= 8'h10 ;
			data[36399] <= 8'h10 ;
			data[36400] <= 8'h10 ;
			data[36401] <= 8'h10 ;
			data[36402] <= 8'h10 ;
			data[36403] <= 8'h10 ;
			data[36404] <= 8'h10 ;
			data[36405] <= 8'h10 ;
			data[36406] <= 8'h10 ;
			data[36407] <= 8'h10 ;
			data[36408] <= 8'h10 ;
			data[36409] <= 8'h10 ;
			data[36410] <= 8'h10 ;
			data[36411] <= 8'h10 ;
			data[36412] <= 8'h10 ;
			data[36413] <= 8'h10 ;
			data[36414] <= 8'h10 ;
			data[36415] <= 8'h10 ;
			data[36416] <= 8'h10 ;
			data[36417] <= 8'h10 ;
			data[36418] <= 8'h10 ;
			data[36419] <= 8'h10 ;
			data[36420] <= 8'h10 ;
			data[36421] <= 8'h10 ;
			data[36422] <= 8'h10 ;
			data[36423] <= 8'h10 ;
			data[36424] <= 8'h10 ;
			data[36425] <= 8'h10 ;
			data[36426] <= 8'h10 ;
			data[36427] <= 8'h10 ;
			data[36428] <= 8'h10 ;
			data[36429] <= 8'h10 ;
			data[36430] <= 8'h10 ;
			data[36431] <= 8'h10 ;
			data[36432] <= 8'h10 ;
			data[36433] <= 8'h10 ;
			data[36434] <= 8'h10 ;
			data[36435] <= 8'h10 ;
			data[36436] <= 8'h10 ;
			data[36437] <= 8'h10 ;
			data[36438] <= 8'h10 ;
			data[36439] <= 8'h10 ;
			data[36440] <= 8'h10 ;
			data[36441] <= 8'h10 ;
			data[36442] <= 8'h10 ;
			data[36443] <= 8'h10 ;
			data[36444] <= 8'h10 ;
			data[36445] <= 8'h10 ;
			data[36446] <= 8'h10 ;
			data[36447] <= 8'h10 ;
			data[36448] <= 8'h10 ;
			data[36449] <= 8'h10 ;
			data[36450] <= 8'h10 ;
			data[36451] <= 8'h10 ;
			data[36452] <= 8'h10 ;
			data[36453] <= 8'h10 ;
			data[36454] <= 8'h10 ;
			data[36455] <= 8'h10 ;
			data[36456] <= 8'h10 ;
			data[36457] <= 8'h10 ;
			data[36458] <= 8'h10 ;
			data[36459] <= 8'h10 ;
			data[36460] <= 8'h10 ;
			data[36461] <= 8'h10 ;
			data[36462] <= 8'h10 ;
			data[36463] <= 8'h10 ;
			data[36464] <= 8'h10 ;
			data[36465] <= 8'h10 ;
			data[36466] <= 8'h10 ;
			data[36467] <= 8'h10 ;
			data[36468] <= 8'h10 ;
			data[36469] <= 8'h10 ;
			data[36470] <= 8'h10 ;
			data[36471] <= 8'h10 ;
			data[36472] <= 8'h10 ;
			data[36473] <= 8'h10 ;
			data[36474] <= 8'h10 ;
			data[36475] <= 8'h10 ;
			data[36476] <= 8'h10 ;
			data[36477] <= 8'h10 ;
			data[36478] <= 8'h10 ;
			data[36479] <= 8'h10 ;
			data[36480] <= 8'h10 ;
			data[36481] <= 8'h10 ;
			data[36482] <= 8'h10 ;
			data[36483] <= 8'h10 ;
			data[36484] <= 8'h10 ;
			data[36485] <= 8'h10 ;
			data[36486] <= 8'h10 ;
			data[36487] <= 8'h10 ;
			data[36488] <= 8'h10 ;
			data[36489] <= 8'h10 ;
			data[36490] <= 8'h10 ;
			data[36491] <= 8'h10 ;
			data[36492] <= 8'h10 ;
			data[36493] <= 8'h10 ;
			data[36494] <= 8'h10 ;
			data[36495] <= 8'h10 ;
			data[36496] <= 8'h10 ;
			data[36497] <= 8'h10 ;
			data[36498] <= 8'h10 ;
			data[36499] <= 8'h10 ;
			data[36500] <= 8'h10 ;
			data[36501] <= 8'h10 ;
			data[36502] <= 8'h10 ;
			data[36503] <= 8'h10 ;
			data[36504] <= 8'h10 ;
			data[36505] <= 8'h10 ;
			data[36506] <= 8'h10 ;
			data[36507] <= 8'h10 ;
			data[36508] <= 8'h10 ;
			data[36509] <= 8'h10 ;
			data[36510] <= 8'h10 ;
			data[36511] <= 8'h10 ;
			data[36512] <= 8'h10 ;
			data[36513] <= 8'h10 ;
			data[36514] <= 8'h10 ;
			data[36515] <= 8'h10 ;
			data[36516] <= 8'h10 ;
			data[36517] <= 8'h10 ;
			data[36518] <= 8'h10 ;
			data[36519] <= 8'h10 ;
			data[36520] <= 8'h10 ;
			data[36521] <= 8'h10 ;
			data[36522] <= 8'h10 ;
			data[36523] <= 8'h10 ;
			data[36524] <= 8'h10 ;
			data[36525] <= 8'h10 ;
			data[36526] <= 8'h10 ;
			data[36527] <= 8'h10 ;
			data[36528] <= 8'h10 ;
			data[36529] <= 8'h10 ;
			data[36530] <= 8'h10 ;
			data[36531] <= 8'h10 ;
			data[36532] <= 8'h10 ;
			data[36533] <= 8'h10 ;
			data[36534] <= 8'h10 ;
			data[36535] <= 8'h10 ;
			data[36536] <= 8'h10 ;
			data[36537] <= 8'h10 ;
			data[36538] <= 8'h10 ;
			data[36539] <= 8'h10 ;
			data[36540] <= 8'h10 ;
			data[36541] <= 8'h10 ;
			data[36542] <= 8'h10 ;
			data[36543] <= 8'h10 ;
			data[36544] <= 8'h10 ;
			data[36545] <= 8'h10 ;
			data[36546] <= 8'h10 ;
			data[36547] <= 8'h10 ;
			data[36548] <= 8'h10 ;
			data[36549] <= 8'h10 ;
			data[36550] <= 8'h10 ;
			data[36551] <= 8'h10 ;
			data[36552] <= 8'h10 ;
			data[36553] <= 8'h10 ;
			data[36554] <= 8'h10 ;
			data[36555] <= 8'h10 ;
			data[36556] <= 8'h10 ;
			data[36557] <= 8'h10 ;
			data[36558] <= 8'h10 ;
			data[36559] <= 8'h10 ;
			data[36560] <= 8'h10 ;
			data[36561] <= 8'h10 ;
			data[36562] <= 8'h10 ;
			data[36563] <= 8'h10 ;
			data[36564] <= 8'h10 ;
			data[36565] <= 8'h10 ;
			data[36566] <= 8'h10 ;
			data[36567] <= 8'h10 ;
			data[36568] <= 8'h10 ;
			data[36569] <= 8'h10 ;
			data[36570] <= 8'h10 ;
			data[36571] <= 8'h10 ;
			data[36572] <= 8'h10 ;
			data[36573] <= 8'h10 ;
			data[36574] <= 8'h10 ;
			data[36575] <= 8'h10 ;
			data[36576] <= 8'h10 ;
			data[36577] <= 8'h10 ;
			data[36578] <= 8'h10 ;
			data[36579] <= 8'h10 ;
			data[36580] <= 8'h10 ;
			data[36581] <= 8'h10 ;
			data[36582] <= 8'h10 ;
			data[36583] <= 8'h10 ;
			data[36584] <= 8'h10 ;
			data[36585] <= 8'h10 ;
			data[36586] <= 8'h10 ;
			data[36587] <= 8'h10 ;
			data[36588] <= 8'h10 ;
			data[36589] <= 8'h10 ;
			data[36590] <= 8'h10 ;
			data[36591] <= 8'h10 ;
			data[36592] <= 8'h10 ;
			data[36593] <= 8'h10 ;
			data[36594] <= 8'h10 ;
			data[36595] <= 8'h10 ;
			data[36596] <= 8'h10 ;
			data[36597] <= 8'h10 ;
			data[36598] <= 8'h10 ;
			data[36599] <= 8'h10 ;
			data[36600] <= 8'h10 ;
			data[36601] <= 8'h10 ;
			data[36602] <= 8'h10 ;
			data[36603] <= 8'h10 ;
			data[36604] <= 8'h10 ;
			data[36605] <= 8'h10 ;
			data[36606] <= 8'h10 ;
			data[36607] <= 8'h10 ;
			data[36608] <= 8'h10 ;
			data[36609] <= 8'h10 ;
			data[36610] <= 8'h10 ;
			data[36611] <= 8'h10 ;
			data[36612] <= 8'h10 ;
			data[36613] <= 8'h10 ;
			data[36614] <= 8'h10 ;
			data[36615] <= 8'h10 ;
			data[36616] <= 8'h10 ;
			data[36617] <= 8'h10 ;
			data[36618] <= 8'h10 ;
			data[36619] <= 8'h10 ;
			data[36620] <= 8'h10 ;
			data[36621] <= 8'h10 ;
			data[36622] <= 8'h10 ;
			data[36623] <= 8'h10 ;
			data[36624] <= 8'h10 ;
			data[36625] <= 8'h10 ;
			data[36626] <= 8'h10 ;
			data[36627] <= 8'h10 ;
			data[36628] <= 8'h10 ;
			data[36629] <= 8'h10 ;
			data[36630] <= 8'h10 ;
			data[36631] <= 8'h10 ;
			data[36632] <= 8'h10 ;
			data[36633] <= 8'h10 ;
			data[36634] <= 8'h10 ;
			data[36635] <= 8'h10 ;
			data[36636] <= 8'h10 ;
			data[36637] <= 8'h10 ;
			data[36638] <= 8'h10 ;
			data[36639] <= 8'h10 ;
			data[36640] <= 8'h10 ;
			data[36641] <= 8'h10 ;
			data[36642] <= 8'h10 ;
			data[36643] <= 8'h10 ;
			data[36644] <= 8'h10 ;
			data[36645] <= 8'h10 ;
			data[36646] <= 8'h10 ;
			data[36647] <= 8'h10 ;
			data[36648] <= 8'h10 ;
			data[36649] <= 8'h10 ;
			data[36650] <= 8'h10 ;
			data[36651] <= 8'h10 ;
			data[36652] <= 8'h10 ;
			data[36653] <= 8'h10 ;
			data[36654] <= 8'h10 ;
			data[36655] <= 8'h10 ;
			data[36656] <= 8'h10 ;
			data[36657] <= 8'h10 ;
			data[36658] <= 8'h10 ;
			data[36659] <= 8'h10 ;
			data[36660] <= 8'h10 ;
			data[36661] <= 8'h10 ;
			data[36662] <= 8'h10 ;
			data[36663] <= 8'h10 ;
			data[36664] <= 8'h10 ;
			data[36665] <= 8'h10 ;
			data[36666] <= 8'h10 ;
			data[36667] <= 8'h10 ;
			data[36668] <= 8'h10 ;
			data[36669] <= 8'h10 ;
			data[36670] <= 8'h10 ;
			data[36671] <= 8'h10 ;
			data[36672] <= 8'h10 ;
			data[36673] <= 8'h10 ;
			data[36674] <= 8'h10 ;
			data[36675] <= 8'h10 ;
			data[36676] <= 8'h10 ;
			data[36677] <= 8'h10 ;
			data[36678] <= 8'h10 ;
			data[36679] <= 8'h10 ;
			data[36680] <= 8'h10 ;
			data[36681] <= 8'h10 ;
			data[36682] <= 8'h10 ;
			data[36683] <= 8'h10 ;
			data[36684] <= 8'h10 ;
			data[36685] <= 8'h10 ;
			data[36686] <= 8'h10 ;
			data[36687] <= 8'h10 ;
			data[36688] <= 8'h10 ;
			data[36689] <= 8'h10 ;
			data[36690] <= 8'h10 ;
			data[36691] <= 8'h10 ;
			data[36692] <= 8'h10 ;
			data[36693] <= 8'h10 ;
			data[36694] <= 8'h10 ;
			data[36695] <= 8'h10 ;
			data[36696] <= 8'h10 ;
			data[36697] <= 8'h10 ;
			data[36698] <= 8'h10 ;
			data[36699] <= 8'h10 ;
			data[36700] <= 8'h10 ;
			data[36701] <= 8'h10 ;
			data[36702] <= 8'h10 ;
			data[36703] <= 8'h10 ;
			data[36704] <= 8'h10 ;
			data[36705] <= 8'h10 ;
			data[36706] <= 8'h10 ;
			data[36707] <= 8'h10 ;
			data[36708] <= 8'h10 ;
			data[36709] <= 8'h10 ;
			data[36710] <= 8'h10 ;
			data[36711] <= 8'h10 ;
			data[36712] <= 8'h10 ;
			data[36713] <= 8'h10 ;
			data[36714] <= 8'h10 ;
			data[36715] <= 8'h10 ;
			data[36716] <= 8'h10 ;
			data[36717] <= 8'h10 ;
			data[36718] <= 8'h10 ;
			data[36719] <= 8'h10 ;
			data[36720] <= 8'h10 ;
			data[36721] <= 8'h10 ;
			data[36722] <= 8'h10 ;
			data[36723] <= 8'h10 ;
			data[36724] <= 8'h10 ;
			data[36725] <= 8'h10 ;
			data[36726] <= 8'h10 ;
			data[36727] <= 8'h10 ;
			data[36728] <= 8'h10 ;
			data[36729] <= 8'h10 ;
			data[36730] <= 8'h10 ;
			data[36731] <= 8'h10 ;
			data[36732] <= 8'h10 ;
			data[36733] <= 8'h10 ;
			data[36734] <= 8'h10 ;
			data[36735] <= 8'h10 ;
			data[36736] <= 8'h10 ;
			data[36737] <= 8'h10 ;
			data[36738] <= 8'h10 ;
			data[36739] <= 8'h10 ;
			data[36740] <= 8'h10 ;
			data[36741] <= 8'h10 ;
			data[36742] <= 8'h10 ;
			data[36743] <= 8'h10 ;
			data[36744] <= 8'h10 ;
			data[36745] <= 8'h10 ;
			data[36746] <= 8'h10 ;
			data[36747] <= 8'h10 ;
			data[36748] <= 8'h10 ;
			data[36749] <= 8'h10 ;
			data[36750] <= 8'h10 ;
			data[36751] <= 8'h10 ;
			data[36752] <= 8'h10 ;
			data[36753] <= 8'h10 ;
			data[36754] <= 8'h10 ;
			data[36755] <= 8'h10 ;
			data[36756] <= 8'h10 ;
			data[36757] <= 8'h10 ;
			data[36758] <= 8'h10 ;
			data[36759] <= 8'h10 ;
			data[36760] <= 8'h10 ;
			data[36761] <= 8'h10 ;
			data[36762] <= 8'h10 ;
			data[36763] <= 8'h10 ;
			data[36764] <= 8'h10 ;
			data[36765] <= 8'h10 ;
			data[36766] <= 8'h10 ;
			data[36767] <= 8'h10 ;
			data[36768] <= 8'h10 ;
			data[36769] <= 8'h10 ;
			data[36770] <= 8'h10 ;
			data[36771] <= 8'h10 ;
			data[36772] <= 8'h10 ;
			data[36773] <= 8'h10 ;
			data[36774] <= 8'h10 ;
			data[36775] <= 8'h10 ;
			data[36776] <= 8'h10 ;
			data[36777] <= 8'h10 ;
			data[36778] <= 8'h10 ;
			data[36779] <= 8'h10 ;
			data[36780] <= 8'h10 ;
			data[36781] <= 8'h10 ;
			data[36782] <= 8'h10 ;
			data[36783] <= 8'h10 ;
			data[36784] <= 8'h10 ;
			data[36785] <= 8'h10 ;
			data[36786] <= 8'h10 ;
			data[36787] <= 8'h10 ;
			data[36788] <= 8'h10 ;
			data[36789] <= 8'h10 ;
			data[36790] <= 8'h10 ;
			data[36791] <= 8'h10 ;
			data[36792] <= 8'h10 ;
			data[36793] <= 8'h10 ;
			data[36794] <= 8'h10 ;
			data[36795] <= 8'h10 ;
			data[36796] <= 8'h10 ;
			data[36797] <= 8'h10 ;
			data[36798] <= 8'h10 ;
			data[36799] <= 8'h10 ;
			data[36800] <= 8'h10 ;
			data[36801] <= 8'h10 ;
			data[36802] <= 8'h10 ;
			data[36803] <= 8'h10 ;
			data[36804] <= 8'h10 ;
			data[36805] <= 8'h10 ;
			data[36806] <= 8'h10 ;
			data[36807] <= 8'h10 ;
			data[36808] <= 8'h10 ;
			data[36809] <= 8'h10 ;
			data[36810] <= 8'h10 ;
			data[36811] <= 8'h10 ;
			data[36812] <= 8'h10 ;
			data[36813] <= 8'h10 ;
			data[36814] <= 8'h10 ;
			data[36815] <= 8'h10 ;
			data[36816] <= 8'h10 ;
			data[36817] <= 8'h10 ;
			data[36818] <= 8'h10 ;
			data[36819] <= 8'h10 ;
			data[36820] <= 8'h10 ;
			data[36821] <= 8'h10 ;
			data[36822] <= 8'h10 ;
			data[36823] <= 8'h10 ;
			data[36824] <= 8'h10 ;
			data[36825] <= 8'h10 ;
			data[36826] <= 8'h10 ;
			data[36827] <= 8'h10 ;
			data[36828] <= 8'h10 ;
			data[36829] <= 8'h10 ;
			data[36830] <= 8'h10 ;
			data[36831] <= 8'h10 ;
			data[36832] <= 8'h10 ;
			data[36833] <= 8'h10 ;
			data[36834] <= 8'h10 ;
			data[36835] <= 8'h10 ;
			data[36836] <= 8'h10 ;
			data[36837] <= 8'h10 ;
			data[36838] <= 8'h10 ;
			data[36839] <= 8'h10 ;
			data[36840] <= 8'h10 ;
			data[36841] <= 8'h10 ;
			data[36842] <= 8'h10 ;
			data[36843] <= 8'h10 ;
			data[36844] <= 8'h10 ;
			data[36845] <= 8'h10 ;
			data[36846] <= 8'h10 ;
			data[36847] <= 8'h10 ;
			data[36848] <= 8'h10 ;
			data[36849] <= 8'h10 ;
			data[36850] <= 8'h10 ;
			data[36851] <= 8'h10 ;
			data[36852] <= 8'h10 ;
			data[36853] <= 8'h10 ;
			data[36854] <= 8'h10 ;
			data[36855] <= 8'h10 ;
			data[36856] <= 8'h10 ;
			data[36857] <= 8'h10 ;
			data[36858] <= 8'h10 ;
			data[36859] <= 8'h10 ;
			data[36860] <= 8'h10 ;
			data[36861] <= 8'h10 ;
			data[36862] <= 8'h10 ;
			data[36863] <= 8'h10 ;
			data[36864] <= 8'h10 ;
			data[36865] <= 8'h10 ;
			data[36866] <= 8'h10 ;
			data[36867] <= 8'h10 ;
			data[36868] <= 8'h10 ;
			data[36869] <= 8'h10 ;
			data[36870] <= 8'h10 ;
			data[36871] <= 8'h10 ;
			data[36872] <= 8'h10 ;
			data[36873] <= 8'h10 ;
			data[36874] <= 8'h10 ;
			data[36875] <= 8'h10 ;
			data[36876] <= 8'h10 ;
			data[36877] <= 8'h10 ;
			data[36878] <= 8'h10 ;
			data[36879] <= 8'h10 ;
			data[36880] <= 8'h10 ;
			data[36881] <= 8'h10 ;
			data[36882] <= 8'h10 ;
			data[36883] <= 8'h10 ;
			data[36884] <= 8'h10 ;
			data[36885] <= 8'h10 ;
			data[36886] <= 8'h10 ;
			data[36887] <= 8'h10 ;
			data[36888] <= 8'h10 ;
			data[36889] <= 8'h10 ;
			data[36890] <= 8'h10 ;
			data[36891] <= 8'h10 ;
			data[36892] <= 8'h10 ;
			data[36893] <= 8'h10 ;
			data[36894] <= 8'h10 ;
			data[36895] <= 8'h10 ;
			data[36896] <= 8'h10 ;
			data[36897] <= 8'h10 ;
			data[36898] <= 8'h10 ;
			data[36899] <= 8'h10 ;
			data[36900] <= 8'h10 ;
			data[36901] <= 8'h10 ;
			data[36902] <= 8'h10 ;
			data[36903] <= 8'h10 ;
			data[36904] <= 8'h10 ;
			data[36905] <= 8'h10 ;
			data[36906] <= 8'h10 ;
			data[36907] <= 8'h10 ;
			data[36908] <= 8'h10 ;
			data[36909] <= 8'h10 ;
			data[36910] <= 8'h10 ;
			data[36911] <= 8'h10 ;
			data[36912] <= 8'h10 ;
			data[36913] <= 8'h10 ;
			data[36914] <= 8'h10 ;
			data[36915] <= 8'h10 ;
			data[36916] <= 8'h10 ;
			data[36917] <= 8'h10 ;
			data[36918] <= 8'h10 ;
			data[36919] <= 8'h10 ;
			data[36920] <= 8'h10 ;
			data[36921] <= 8'h10 ;
			data[36922] <= 8'h10 ;
			data[36923] <= 8'h10 ;
			data[36924] <= 8'h10 ;
			data[36925] <= 8'h10 ;
			data[36926] <= 8'h10 ;
			data[36927] <= 8'h10 ;
			data[36928] <= 8'h10 ;
			data[36929] <= 8'h10 ;
			data[36930] <= 8'h10 ;
			data[36931] <= 8'h10 ;
			data[36932] <= 8'h10 ;
			data[36933] <= 8'h10 ;
			data[36934] <= 8'h10 ;
			data[36935] <= 8'h10 ;
			data[36936] <= 8'h10 ;
			data[36937] <= 8'h10 ;
			data[36938] <= 8'h10 ;
			data[36939] <= 8'h10 ;
			data[36940] <= 8'h10 ;
			data[36941] <= 8'h10 ;
			data[36942] <= 8'h10 ;
			data[36943] <= 8'h10 ;
			data[36944] <= 8'h10 ;
			data[36945] <= 8'h10 ;
			data[36946] <= 8'h10 ;
			data[36947] <= 8'h10 ;
			data[36948] <= 8'h10 ;
			data[36949] <= 8'h10 ;
			data[36950] <= 8'h10 ;
			data[36951] <= 8'h10 ;
			data[36952] <= 8'h10 ;
			data[36953] <= 8'h10 ;
			data[36954] <= 8'h10 ;
			data[36955] <= 8'h10 ;
			data[36956] <= 8'h10 ;
			data[36957] <= 8'h10 ;
			data[36958] <= 8'h10 ;
			data[36959] <= 8'h10 ;
			data[36960] <= 8'h10 ;
			data[36961] <= 8'h10 ;
			data[36962] <= 8'h10 ;
			data[36963] <= 8'h10 ;
			data[36964] <= 8'h10 ;
			data[36965] <= 8'h10 ;
			data[36966] <= 8'h10 ;
			data[36967] <= 8'h10 ;
			data[36968] <= 8'h10 ;
			data[36969] <= 8'h10 ;
			data[36970] <= 8'h10 ;
			data[36971] <= 8'h10 ;
			data[36972] <= 8'h10 ;
			data[36973] <= 8'h10 ;
			data[36974] <= 8'h10 ;
			data[36975] <= 8'h10 ;
			data[36976] <= 8'h10 ;
			data[36977] <= 8'h10 ;
			data[36978] <= 8'h10 ;
			data[36979] <= 8'h10 ;
			data[36980] <= 8'h10 ;
			data[36981] <= 8'h10 ;
			data[36982] <= 8'h10 ;
			data[36983] <= 8'h10 ;
			data[36984] <= 8'h10 ;
			data[36985] <= 8'h10 ;
			data[36986] <= 8'h10 ;
			data[36987] <= 8'h10 ;
			data[36988] <= 8'h10 ;
			data[36989] <= 8'h10 ;
			data[36990] <= 8'h10 ;
			data[36991] <= 8'h10 ;
			data[36992] <= 8'h10 ;
			data[36993] <= 8'h10 ;
			data[36994] <= 8'h10 ;
			data[36995] <= 8'h10 ;
			data[36996] <= 8'h10 ;
			data[36997] <= 8'h10 ;
			data[36998] <= 8'h10 ;
			data[36999] <= 8'h10 ;
			data[37000] <= 8'h10 ;
			data[37001] <= 8'h10 ;
			data[37002] <= 8'h10 ;
			data[37003] <= 8'h10 ;
			data[37004] <= 8'h10 ;
			data[37005] <= 8'h10 ;
			data[37006] <= 8'h10 ;
			data[37007] <= 8'h10 ;
			data[37008] <= 8'h10 ;
			data[37009] <= 8'h10 ;
			data[37010] <= 8'h10 ;
			data[37011] <= 8'h10 ;
			data[37012] <= 8'h10 ;
			data[37013] <= 8'h10 ;
			data[37014] <= 8'h10 ;
			data[37015] <= 8'h10 ;
			data[37016] <= 8'h10 ;
			data[37017] <= 8'h10 ;
			data[37018] <= 8'h10 ;
			data[37019] <= 8'h10 ;
			data[37020] <= 8'h10 ;
			data[37021] <= 8'h10 ;
			data[37022] <= 8'h10 ;
			data[37023] <= 8'h10 ;
			data[37024] <= 8'h10 ;
			data[37025] <= 8'h10 ;
			data[37026] <= 8'h10 ;
			data[37027] <= 8'h10 ;
			data[37028] <= 8'h10 ;
			data[37029] <= 8'h10 ;
			data[37030] <= 8'h10 ;
			data[37031] <= 8'h10 ;
			data[37032] <= 8'h10 ;
			data[37033] <= 8'h10 ;
			data[37034] <= 8'h10 ;
			data[37035] <= 8'h10 ;
			data[37036] <= 8'h10 ;
			data[37037] <= 8'h10 ;
			data[37038] <= 8'h10 ;
			data[37039] <= 8'h10 ;
			data[37040] <= 8'h10 ;
			data[37041] <= 8'h10 ;
			data[37042] <= 8'h10 ;
			data[37043] <= 8'h10 ;
			data[37044] <= 8'h10 ;
			data[37045] <= 8'h10 ;
			data[37046] <= 8'h10 ;
			data[37047] <= 8'h10 ;
			data[37048] <= 8'h10 ;
			data[37049] <= 8'h10 ;
			data[37050] <= 8'h10 ;
			data[37051] <= 8'h10 ;
			data[37052] <= 8'h10 ;
			data[37053] <= 8'h10 ;
			data[37054] <= 8'h10 ;
			data[37055] <= 8'h10 ;
			data[37056] <= 8'h10 ;
			data[37057] <= 8'h10 ;
			data[37058] <= 8'h10 ;
			data[37059] <= 8'h10 ;
			data[37060] <= 8'h10 ;
			data[37061] <= 8'h10 ;
			data[37062] <= 8'h10 ;
			data[37063] <= 8'h10 ;
			data[37064] <= 8'h10 ;
			data[37065] <= 8'h10 ;
			data[37066] <= 8'h10 ;
			data[37067] <= 8'h10 ;
			data[37068] <= 8'h10 ;
			data[37069] <= 8'h10 ;
			data[37070] <= 8'h10 ;
			data[37071] <= 8'h10 ;
			data[37072] <= 8'h10 ;
			data[37073] <= 8'h10 ;
			data[37074] <= 8'h10 ;
			data[37075] <= 8'h10 ;
			data[37076] <= 8'h10 ;
			data[37077] <= 8'h10 ;
			data[37078] <= 8'h10 ;
			data[37079] <= 8'h10 ;
			data[37080] <= 8'h10 ;
			data[37081] <= 8'h10 ;
			data[37082] <= 8'h10 ;
			data[37083] <= 8'h10 ;
			data[37084] <= 8'h10 ;
			data[37085] <= 8'h10 ;
			data[37086] <= 8'h10 ;
			data[37087] <= 8'h10 ;
			data[37088] <= 8'h10 ;
			data[37089] <= 8'h10 ;
			data[37090] <= 8'h10 ;
			data[37091] <= 8'h10 ;
			data[37092] <= 8'h10 ;
			data[37093] <= 8'h10 ;
			data[37094] <= 8'h10 ;
			data[37095] <= 8'h10 ;
			data[37096] <= 8'h10 ;
			data[37097] <= 8'h10 ;
			data[37098] <= 8'h10 ;
			data[37099] <= 8'h10 ;
			data[37100] <= 8'h10 ;
			data[37101] <= 8'h10 ;
			data[37102] <= 8'h10 ;
			data[37103] <= 8'h10 ;
			data[37104] <= 8'h10 ;
			data[37105] <= 8'h10 ;
			data[37106] <= 8'h10 ;
			data[37107] <= 8'h10 ;
			data[37108] <= 8'h10 ;
			data[37109] <= 8'h10 ;
			data[37110] <= 8'h10 ;
			data[37111] <= 8'h10 ;
			data[37112] <= 8'h10 ;
			data[37113] <= 8'h10 ;
			data[37114] <= 8'h10 ;
			data[37115] <= 8'h10 ;
			data[37116] <= 8'h10 ;
			data[37117] <= 8'h10 ;
			data[37118] <= 8'h10 ;
			data[37119] <= 8'h10 ;
			data[37120] <= 8'h10 ;
			data[37121] <= 8'h10 ;
			data[37122] <= 8'h10 ;
			data[37123] <= 8'h10 ;
			data[37124] <= 8'h10 ;
			data[37125] <= 8'h10 ;
			data[37126] <= 8'h10 ;
			data[37127] <= 8'h10 ;
			data[37128] <= 8'h10 ;
			data[37129] <= 8'h10 ;
			data[37130] <= 8'h10 ;
			data[37131] <= 8'h10 ;
			data[37132] <= 8'h10 ;
			data[37133] <= 8'h10 ;
			data[37134] <= 8'h10 ;
			data[37135] <= 8'h10 ;
			data[37136] <= 8'h10 ;
			data[37137] <= 8'h10 ;
			data[37138] <= 8'h10 ;
			data[37139] <= 8'h10 ;
			data[37140] <= 8'h10 ;
			data[37141] <= 8'h10 ;
			data[37142] <= 8'h10 ;
			data[37143] <= 8'h10 ;
			data[37144] <= 8'h10 ;
			data[37145] <= 8'h10 ;
			data[37146] <= 8'h10 ;
			data[37147] <= 8'h10 ;
			data[37148] <= 8'h10 ;
			data[37149] <= 8'h10 ;
			data[37150] <= 8'h10 ;
			data[37151] <= 8'h10 ;
			data[37152] <= 8'h10 ;
			data[37153] <= 8'h10 ;
			data[37154] <= 8'h10 ;
			data[37155] <= 8'h10 ;
			data[37156] <= 8'h10 ;
			data[37157] <= 8'h10 ;
			data[37158] <= 8'h10 ;
			data[37159] <= 8'h10 ;
			data[37160] <= 8'h10 ;
			data[37161] <= 8'h10 ;
			data[37162] <= 8'h10 ;
			data[37163] <= 8'h10 ;
			data[37164] <= 8'h10 ;
			data[37165] <= 8'h10 ;
			data[37166] <= 8'h10 ;
			data[37167] <= 8'h10 ;
			data[37168] <= 8'h10 ;
			data[37169] <= 8'h10 ;
			data[37170] <= 8'h10 ;
			data[37171] <= 8'h10 ;
			data[37172] <= 8'h10 ;
			data[37173] <= 8'h10 ;
			data[37174] <= 8'h10 ;
			data[37175] <= 8'h10 ;
			data[37176] <= 8'h10 ;
			data[37177] <= 8'h10 ;
			data[37178] <= 8'h10 ;
			data[37179] <= 8'h10 ;
			data[37180] <= 8'h10 ;
			data[37181] <= 8'h10 ;
			data[37182] <= 8'h10 ;
			data[37183] <= 8'h10 ;
			data[37184] <= 8'h10 ;
			data[37185] <= 8'h10 ;
			data[37186] <= 8'h10 ;
			data[37187] <= 8'h10 ;
			data[37188] <= 8'h10 ;
			data[37189] <= 8'h10 ;
			data[37190] <= 8'h10 ;
			data[37191] <= 8'h10 ;
			data[37192] <= 8'h10 ;
			data[37193] <= 8'h10 ;
			data[37194] <= 8'h10 ;
			data[37195] <= 8'h10 ;
			data[37196] <= 8'h10 ;
			data[37197] <= 8'h10 ;
			data[37198] <= 8'h10 ;
			data[37199] <= 8'h10 ;
			data[37200] <= 8'h10 ;
			data[37201] <= 8'h10 ;
			data[37202] <= 8'h10 ;
			data[37203] <= 8'h10 ;
			data[37204] <= 8'h10 ;
			data[37205] <= 8'h10 ;
			data[37206] <= 8'h10 ;
			data[37207] <= 8'h10 ;
			data[37208] <= 8'h10 ;
			data[37209] <= 8'h10 ;
			data[37210] <= 8'h10 ;
			data[37211] <= 8'h10 ;
			data[37212] <= 8'h10 ;
			data[37213] <= 8'h10 ;
			data[37214] <= 8'h10 ;
			data[37215] <= 8'h10 ;
			data[37216] <= 8'h10 ;
			data[37217] <= 8'h10 ;
			data[37218] <= 8'h10 ;
			data[37219] <= 8'h10 ;
			data[37220] <= 8'h10 ;
			data[37221] <= 8'h10 ;
			data[37222] <= 8'h10 ;
			data[37223] <= 8'h10 ;
			data[37224] <= 8'h10 ;
			data[37225] <= 8'h10 ;
			data[37226] <= 8'h10 ;
			data[37227] <= 8'h10 ;
			data[37228] <= 8'h10 ;
			data[37229] <= 8'h10 ;
			data[37230] <= 8'h10 ;
			data[37231] <= 8'h10 ;
			data[37232] <= 8'h10 ;
			data[37233] <= 8'h10 ;
			data[37234] <= 8'h10 ;
			data[37235] <= 8'h10 ;
			data[37236] <= 8'h10 ;
			data[37237] <= 8'h10 ;
			data[37238] <= 8'h10 ;
			data[37239] <= 8'h10 ;
			data[37240] <= 8'h10 ;
			data[37241] <= 8'h10 ;
			data[37242] <= 8'h10 ;
			data[37243] <= 8'h10 ;
			data[37244] <= 8'h10 ;
			data[37245] <= 8'h10 ;
			data[37246] <= 8'h10 ;
			data[37247] <= 8'h10 ;
			data[37248] <= 8'h10 ;
			data[37249] <= 8'h10 ;
			data[37250] <= 8'h10 ;
			data[37251] <= 8'h10 ;
			data[37252] <= 8'h10 ;
			data[37253] <= 8'h10 ;
			data[37254] <= 8'h10 ;
			data[37255] <= 8'h10 ;
			data[37256] <= 8'h10 ;
			data[37257] <= 8'h10 ;
			data[37258] <= 8'h10 ;
			data[37259] <= 8'h10 ;
			data[37260] <= 8'h10 ;
			data[37261] <= 8'h10 ;
			data[37262] <= 8'h10 ;
			data[37263] <= 8'h10 ;
			data[37264] <= 8'h10 ;
			data[37265] <= 8'h10 ;
			data[37266] <= 8'h10 ;
			data[37267] <= 8'h10 ;
			data[37268] <= 8'h10 ;
			data[37269] <= 8'h10 ;
			data[37270] <= 8'h10 ;
			data[37271] <= 8'h10 ;
			data[37272] <= 8'h10 ;
			data[37273] <= 8'h10 ;
			data[37274] <= 8'h10 ;
			data[37275] <= 8'h10 ;
			data[37276] <= 8'h10 ;
			data[37277] <= 8'h10 ;
			data[37278] <= 8'h10 ;
			data[37279] <= 8'h10 ;
			data[37280] <= 8'h10 ;
			data[37281] <= 8'h10 ;
			data[37282] <= 8'h10 ;
			data[37283] <= 8'h10 ;
			data[37284] <= 8'h10 ;
			data[37285] <= 8'h10 ;
			data[37286] <= 8'h10 ;
			data[37287] <= 8'h10 ;
			data[37288] <= 8'h10 ;
			data[37289] <= 8'h10 ;
			data[37290] <= 8'h10 ;
			data[37291] <= 8'h10 ;
			data[37292] <= 8'h10 ;
			data[37293] <= 8'h10 ;
			data[37294] <= 8'h10 ;
			data[37295] <= 8'h10 ;
			data[37296] <= 8'h10 ;
			data[37297] <= 8'h10 ;
			data[37298] <= 8'h10 ;
			data[37299] <= 8'h10 ;
			data[37300] <= 8'h10 ;
			data[37301] <= 8'h10 ;
			data[37302] <= 8'h10 ;
			data[37303] <= 8'h10 ;
			data[37304] <= 8'h10 ;
			data[37305] <= 8'h10 ;
			data[37306] <= 8'h10 ;
			data[37307] <= 8'h10 ;
			data[37308] <= 8'h10 ;
			data[37309] <= 8'h10 ;
			data[37310] <= 8'h10 ;
			data[37311] <= 8'h10 ;
			data[37312] <= 8'h10 ;
			data[37313] <= 8'h10 ;
			data[37314] <= 8'h10 ;
			data[37315] <= 8'h10 ;
			data[37316] <= 8'h10 ;
			data[37317] <= 8'h10 ;
			data[37318] <= 8'h10 ;
			data[37319] <= 8'h10 ;
			data[37320] <= 8'h10 ;
			data[37321] <= 8'h10 ;
			data[37322] <= 8'h10 ;
			data[37323] <= 8'h10 ;
			data[37324] <= 8'h10 ;
			data[37325] <= 8'h10 ;
			data[37326] <= 8'h10 ;
			data[37327] <= 8'h10 ;
			data[37328] <= 8'h10 ;
			data[37329] <= 8'h10 ;
			data[37330] <= 8'h10 ;
			data[37331] <= 8'h10 ;
			data[37332] <= 8'h10 ;
			data[37333] <= 8'h10 ;
			data[37334] <= 8'h10 ;
			data[37335] <= 8'h10 ;
			data[37336] <= 8'h10 ;
			data[37337] <= 8'h10 ;
			data[37338] <= 8'h10 ;
			data[37339] <= 8'h10 ;
			data[37340] <= 8'h10 ;
			data[37341] <= 8'h10 ;
			data[37342] <= 8'h10 ;
			data[37343] <= 8'h10 ;
			data[37344] <= 8'h10 ;
			data[37345] <= 8'h10 ;
			data[37346] <= 8'h10 ;
			data[37347] <= 8'h10 ;
			data[37348] <= 8'h10 ;
			data[37349] <= 8'h10 ;
			data[37350] <= 8'h10 ;
			data[37351] <= 8'h10 ;
			data[37352] <= 8'h10 ;
			data[37353] <= 8'h10 ;
			data[37354] <= 8'h10 ;
			data[37355] <= 8'h10 ;
			data[37356] <= 8'h10 ;
			data[37357] <= 8'h10 ;
			data[37358] <= 8'h10 ;
			data[37359] <= 8'h10 ;
			data[37360] <= 8'h10 ;
			data[37361] <= 8'h10 ;
			data[37362] <= 8'h10 ;
			data[37363] <= 8'h10 ;
			data[37364] <= 8'h10 ;
			data[37365] <= 8'h10 ;
			data[37366] <= 8'h10 ;
			data[37367] <= 8'h10 ;
			data[37368] <= 8'h10 ;
			data[37369] <= 8'h10 ;
			data[37370] <= 8'h10 ;
			data[37371] <= 8'h10 ;
			data[37372] <= 8'h10 ;
			data[37373] <= 8'h10 ;
			data[37374] <= 8'h10 ;
			data[37375] <= 8'h10 ;
			data[37376] <= 8'h10 ;
			data[37377] <= 8'h10 ;
			data[37378] <= 8'h10 ;
			data[37379] <= 8'h10 ;
			data[37380] <= 8'h10 ;
			data[37381] <= 8'h10 ;
			data[37382] <= 8'h10 ;
			data[37383] <= 8'h10 ;
			data[37384] <= 8'h10 ;
			data[37385] <= 8'h10 ;
			data[37386] <= 8'h10 ;
			data[37387] <= 8'h10 ;
			data[37388] <= 8'h10 ;
			data[37389] <= 8'h10 ;
			data[37390] <= 8'h10 ;
			data[37391] <= 8'h10 ;
			data[37392] <= 8'h10 ;
			data[37393] <= 8'h10 ;
			data[37394] <= 8'h10 ;
			data[37395] <= 8'h10 ;
			data[37396] <= 8'h10 ;
			data[37397] <= 8'h10 ;
			data[37398] <= 8'h10 ;
			data[37399] <= 8'h10 ;
			data[37400] <= 8'h10 ;
			data[37401] <= 8'h10 ;
			data[37402] <= 8'h10 ;
			data[37403] <= 8'h10 ;
			data[37404] <= 8'h10 ;
			data[37405] <= 8'h10 ;
			data[37406] <= 8'h10 ;
			data[37407] <= 8'h10 ;
			data[37408] <= 8'h10 ;
			data[37409] <= 8'h10 ;
			data[37410] <= 8'h10 ;
			data[37411] <= 8'h10 ;
			data[37412] <= 8'h10 ;
			data[37413] <= 8'h10 ;
			data[37414] <= 8'h10 ;
			data[37415] <= 8'h10 ;
			data[37416] <= 8'h10 ;
			data[37417] <= 8'h10 ;
			data[37418] <= 8'h10 ;
			data[37419] <= 8'h10 ;
			data[37420] <= 8'h10 ;
			data[37421] <= 8'h10 ;
			data[37422] <= 8'h10 ;
			data[37423] <= 8'h10 ;
			data[37424] <= 8'h10 ;
			data[37425] <= 8'h10 ;
			data[37426] <= 8'h10 ;
			data[37427] <= 8'h10 ;
			data[37428] <= 8'h10 ;
			data[37429] <= 8'h10 ;
			data[37430] <= 8'h10 ;
			data[37431] <= 8'h10 ;
			data[37432] <= 8'h10 ;
			data[37433] <= 8'h10 ;
			data[37434] <= 8'h10 ;
			data[37435] <= 8'h10 ;
			data[37436] <= 8'h10 ;
			data[37437] <= 8'h10 ;
			data[37438] <= 8'h10 ;
			data[37439] <= 8'h10 ;
			data[37440] <= 8'h10 ;
			data[37441] <= 8'h10 ;
			data[37442] <= 8'h10 ;
			data[37443] <= 8'h10 ;
			data[37444] <= 8'h10 ;
			data[37445] <= 8'h10 ;
			data[37446] <= 8'h10 ;
			data[37447] <= 8'h10 ;
			data[37448] <= 8'h10 ;
			data[37449] <= 8'h10 ;
			data[37450] <= 8'h10 ;
			data[37451] <= 8'h10 ;
			data[37452] <= 8'h10 ;
			data[37453] <= 8'h10 ;
			data[37454] <= 8'h10 ;
			data[37455] <= 8'h10 ;
			data[37456] <= 8'h10 ;
			data[37457] <= 8'h10 ;
			data[37458] <= 8'h10 ;
			data[37459] <= 8'h10 ;
			data[37460] <= 8'h10 ;
			data[37461] <= 8'h10 ;
			data[37462] <= 8'h10 ;
			data[37463] <= 8'h10 ;
			data[37464] <= 8'h10 ;
			data[37465] <= 8'h10 ;
			data[37466] <= 8'h10 ;
			data[37467] <= 8'h10 ;
			data[37468] <= 8'h10 ;
			data[37469] <= 8'h10 ;
			data[37470] <= 8'h10 ;
			data[37471] <= 8'h10 ;
			data[37472] <= 8'h10 ;
			data[37473] <= 8'h10 ;
			data[37474] <= 8'h10 ;
			data[37475] <= 8'h10 ;
			data[37476] <= 8'h10 ;
			data[37477] <= 8'h10 ;
			data[37478] <= 8'h10 ;
			data[37479] <= 8'h10 ;
			data[37480] <= 8'h10 ;
			data[37481] <= 8'h10 ;
			data[37482] <= 8'h10 ;
			data[37483] <= 8'h10 ;
			data[37484] <= 8'h10 ;
			data[37485] <= 8'h10 ;
			data[37486] <= 8'h10 ;
			data[37487] <= 8'h10 ;
			data[37488] <= 8'h10 ;
			data[37489] <= 8'h10 ;
			data[37490] <= 8'h10 ;
			data[37491] <= 8'h10 ;
			data[37492] <= 8'h10 ;
			data[37493] <= 8'h10 ;
			data[37494] <= 8'h10 ;
			data[37495] <= 8'h10 ;
			data[37496] <= 8'h10 ;
			data[37497] <= 8'h10 ;
			data[37498] <= 8'h10 ;
			data[37499] <= 8'h10 ;
			data[37500] <= 8'h10 ;
			data[37501] <= 8'h10 ;
			data[37502] <= 8'h10 ;
			data[37503] <= 8'h10 ;
			data[37504] <= 8'h10 ;
			data[37505] <= 8'h10 ;
			data[37506] <= 8'h10 ;
			data[37507] <= 8'h10 ;
			data[37508] <= 8'h10 ;
			data[37509] <= 8'h10 ;
			data[37510] <= 8'h10 ;
			data[37511] <= 8'h10 ;
			data[37512] <= 8'h10 ;
			data[37513] <= 8'h10 ;
			data[37514] <= 8'h10 ;
			data[37515] <= 8'h10 ;
			data[37516] <= 8'h10 ;
			data[37517] <= 8'h10 ;
			data[37518] <= 8'h10 ;
			data[37519] <= 8'h10 ;
			data[37520] <= 8'h10 ;
			data[37521] <= 8'h10 ;
			data[37522] <= 8'h10 ;
			data[37523] <= 8'h10 ;
			data[37524] <= 8'h10 ;
			data[37525] <= 8'h10 ;
			data[37526] <= 8'h10 ;
			data[37527] <= 8'h10 ;
			data[37528] <= 8'h10 ;
			data[37529] <= 8'h10 ;
			data[37530] <= 8'h10 ;
			data[37531] <= 8'h10 ;
			data[37532] <= 8'h10 ;
			data[37533] <= 8'h10 ;
			data[37534] <= 8'h10 ;
			data[37535] <= 8'h10 ;
			data[37536] <= 8'h10 ;
			data[37537] <= 8'h10 ;
			data[37538] <= 8'h10 ;
			data[37539] <= 8'h10 ;
			data[37540] <= 8'h10 ;
			data[37541] <= 8'h10 ;
			data[37542] <= 8'h10 ;
			data[37543] <= 8'h10 ;
			data[37544] <= 8'h10 ;
			data[37545] <= 8'h10 ;
			data[37546] <= 8'h10 ;
			data[37547] <= 8'h10 ;
			data[37548] <= 8'h10 ;
			data[37549] <= 8'h10 ;
			data[37550] <= 8'h10 ;
			data[37551] <= 8'h10 ;
			data[37552] <= 8'h10 ;
			data[37553] <= 8'h10 ;
			data[37554] <= 8'h10 ;
			data[37555] <= 8'h10 ;
			data[37556] <= 8'h10 ;
			data[37557] <= 8'h10 ;
			data[37558] <= 8'h10 ;
			data[37559] <= 8'h10 ;
			data[37560] <= 8'h10 ;
			data[37561] <= 8'h10 ;
			data[37562] <= 8'h10 ;
			data[37563] <= 8'h10 ;
			data[37564] <= 8'h10 ;
			data[37565] <= 8'h10 ;
			data[37566] <= 8'h10 ;
			data[37567] <= 8'h10 ;
			data[37568] <= 8'h10 ;
			data[37569] <= 8'h10 ;
			data[37570] <= 8'h10 ;
			data[37571] <= 8'h10 ;
			data[37572] <= 8'h10 ;
			data[37573] <= 8'h10 ;
			data[37574] <= 8'h10 ;
			data[37575] <= 8'h10 ;
			data[37576] <= 8'h10 ;
			data[37577] <= 8'h10 ;
			data[37578] <= 8'h10 ;
			data[37579] <= 8'h10 ;
			data[37580] <= 8'h10 ;
			data[37581] <= 8'h10 ;
			data[37582] <= 8'h10 ;
			data[37583] <= 8'h10 ;
			data[37584] <= 8'h10 ;
			data[37585] <= 8'h10 ;
			data[37586] <= 8'h10 ;
			data[37587] <= 8'h10 ;
			data[37588] <= 8'h10 ;
			data[37589] <= 8'h10 ;
			data[37590] <= 8'h10 ;
			data[37591] <= 8'h10 ;
			data[37592] <= 8'h10 ;
			data[37593] <= 8'h10 ;
			data[37594] <= 8'h10 ;
			data[37595] <= 8'h10 ;
			data[37596] <= 8'h10 ;
			data[37597] <= 8'h10 ;
			data[37598] <= 8'h10 ;
			data[37599] <= 8'h10 ;
			data[37600] <= 8'h10 ;
			data[37601] <= 8'h10 ;
			data[37602] <= 8'h10 ;
			data[37603] <= 8'h10 ;
			data[37604] <= 8'h10 ;
			data[37605] <= 8'h10 ;
			data[37606] <= 8'h10 ;
			data[37607] <= 8'h10 ;
			data[37608] <= 8'h10 ;
			data[37609] <= 8'h10 ;
			data[37610] <= 8'h10 ;
			data[37611] <= 8'h10 ;
			data[37612] <= 8'h10 ;
			data[37613] <= 8'h10 ;
			data[37614] <= 8'h10 ;
			data[37615] <= 8'h10 ;
			data[37616] <= 8'h10 ;
			data[37617] <= 8'h10 ;
			data[37618] <= 8'h10 ;
			data[37619] <= 8'h10 ;
			data[37620] <= 8'h10 ;
			data[37621] <= 8'h10 ;
			data[37622] <= 8'h10 ;
			data[37623] <= 8'h10 ;
			data[37624] <= 8'h10 ;
			data[37625] <= 8'h10 ;
			data[37626] <= 8'h10 ;
			data[37627] <= 8'h10 ;
			data[37628] <= 8'h10 ;
			data[37629] <= 8'h10 ;
			data[37630] <= 8'h10 ;
			data[37631] <= 8'h10 ;
			data[37632] <= 8'h10 ;
			data[37633] <= 8'h10 ;
			data[37634] <= 8'h10 ;
			data[37635] <= 8'h10 ;
			data[37636] <= 8'h10 ;
			data[37637] <= 8'h10 ;
			data[37638] <= 8'h10 ;
			data[37639] <= 8'h10 ;
			data[37640] <= 8'h10 ;
			data[37641] <= 8'h10 ;
			data[37642] <= 8'h10 ;
			data[37643] <= 8'h10 ;
			data[37644] <= 8'h10 ;
			data[37645] <= 8'h10 ;
			data[37646] <= 8'h10 ;
			data[37647] <= 8'h10 ;
			data[37648] <= 8'h10 ;
			data[37649] <= 8'h10 ;
			data[37650] <= 8'h10 ;
			data[37651] <= 8'h10 ;
			data[37652] <= 8'h10 ;
			data[37653] <= 8'h10 ;
			data[37654] <= 8'h10 ;
			data[37655] <= 8'h10 ;
			data[37656] <= 8'h10 ;
			data[37657] <= 8'h10 ;
			data[37658] <= 8'h10 ;
			data[37659] <= 8'h10 ;
			data[37660] <= 8'h10 ;
			data[37661] <= 8'h10 ;
			data[37662] <= 8'h10 ;
			data[37663] <= 8'h10 ;
			data[37664] <= 8'h10 ;
			data[37665] <= 8'h10 ;
			data[37666] <= 8'h10 ;
			data[37667] <= 8'h10 ;
			data[37668] <= 8'h10 ;
			data[37669] <= 8'h10 ;
			data[37670] <= 8'h10 ;
			data[37671] <= 8'h10 ;
			data[37672] <= 8'h10 ;
			data[37673] <= 8'h10 ;
			data[37674] <= 8'h10 ;
			data[37675] <= 8'h10 ;
			data[37676] <= 8'h10 ;
			data[37677] <= 8'h10 ;
			data[37678] <= 8'h10 ;
			data[37679] <= 8'h10 ;
			data[37680] <= 8'h10 ;
			data[37681] <= 8'h10 ;
			data[37682] <= 8'h10 ;
			data[37683] <= 8'h10 ;
			data[37684] <= 8'h10 ;
			data[37685] <= 8'h10 ;
			data[37686] <= 8'h10 ;
			data[37687] <= 8'h10 ;
			data[37688] <= 8'h10 ;
			data[37689] <= 8'h10 ;
			data[37690] <= 8'h10 ;
			data[37691] <= 8'h10 ;
			data[37692] <= 8'h10 ;
			data[37693] <= 8'h10 ;
			data[37694] <= 8'h10 ;
			data[37695] <= 8'h10 ;
			data[37696] <= 8'h10 ;
			data[37697] <= 8'h10 ;
			data[37698] <= 8'h10 ;
			data[37699] <= 8'h10 ;
			data[37700] <= 8'h10 ;
			data[37701] <= 8'h10 ;
			data[37702] <= 8'h10 ;
			data[37703] <= 8'h10 ;
			data[37704] <= 8'h10 ;
			data[37705] <= 8'h10 ;
			data[37706] <= 8'h10 ;
			data[37707] <= 8'h10 ;
			data[37708] <= 8'h10 ;
			data[37709] <= 8'h10 ;
			data[37710] <= 8'h10 ;
			data[37711] <= 8'h10 ;
			data[37712] <= 8'h10 ;
			data[37713] <= 8'h10 ;
			data[37714] <= 8'h10 ;
			data[37715] <= 8'h10 ;
			data[37716] <= 8'h10 ;
			data[37717] <= 8'h10 ;
			data[37718] <= 8'h10 ;
			data[37719] <= 8'h10 ;
			data[37720] <= 8'h10 ;
			data[37721] <= 8'h10 ;
			data[37722] <= 8'h10 ;
			data[37723] <= 8'h10 ;
			data[37724] <= 8'h10 ;
			data[37725] <= 8'h10 ;
			data[37726] <= 8'h10 ;
			data[37727] <= 8'h10 ;
			data[37728] <= 8'h10 ;
			data[37729] <= 8'h10 ;
			data[37730] <= 8'h10 ;
			data[37731] <= 8'h10 ;
			data[37732] <= 8'h10 ;
			data[37733] <= 8'h10 ;
			data[37734] <= 8'h10 ;
			data[37735] <= 8'h10 ;
			data[37736] <= 8'h10 ;
			data[37737] <= 8'h10 ;
			data[37738] <= 8'h10 ;
			data[37739] <= 8'h10 ;
			data[37740] <= 8'h10 ;
			data[37741] <= 8'h10 ;
			data[37742] <= 8'h10 ;
			data[37743] <= 8'h10 ;
			data[37744] <= 8'h10 ;
			data[37745] <= 8'h10 ;
			data[37746] <= 8'h10 ;
			data[37747] <= 8'h10 ;
			data[37748] <= 8'h10 ;
			data[37749] <= 8'h10 ;
			data[37750] <= 8'h10 ;
			data[37751] <= 8'h10 ;
			data[37752] <= 8'h10 ;
			data[37753] <= 8'h10 ;
			data[37754] <= 8'h10 ;
			data[37755] <= 8'h10 ;
			data[37756] <= 8'h10 ;
			data[37757] <= 8'h10 ;
			data[37758] <= 8'h10 ;
			data[37759] <= 8'h10 ;
			data[37760] <= 8'h10 ;
			data[37761] <= 8'h10 ;
			data[37762] <= 8'h10 ;
			data[37763] <= 8'h10 ;
			data[37764] <= 8'h10 ;
			data[37765] <= 8'h10 ;
			data[37766] <= 8'h10 ;
			data[37767] <= 8'h10 ;
			data[37768] <= 8'h10 ;
			data[37769] <= 8'h10 ;
			data[37770] <= 8'h10 ;
			data[37771] <= 8'h10 ;
			data[37772] <= 8'h10 ;
			data[37773] <= 8'h10 ;
			data[37774] <= 8'h10 ;
			data[37775] <= 8'h10 ;
			data[37776] <= 8'h10 ;
			data[37777] <= 8'h10 ;
			data[37778] <= 8'h10 ;
			data[37779] <= 8'h10 ;
			data[37780] <= 8'h10 ;
			data[37781] <= 8'h10 ;
			data[37782] <= 8'h10 ;
			data[37783] <= 8'h10 ;
			data[37784] <= 8'h10 ;
			data[37785] <= 8'h10 ;
			data[37786] <= 8'h10 ;
			data[37787] <= 8'h10 ;
			data[37788] <= 8'h10 ;
			data[37789] <= 8'h10 ;
			data[37790] <= 8'h10 ;
			data[37791] <= 8'h10 ;
			data[37792] <= 8'h10 ;
			data[37793] <= 8'h10 ;
			data[37794] <= 8'h10 ;
			data[37795] <= 8'h10 ;
			data[37796] <= 8'h10 ;
			data[37797] <= 8'h10 ;
			data[37798] <= 8'h10 ;
			data[37799] <= 8'h10 ;
			data[37800] <= 8'h10 ;
			data[37801] <= 8'h10 ;
			data[37802] <= 8'h10 ;
			data[37803] <= 8'h10 ;
			data[37804] <= 8'h10 ;
			data[37805] <= 8'h10 ;
			data[37806] <= 8'h10 ;
			data[37807] <= 8'h10 ;
			data[37808] <= 8'h10 ;
			data[37809] <= 8'h10 ;
			data[37810] <= 8'h10 ;
			data[37811] <= 8'h10 ;
			data[37812] <= 8'h10 ;
			data[37813] <= 8'h10 ;
			data[37814] <= 8'h10 ;
			data[37815] <= 8'h10 ;
			data[37816] <= 8'h10 ;
			data[37817] <= 8'h10 ;
			data[37818] <= 8'h10 ;
			data[37819] <= 8'h10 ;
			data[37820] <= 8'h10 ;
			data[37821] <= 8'h10 ;
			data[37822] <= 8'h10 ;
			data[37823] <= 8'h10 ;
			data[37824] <= 8'h10 ;
			data[37825] <= 8'h10 ;
			data[37826] <= 8'h10 ;
			data[37827] <= 8'h10 ;
			data[37828] <= 8'h10 ;
			data[37829] <= 8'h10 ;
			data[37830] <= 8'h10 ;
			data[37831] <= 8'h10 ;
			data[37832] <= 8'h10 ;
			data[37833] <= 8'h10 ;
			data[37834] <= 8'h10 ;
			data[37835] <= 8'h10 ;
			data[37836] <= 8'h10 ;
			data[37837] <= 8'h10 ;
			data[37838] <= 8'h10 ;
			data[37839] <= 8'h10 ;
			data[37840] <= 8'h10 ;
			data[37841] <= 8'h10 ;
			data[37842] <= 8'h10 ;
			data[37843] <= 8'h10 ;
			data[37844] <= 8'h10 ;
			data[37845] <= 8'h10 ;
			data[37846] <= 8'h10 ;
			data[37847] <= 8'h10 ;
			data[37848] <= 8'h10 ;
			data[37849] <= 8'h10 ;
			data[37850] <= 8'h10 ;
			data[37851] <= 8'h10 ;
			data[37852] <= 8'h10 ;
			data[37853] <= 8'h10 ;
			data[37854] <= 8'h10 ;
			data[37855] <= 8'h10 ;
			data[37856] <= 8'h10 ;
			data[37857] <= 8'h10 ;
			data[37858] <= 8'h10 ;
			data[37859] <= 8'h10 ;
			data[37860] <= 8'h10 ;
			data[37861] <= 8'h10 ;
			data[37862] <= 8'h10 ;
			data[37863] <= 8'h10 ;
			data[37864] <= 8'h10 ;
			data[37865] <= 8'h10 ;
			data[37866] <= 8'h10 ;
			data[37867] <= 8'h10 ;
			data[37868] <= 8'h10 ;
			data[37869] <= 8'h10 ;
			data[37870] <= 8'h10 ;
			data[37871] <= 8'h10 ;
			data[37872] <= 8'h10 ;
			data[37873] <= 8'h10 ;
			data[37874] <= 8'h10 ;
			data[37875] <= 8'h10 ;
			data[37876] <= 8'h10 ;
			data[37877] <= 8'h10 ;
			data[37878] <= 8'h10 ;
			data[37879] <= 8'h10 ;
			data[37880] <= 8'h10 ;
			data[37881] <= 8'h10 ;
			data[37882] <= 8'h10 ;
			data[37883] <= 8'h10 ;
			data[37884] <= 8'h10 ;
			data[37885] <= 8'h10 ;
			data[37886] <= 8'h10 ;
			data[37887] <= 8'h10 ;
			data[37888] <= 8'h10 ;
			data[37889] <= 8'h10 ;
			data[37890] <= 8'h10 ;
			data[37891] <= 8'h10 ;
			data[37892] <= 8'h10 ;
			data[37893] <= 8'h10 ;
			data[37894] <= 8'h10 ;
			data[37895] <= 8'h10 ;
			data[37896] <= 8'h10 ;
			data[37897] <= 8'h10 ;
			data[37898] <= 8'h10 ;
			data[37899] <= 8'h10 ;
			data[37900] <= 8'h10 ;
			data[37901] <= 8'h10 ;
			data[37902] <= 8'h10 ;
			data[37903] <= 8'h10 ;
			data[37904] <= 8'h10 ;
			data[37905] <= 8'h10 ;
			data[37906] <= 8'h10 ;
			data[37907] <= 8'h10 ;
			data[37908] <= 8'h10 ;
			data[37909] <= 8'h10 ;
			data[37910] <= 8'h10 ;
			data[37911] <= 8'h10 ;
			data[37912] <= 8'h10 ;
			data[37913] <= 8'h10 ;
			data[37914] <= 8'h10 ;
			data[37915] <= 8'h10 ;
			data[37916] <= 8'h10 ;
			data[37917] <= 8'h10 ;
			data[37918] <= 8'h10 ;
			data[37919] <= 8'h10 ;
			data[37920] <= 8'h10 ;
			data[37921] <= 8'h10 ;
			data[37922] <= 8'h10 ;
			data[37923] <= 8'h10 ;
			data[37924] <= 8'h10 ;
			data[37925] <= 8'h10 ;
			data[37926] <= 8'h10 ;
			data[37927] <= 8'h10 ;
			data[37928] <= 8'h10 ;
			data[37929] <= 8'h10 ;
			data[37930] <= 8'h10 ;
			data[37931] <= 8'h10 ;
			data[37932] <= 8'h10 ;
			data[37933] <= 8'h10 ;
			data[37934] <= 8'h10 ;
			data[37935] <= 8'h10 ;
			data[37936] <= 8'h10 ;
			data[37937] <= 8'h10 ;
			data[37938] <= 8'h10 ;
			data[37939] <= 8'h10 ;
			data[37940] <= 8'h10 ;
			data[37941] <= 8'h10 ;
			data[37942] <= 8'h10 ;
			data[37943] <= 8'h10 ;
			data[37944] <= 8'h10 ;
			data[37945] <= 8'h10 ;
			data[37946] <= 8'h10 ;
			data[37947] <= 8'h10 ;
			data[37948] <= 8'h10 ;
			data[37949] <= 8'h10 ;
			data[37950] <= 8'h10 ;
			data[37951] <= 8'h10 ;
			data[37952] <= 8'h10 ;
			data[37953] <= 8'h10 ;
			data[37954] <= 8'h10 ;
			data[37955] <= 8'h10 ;
			data[37956] <= 8'h10 ;
			data[37957] <= 8'h10 ;
			data[37958] <= 8'h10 ;
			data[37959] <= 8'h10 ;
			data[37960] <= 8'h10 ;
			data[37961] <= 8'h10 ;
			data[37962] <= 8'h10 ;
			data[37963] <= 8'h10 ;
			data[37964] <= 8'h10 ;
			data[37965] <= 8'h10 ;
			data[37966] <= 8'h10 ;
			data[37967] <= 8'h10 ;
			data[37968] <= 8'h10 ;
			data[37969] <= 8'h10 ;
			data[37970] <= 8'h10 ;
			data[37971] <= 8'h10 ;
			data[37972] <= 8'h10 ;
			data[37973] <= 8'h10 ;
			data[37974] <= 8'h10 ;
			data[37975] <= 8'h10 ;
			data[37976] <= 8'h10 ;
			data[37977] <= 8'h10 ;
			data[37978] <= 8'h10 ;
			data[37979] <= 8'h10 ;
			data[37980] <= 8'h10 ;
			data[37981] <= 8'h10 ;
			data[37982] <= 8'h10 ;
			data[37983] <= 8'h10 ;
			data[37984] <= 8'h10 ;
			data[37985] <= 8'h10 ;
			data[37986] <= 8'h10 ;
			data[37987] <= 8'h10 ;
			data[37988] <= 8'h10 ;
			data[37989] <= 8'h10 ;
			data[37990] <= 8'h10 ;
			data[37991] <= 8'h10 ;
			data[37992] <= 8'h10 ;
			data[37993] <= 8'h10 ;
			data[37994] <= 8'h10 ;
			data[37995] <= 8'h10 ;
			data[37996] <= 8'h10 ;
			data[37997] <= 8'h10 ;
			data[37998] <= 8'h10 ;
			data[37999] <= 8'h10 ;
			data[38000] <= 8'h10 ;
			data[38001] <= 8'h10 ;
			data[38002] <= 8'h10 ;
			data[38003] <= 8'h10 ;
			data[38004] <= 8'h10 ;
			data[38005] <= 8'h10 ;
			data[38006] <= 8'h10 ;
			data[38007] <= 8'h10 ;
			data[38008] <= 8'h10 ;
			data[38009] <= 8'h10 ;
			data[38010] <= 8'h10 ;
			data[38011] <= 8'h10 ;
			data[38012] <= 8'h10 ;
			data[38013] <= 8'h10 ;
			data[38014] <= 8'h10 ;
			data[38015] <= 8'h10 ;
			data[38016] <= 8'h10 ;
			data[38017] <= 8'h10 ;
			data[38018] <= 8'h10 ;
			data[38019] <= 8'h10 ;
			data[38020] <= 8'h10 ;
			data[38021] <= 8'h10 ;
			data[38022] <= 8'h10 ;
			data[38023] <= 8'h10 ;
			data[38024] <= 8'h10 ;
			data[38025] <= 8'h10 ;
			data[38026] <= 8'h10 ;
			data[38027] <= 8'h10 ;
			data[38028] <= 8'h10 ;
			data[38029] <= 8'h10 ;
			data[38030] <= 8'h10 ;
			data[38031] <= 8'h10 ;
			data[38032] <= 8'h10 ;
			data[38033] <= 8'h10 ;
			data[38034] <= 8'h10 ;
			data[38035] <= 8'h10 ;
			data[38036] <= 8'h10 ;
			data[38037] <= 8'h10 ;
			data[38038] <= 8'h10 ;
			data[38039] <= 8'h10 ;
			data[38040] <= 8'h10 ;
			data[38041] <= 8'h10 ;
			data[38042] <= 8'h10 ;
			data[38043] <= 8'h10 ;
			data[38044] <= 8'h10 ;
			data[38045] <= 8'h10 ;
			data[38046] <= 8'h10 ;
			data[38047] <= 8'h10 ;
			data[38048] <= 8'h10 ;
			data[38049] <= 8'h10 ;
			data[38050] <= 8'h10 ;
			data[38051] <= 8'h10 ;
			data[38052] <= 8'h10 ;
			data[38053] <= 8'h10 ;
			data[38054] <= 8'h10 ;
			data[38055] <= 8'h10 ;
			data[38056] <= 8'h10 ;
			data[38057] <= 8'h10 ;
			data[38058] <= 8'h10 ;
			data[38059] <= 8'h10 ;
			data[38060] <= 8'h10 ;
			data[38061] <= 8'h10 ;
			data[38062] <= 8'h10 ;
			data[38063] <= 8'h10 ;
			data[38064] <= 8'h10 ;
			data[38065] <= 8'h10 ;
			data[38066] <= 8'h10 ;
			data[38067] <= 8'h10 ;
			data[38068] <= 8'h10 ;
			data[38069] <= 8'h10 ;
			data[38070] <= 8'h10 ;
			data[38071] <= 8'h10 ;
			data[38072] <= 8'h10 ;
			data[38073] <= 8'h10 ;
			data[38074] <= 8'h10 ;
			data[38075] <= 8'h10 ;
			data[38076] <= 8'h10 ;
			data[38077] <= 8'h10 ;
			data[38078] <= 8'h10 ;
			data[38079] <= 8'h10 ;
			data[38080] <= 8'h10 ;
			data[38081] <= 8'h10 ;
			data[38082] <= 8'h10 ;
			data[38083] <= 8'h10 ;
			data[38084] <= 8'h10 ;
			data[38085] <= 8'h10 ;
			data[38086] <= 8'h10 ;
			data[38087] <= 8'h10 ;
			data[38088] <= 8'h10 ;
			data[38089] <= 8'h10 ;
			data[38090] <= 8'h10 ;
			data[38091] <= 8'h10 ;
			data[38092] <= 8'h10 ;
			data[38093] <= 8'h10 ;
			data[38094] <= 8'h10 ;
			data[38095] <= 8'h10 ;
			data[38096] <= 8'h10 ;
			data[38097] <= 8'h10 ;
			data[38098] <= 8'h10 ;
			data[38099] <= 8'h10 ;
			data[38100] <= 8'h10 ;
			data[38101] <= 8'h10 ;
			data[38102] <= 8'h10 ;
			data[38103] <= 8'h10 ;
			data[38104] <= 8'h10 ;
			data[38105] <= 8'h10 ;
			data[38106] <= 8'h10 ;
			data[38107] <= 8'h10 ;
			data[38108] <= 8'h10 ;
			data[38109] <= 8'h10 ;
			data[38110] <= 8'h10 ;
			data[38111] <= 8'h10 ;
			data[38112] <= 8'h10 ;
			data[38113] <= 8'h10 ;
			data[38114] <= 8'h10 ;
			data[38115] <= 8'h10 ;
			data[38116] <= 8'h10 ;
			data[38117] <= 8'h10 ;
			data[38118] <= 8'h10 ;
			data[38119] <= 8'h10 ;
			data[38120] <= 8'h10 ;
			data[38121] <= 8'h10 ;
			data[38122] <= 8'h10 ;
			data[38123] <= 8'h10 ;
			data[38124] <= 8'h10 ;
			data[38125] <= 8'h10 ;
			data[38126] <= 8'h10 ;
			data[38127] <= 8'h10 ;
			data[38128] <= 8'h10 ;
			data[38129] <= 8'h10 ;
			data[38130] <= 8'h10 ;
			data[38131] <= 8'h10 ;
			data[38132] <= 8'h10 ;
			data[38133] <= 8'h10 ;
			data[38134] <= 8'h10 ;
			data[38135] <= 8'h10 ;
			data[38136] <= 8'h10 ;
			data[38137] <= 8'h10 ;
			data[38138] <= 8'h10 ;
			data[38139] <= 8'h10 ;
			data[38140] <= 8'h10 ;
			data[38141] <= 8'h10 ;
			data[38142] <= 8'h10 ;
			data[38143] <= 8'h10 ;
			data[38144] <= 8'h10 ;
			data[38145] <= 8'h10 ;
			data[38146] <= 8'h10 ;
			data[38147] <= 8'h10 ;
			data[38148] <= 8'h10 ;
			data[38149] <= 8'h10 ;
			data[38150] <= 8'h10 ;
			data[38151] <= 8'h10 ;
			data[38152] <= 8'h10 ;
			data[38153] <= 8'h10 ;
			data[38154] <= 8'h10 ;
			data[38155] <= 8'h10 ;
			data[38156] <= 8'h10 ;
			data[38157] <= 8'h10 ;
			data[38158] <= 8'h10 ;
			data[38159] <= 8'h10 ;
			data[38160] <= 8'h10 ;
			data[38161] <= 8'h10 ;
			data[38162] <= 8'h10 ;
			data[38163] <= 8'h10 ;
			data[38164] <= 8'h10 ;
			data[38165] <= 8'h10 ;
			data[38166] <= 8'h10 ;
			data[38167] <= 8'h10 ;
			data[38168] <= 8'h10 ;
			data[38169] <= 8'h10 ;
			data[38170] <= 8'h10 ;
			data[38171] <= 8'h10 ;
			data[38172] <= 8'h10 ;
			data[38173] <= 8'h10 ;
			data[38174] <= 8'h10 ;
			data[38175] <= 8'h10 ;
			data[38176] <= 8'h10 ;
			data[38177] <= 8'h10 ;
			data[38178] <= 8'h10 ;
			data[38179] <= 8'h10 ;
			data[38180] <= 8'h10 ;
			data[38181] <= 8'h10 ;
			data[38182] <= 8'h10 ;
			data[38183] <= 8'h10 ;
			data[38184] <= 8'h10 ;
			data[38185] <= 8'h10 ;
			data[38186] <= 8'h10 ;
			data[38187] <= 8'h10 ;
			data[38188] <= 8'h10 ;
			data[38189] <= 8'h10 ;
			data[38190] <= 8'h10 ;
			data[38191] <= 8'h10 ;
			data[38192] <= 8'h10 ;
			data[38193] <= 8'h10 ;
			data[38194] <= 8'h10 ;
			data[38195] <= 8'h10 ;
			data[38196] <= 8'h10 ;
			data[38197] <= 8'h10 ;
			data[38198] <= 8'h10 ;
			data[38199] <= 8'h10 ;
			data[38200] <= 8'h10 ;
			data[38201] <= 8'h10 ;
			data[38202] <= 8'h10 ;
			data[38203] <= 8'h10 ;
			data[38204] <= 8'h10 ;
			data[38205] <= 8'h10 ;
			data[38206] <= 8'h10 ;
			data[38207] <= 8'h10 ;
			data[38208] <= 8'h10 ;
			data[38209] <= 8'h10 ;
			data[38210] <= 8'h10 ;
			data[38211] <= 8'h10 ;
			data[38212] <= 8'h10 ;
			data[38213] <= 8'h10 ;
			data[38214] <= 8'h10 ;
			data[38215] <= 8'h10 ;
			data[38216] <= 8'h10 ;
			data[38217] <= 8'h10 ;
			data[38218] <= 8'h10 ;
			data[38219] <= 8'h10 ;
			data[38220] <= 8'h10 ;
			data[38221] <= 8'h10 ;
			data[38222] <= 8'h10 ;
			data[38223] <= 8'h10 ;
			data[38224] <= 8'h10 ;
			data[38225] <= 8'h10 ;
			data[38226] <= 8'h10 ;
			data[38227] <= 8'h10 ;
			data[38228] <= 8'h10 ;
			data[38229] <= 8'h10 ;
			data[38230] <= 8'h10 ;
			data[38231] <= 8'h10 ;
			data[38232] <= 8'h10 ;
			data[38233] <= 8'h10 ;
			data[38234] <= 8'h10 ;
			data[38235] <= 8'h10 ;
			data[38236] <= 8'h10 ;
			data[38237] <= 8'h10 ;
			data[38238] <= 8'h10 ;
			data[38239] <= 8'h10 ;
			data[38240] <= 8'h10 ;
			data[38241] <= 8'h10 ;
			data[38242] <= 8'h10 ;
			data[38243] <= 8'h10 ;
			data[38244] <= 8'h10 ;
			data[38245] <= 8'h10 ;
			data[38246] <= 8'h10 ;
			data[38247] <= 8'h10 ;
			data[38248] <= 8'h10 ;
			data[38249] <= 8'h10 ;
			data[38250] <= 8'h10 ;
			data[38251] <= 8'h10 ;
			data[38252] <= 8'h10 ;
			data[38253] <= 8'h10 ;
			data[38254] <= 8'h10 ;
			data[38255] <= 8'h10 ;
			data[38256] <= 8'h10 ;
			data[38257] <= 8'h10 ;
			data[38258] <= 8'h10 ;
			data[38259] <= 8'h10 ;
			data[38260] <= 8'h10 ;
			data[38261] <= 8'h10 ;
			data[38262] <= 8'h10 ;
			data[38263] <= 8'h10 ;
			data[38264] <= 8'h10 ;
			data[38265] <= 8'h10 ;
			data[38266] <= 8'h10 ;
			data[38267] <= 8'h10 ;
			data[38268] <= 8'h10 ;
			data[38269] <= 8'h10 ;
			data[38270] <= 8'h10 ;
			data[38271] <= 8'h10 ;
			data[38272] <= 8'h10 ;
			data[38273] <= 8'h10 ;
			data[38274] <= 8'h10 ;
			data[38275] <= 8'h10 ;
			data[38276] <= 8'h10 ;
			data[38277] <= 8'h10 ;
			data[38278] <= 8'h10 ;
			data[38279] <= 8'h10 ;
			data[38280] <= 8'h10 ;
			data[38281] <= 8'h10 ;
			data[38282] <= 8'h10 ;
			data[38283] <= 8'h10 ;
			data[38284] <= 8'h10 ;
			data[38285] <= 8'h10 ;
			data[38286] <= 8'h10 ;
			data[38287] <= 8'h10 ;
			data[38288] <= 8'h10 ;
			data[38289] <= 8'h10 ;
			data[38290] <= 8'h10 ;
			data[38291] <= 8'h10 ;
			data[38292] <= 8'h10 ;
			data[38293] <= 8'h10 ;
			data[38294] <= 8'h10 ;
			data[38295] <= 8'h10 ;
			data[38296] <= 8'h10 ;
			data[38297] <= 8'h10 ;
			data[38298] <= 8'h10 ;
			data[38299] <= 8'h10 ;
			data[38300] <= 8'h10 ;
			data[38301] <= 8'h10 ;
			data[38302] <= 8'h10 ;
			data[38303] <= 8'h10 ;
			data[38304] <= 8'h10 ;
			data[38305] <= 8'h10 ;
			data[38306] <= 8'h10 ;
			data[38307] <= 8'h10 ;
			data[38308] <= 8'h10 ;
			data[38309] <= 8'h10 ;
			data[38310] <= 8'h10 ;
			data[38311] <= 8'h10 ;
			data[38312] <= 8'h10 ;
			data[38313] <= 8'h10 ;
			data[38314] <= 8'h10 ;
			data[38315] <= 8'h10 ;
			data[38316] <= 8'h10 ;
			data[38317] <= 8'h10 ;
			data[38318] <= 8'h10 ;
			data[38319] <= 8'h10 ;
			data[38320] <= 8'h10 ;
			data[38321] <= 8'h10 ;
			data[38322] <= 8'h10 ;
			data[38323] <= 8'h10 ;
			data[38324] <= 8'h10 ;
			data[38325] <= 8'h10 ;
			data[38326] <= 8'h10 ;
			data[38327] <= 8'h10 ;
			data[38328] <= 8'h10 ;
			data[38329] <= 8'h10 ;
			data[38330] <= 8'h10 ;
			data[38331] <= 8'h10 ;
			data[38332] <= 8'h10 ;
			data[38333] <= 8'h10 ;
			data[38334] <= 8'h10 ;
			data[38335] <= 8'h10 ;
			data[38336] <= 8'h10 ;
			data[38337] <= 8'h10 ;
			data[38338] <= 8'h10 ;
			data[38339] <= 8'h10 ;
			data[38340] <= 8'h10 ;
			data[38341] <= 8'h10 ;
			data[38342] <= 8'h10 ;
			data[38343] <= 8'h10 ;
			data[38344] <= 8'h10 ;
			data[38345] <= 8'h10 ;
			data[38346] <= 8'h10 ;
			data[38347] <= 8'h10 ;
			data[38348] <= 8'h10 ;
			data[38349] <= 8'h10 ;
			data[38350] <= 8'h10 ;
			data[38351] <= 8'h10 ;
			data[38352] <= 8'h10 ;
			data[38353] <= 8'h10 ;
			data[38354] <= 8'h10 ;
			data[38355] <= 8'h10 ;
			data[38356] <= 8'h10 ;
			data[38357] <= 8'h10 ;
			data[38358] <= 8'h10 ;
			data[38359] <= 8'h10 ;
			data[38360] <= 8'h10 ;
			data[38361] <= 8'h10 ;
			data[38362] <= 8'h10 ;
			data[38363] <= 8'h10 ;
			data[38364] <= 8'h10 ;
			data[38365] <= 8'h10 ;
			data[38366] <= 8'h10 ;
			data[38367] <= 8'h10 ;
			data[38368] <= 8'h10 ;
			data[38369] <= 8'h10 ;
			data[38370] <= 8'h10 ;
			data[38371] <= 8'h10 ;
			data[38372] <= 8'h10 ;
			data[38373] <= 8'h10 ;
			data[38374] <= 8'h10 ;
			data[38375] <= 8'h10 ;
			data[38376] <= 8'h10 ;
			data[38377] <= 8'h10 ;
			data[38378] <= 8'h10 ;
			data[38379] <= 8'h10 ;
			data[38380] <= 8'h10 ;
			data[38381] <= 8'h10 ;
			data[38382] <= 8'h10 ;
			data[38383] <= 8'h10 ;
			data[38384] <= 8'h10 ;
			data[38385] <= 8'h10 ;
			data[38386] <= 8'h10 ;
			data[38387] <= 8'h10 ;
			data[38388] <= 8'h10 ;
			data[38389] <= 8'h10 ;
			data[38390] <= 8'h10 ;
			data[38391] <= 8'h10 ;
			data[38392] <= 8'h10 ;
			data[38393] <= 8'h10 ;
			data[38394] <= 8'h10 ;
			data[38395] <= 8'h10 ;
			data[38396] <= 8'h10 ;
			data[38397] <= 8'h10 ;
			data[38398] <= 8'h10 ;
			data[38399] <= 8'h10 ;
			data[38400] <= 8'h10 ;
			data[38401] <= 8'h10 ;
			data[38402] <= 8'h10 ;
			data[38403] <= 8'h10 ;
			data[38404] <= 8'h10 ;
			data[38405] <= 8'h10 ;
			data[38406] <= 8'h10 ;
			data[38407] <= 8'h10 ;
			data[38408] <= 8'h10 ;
			data[38409] <= 8'h10 ;
			data[38410] <= 8'h10 ;
			data[38411] <= 8'h10 ;
			data[38412] <= 8'h10 ;
			data[38413] <= 8'h10 ;
			data[38414] <= 8'h10 ;
			data[38415] <= 8'h10 ;
			data[38416] <= 8'h10 ;
			data[38417] <= 8'h10 ;
			data[38418] <= 8'h10 ;
			data[38419] <= 8'h10 ;
			data[38420] <= 8'h10 ;
			data[38421] <= 8'h10 ;
			data[38422] <= 8'h10 ;
			data[38423] <= 8'h10 ;
			data[38424] <= 8'h10 ;
			data[38425] <= 8'h10 ;
			data[38426] <= 8'h10 ;
			data[38427] <= 8'h10 ;
			data[38428] <= 8'h10 ;
			data[38429] <= 8'h10 ;
			data[38430] <= 8'h10 ;
			data[38431] <= 8'h10 ;
			data[38432] <= 8'h10 ;
			data[38433] <= 8'h10 ;
			data[38434] <= 8'h10 ;
			data[38435] <= 8'h10 ;
			data[38436] <= 8'h10 ;
			data[38437] <= 8'h10 ;
			data[38438] <= 8'h10 ;
			data[38439] <= 8'h10 ;
			data[38440] <= 8'h10 ;
			data[38441] <= 8'h10 ;
			data[38442] <= 8'h10 ;
			data[38443] <= 8'h10 ;
			data[38444] <= 8'h10 ;
			data[38445] <= 8'h10 ;
			data[38446] <= 8'h10 ;
			data[38447] <= 8'h10 ;
			data[38448] <= 8'h10 ;
			data[38449] <= 8'h10 ;
			data[38450] <= 8'h10 ;
			data[38451] <= 8'h10 ;
			data[38452] <= 8'h10 ;
			data[38453] <= 8'h10 ;
			data[38454] <= 8'h10 ;
			data[38455] <= 8'h10 ;
			data[38456] <= 8'h10 ;
			data[38457] <= 8'h10 ;
			data[38458] <= 8'h10 ;
			data[38459] <= 8'h10 ;
			data[38460] <= 8'h10 ;
			data[38461] <= 8'h10 ;
			data[38462] <= 8'h10 ;
			data[38463] <= 8'h10 ;
			data[38464] <= 8'h10 ;
			data[38465] <= 8'h10 ;
			data[38466] <= 8'h10 ;
			data[38467] <= 8'h10 ;
			data[38468] <= 8'h10 ;
			data[38469] <= 8'h10 ;
			data[38470] <= 8'h10 ;
			data[38471] <= 8'h10 ;
			data[38472] <= 8'h10 ;
			data[38473] <= 8'h10 ;
			data[38474] <= 8'h10 ;
			data[38475] <= 8'h10 ;
			data[38476] <= 8'h10 ;
			data[38477] <= 8'h10 ;
			data[38478] <= 8'h10 ;
			data[38479] <= 8'h10 ;
			data[38480] <= 8'h10 ;
			data[38481] <= 8'h10 ;
			data[38482] <= 8'h10 ;
			data[38483] <= 8'h10 ;
			data[38484] <= 8'h10 ;
			data[38485] <= 8'h10 ;
			data[38486] <= 8'h10 ;
			data[38487] <= 8'h10 ;
			data[38488] <= 8'h10 ;
			data[38489] <= 8'h10 ;
			data[38490] <= 8'h10 ;
			data[38491] <= 8'h10 ;
			data[38492] <= 8'h10 ;
			data[38493] <= 8'h10 ;
			data[38494] <= 8'h10 ;
			data[38495] <= 8'h10 ;
			data[38496] <= 8'h10 ;
			data[38497] <= 8'h10 ;
			data[38498] <= 8'h10 ;
			data[38499] <= 8'h10 ;
			data[38500] <= 8'h10 ;
			data[38501] <= 8'h10 ;
			data[38502] <= 8'h10 ;
			data[38503] <= 8'h10 ;
			data[38504] <= 8'h10 ;
			data[38505] <= 8'h10 ;
			data[38506] <= 8'h10 ;
			data[38507] <= 8'h10 ;
			data[38508] <= 8'h10 ;
			data[38509] <= 8'h10 ;
			data[38510] <= 8'h10 ;
			data[38511] <= 8'h10 ;
			data[38512] <= 8'h10 ;
			data[38513] <= 8'h10 ;
			data[38514] <= 8'h10 ;
			data[38515] <= 8'h10 ;
			data[38516] <= 8'h10 ;
			data[38517] <= 8'h10 ;
			data[38518] <= 8'h10 ;
			data[38519] <= 8'h10 ;
			data[38520] <= 8'h10 ;
			data[38521] <= 8'h10 ;
			data[38522] <= 8'h10 ;
			data[38523] <= 8'h10 ;
			data[38524] <= 8'h10 ;
			data[38525] <= 8'h10 ;
			data[38526] <= 8'h10 ;
			data[38527] <= 8'h10 ;
			data[38528] <= 8'h10 ;
			data[38529] <= 8'h10 ;
			data[38530] <= 8'h10 ;
			data[38531] <= 8'h10 ;
			data[38532] <= 8'h10 ;
			data[38533] <= 8'h10 ;
			data[38534] <= 8'h10 ;
			data[38535] <= 8'h10 ;
			data[38536] <= 8'h10 ;
			data[38537] <= 8'h10 ;
			data[38538] <= 8'h10 ;
			data[38539] <= 8'h10 ;
			data[38540] <= 8'h10 ;
			data[38541] <= 8'h10 ;
			data[38542] <= 8'h10 ;
			data[38543] <= 8'h10 ;
			data[38544] <= 8'h10 ;
			data[38545] <= 8'h10 ;
			data[38546] <= 8'h10 ;
			data[38547] <= 8'h10 ;
			data[38548] <= 8'h10 ;
			data[38549] <= 8'h10 ;
			data[38550] <= 8'h10 ;
			data[38551] <= 8'h10 ;
			data[38552] <= 8'h10 ;
			data[38553] <= 8'h10 ;
			data[38554] <= 8'h10 ;
			data[38555] <= 8'h10 ;
			data[38556] <= 8'h10 ;
			data[38557] <= 8'h10 ;
			data[38558] <= 8'h10 ;
			data[38559] <= 8'h10 ;
			data[38560] <= 8'h10 ;
			data[38561] <= 8'h10 ;
			data[38562] <= 8'h10 ;
			data[38563] <= 8'h10 ;
			data[38564] <= 8'h10 ;
			data[38565] <= 8'h10 ;
			data[38566] <= 8'h10 ;
			data[38567] <= 8'h10 ;
			data[38568] <= 8'h10 ;
			data[38569] <= 8'h10 ;
			data[38570] <= 8'h10 ;
			data[38571] <= 8'h10 ;
			data[38572] <= 8'h10 ;
			data[38573] <= 8'h10 ;
			data[38574] <= 8'h10 ;
			data[38575] <= 8'h10 ;
			data[38576] <= 8'h10 ;
			data[38577] <= 8'h10 ;
			data[38578] <= 8'h10 ;
			data[38579] <= 8'h10 ;
			data[38580] <= 8'h10 ;
			data[38581] <= 8'h10 ;
			data[38582] <= 8'h10 ;
			data[38583] <= 8'h10 ;
			data[38584] <= 8'h10 ;
			data[38585] <= 8'h10 ;
			data[38586] <= 8'h10 ;
			data[38587] <= 8'h10 ;
			data[38588] <= 8'h10 ;
			data[38589] <= 8'h10 ;
			data[38590] <= 8'h10 ;
			data[38591] <= 8'h10 ;
			data[38592] <= 8'h10 ;
			data[38593] <= 8'h10 ;
			data[38594] <= 8'h10 ;
			data[38595] <= 8'h10 ;
			data[38596] <= 8'h10 ;
			data[38597] <= 8'h10 ;
			data[38598] <= 8'h10 ;
			data[38599] <= 8'h10 ;
			data[38600] <= 8'h10 ;
			data[38601] <= 8'h10 ;
			data[38602] <= 8'h10 ;
			data[38603] <= 8'h10 ;
			data[38604] <= 8'h10 ;
			data[38605] <= 8'h10 ;
			data[38606] <= 8'h10 ;
			data[38607] <= 8'h10 ;
			data[38608] <= 8'h10 ;
			data[38609] <= 8'h10 ;
			data[38610] <= 8'h10 ;
			data[38611] <= 8'h10 ;
			data[38612] <= 8'h10 ;
			data[38613] <= 8'h10 ;
			data[38614] <= 8'h10 ;
			data[38615] <= 8'h10 ;
			data[38616] <= 8'h10 ;
			data[38617] <= 8'h10 ;
			data[38618] <= 8'h10 ;
			data[38619] <= 8'h10 ;
			data[38620] <= 8'h10 ;
			data[38621] <= 8'h10 ;
			data[38622] <= 8'h10 ;
			data[38623] <= 8'h10 ;
			data[38624] <= 8'h10 ;
			data[38625] <= 8'h10 ;
			data[38626] <= 8'h10 ;
			data[38627] <= 8'h10 ;
			data[38628] <= 8'h10 ;
			data[38629] <= 8'h10 ;
			data[38630] <= 8'h10 ;
			data[38631] <= 8'h10 ;
			data[38632] <= 8'h10 ;
			data[38633] <= 8'h10 ;
			data[38634] <= 8'h10 ;
			data[38635] <= 8'h10 ;
			data[38636] <= 8'h10 ;
			data[38637] <= 8'h10 ;
			data[38638] <= 8'h10 ;
			data[38639] <= 8'h10 ;
			data[38640] <= 8'h10 ;
			data[38641] <= 8'h10 ;
			data[38642] <= 8'h10 ;
			data[38643] <= 8'h10 ;
			data[38644] <= 8'h10 ;
			data[38645] <= 8'h10 ;
			data[38646] <= 8'h10 ;
			data[38647] <= 8'h10 ;
			data[38648] <= 8'h10 ;
			data[38649] <= 8'h10 ;
			data[38650] <= 8'h10 ;
			data[38651] <= 8'h10 ;
			data[38652] <= 8'h10 ;
			data[38653] <= 8'h10 ;
			data[38654] <= 8'h10 ;
			data[38655] <= 8'h10 ;
			data[38656] <= 8'h10 ;
			data[38657] <= 8'h10 ;
			data[38658] <= 8'h10 ;
			data[38659] <= 8'h10 ;
			data[38660] <= 8'h10 ;
			data[38661] <= 8'h10 ;
			data[38662] <= 8'h10 ;
			data[38663] <= 8'h10 ;
			data[38664] <= 8'h10 ;
			data[38665] <= 8'h10 ;
			data[38666] <= 8'h10 ;
			data[38667] <= 8'h10 ;
			data[38668] <= 8'h10 ;
			data[38669] <= 8'h10 ;
			data[38670] <= 8'h10 ;
			data[38671] <= 8'h10 ;
			data[38672] <= 8'h10 ;
			data[38673] <= 8'h10 ;
			data[38674] <= 8'h10 ;
			data[38675] <= 8'h10 ;
			data[38676] <= 8'h10 ;
			data[38677] <= 8'h10 ;
			data[38678] <= 8'h10 ;
			data[38679] <= 8'h10 ;
			data[38680] <= 8'h10 ;
			data[38681] <= 8'h10 ;
			data[38682] <= 8'h10 ;
			data[38683] <= 8'h10 ;
			data[38684] <= 8'h10 ;
			data[38685] <= 8'h10 ;
			data[38686] <= 8'h10 ;
			data[38687] <= 8'h10 ;
			data[38688] <= 8'h10 ;
			data[38689] <= 8'h10 ;
			data[38690] <= 8'h10 ;
			data[38691] <= 8'h10 ;
			data[38692] <= 8'h10 ;
			data[38693] <= 8'h10 ;
			data[38694] <= 8'h10 ;
			data[38695] <= 8'h10 ;
			data[38696] <= 8'h10 ;
			data[38697] <= 8'h10 ;
			data[38698] <= 8'h10 ;
			data[38699] <= 8'h10 ;
			data[38700] <= 8'h10 ;
			data[38701] <= 8'h10 ;
			data[38702] <= 8'h10 ;
			data[38703] <= 8'h10 ;
			data[38704] <= 8'h10 ;
			data[38705] <= 8'h10 ;
			data[38706] <= 8'h10 ;
			data[38707] <= 8'h10 ;
			data[38708] <= 8'h10 ;
			data[38709] <= 8'h10 ;
			data[38710] <= 8'h10 ;
			data[38711] <= 8'h10 ;
			data[38712] <= 8'h10 ;
			data[38713] <= 8'h10 ;
			data[38714] <= 8'h10 ;
			data[38715] <= 8'h10 ;
			data[38716] <= 8'h10 ;
			data[38717] <= 8'h10 ;
			data[38718] <= 8'h10 ;
			data[38719] <= 8'h10 ;
			data[38720] <= 8'h10 ;
			data[38721] <= 8'h10 ;
			data[38722] <= 8'h10 ;
			data[38723] <= 8'h10 ;
			data[38724] <= 8'h10 ;
			data[38725] <= 8'h10 ;
			data[38726] <= 8'h10 ;
			data[38727] <= 8'h10 ;
			data[38728] <= 8'h10 ;
			data[38729] <= 8'h10 ;
			data[38730] <= 8'h10 ;
			data[38731] <= 8'h10 ;
			data[38732] <= 8'h10 ;
			data[38733] <= 8'h10 ;
			data[38734] <= 8'h10 ;
			data[38735] <= 8'h10 ;
			data[38736] <= 8'h10 ;
			data[38737] <= 8'h10 ;
			data[38738] <= 8'h10 ;
			data[38739] <= 8'h10 ;
			data[38740] <= 8'h10 ;
			data[38741] <= 8'h10 ;
			data[38742] <= 8'h10 ;
			data[38743] <= 8'h10 ;
			data[38744] <= 8'h10 ;
			data[38745] <= 8'h10 ;
			data[38746] <= 8'h10 ;
			data[38747] <= 8'h10 ;
			data[38748] <= 8'h10 ;
			data[38749] <= 8'h10 ;
			data[38750] <= 8'h10 ;
			data[38751] <= 8'h10 ;
			data[38752] <= 8'h10 ;
			data[38753] <= 8'h10 ;
			data[38754] <= 8'h10 ;
			data[38755] <= 8'h10 ;
			data[38756] <= 8'h10 ;
			data[38757] <= 8'h10 ;
			data[38758] <= 8'h10 ;
			data[38759] <= 8'h10 ;
			data[38760] <= 8'h10 ;
			data[38761] <= 8'h10 ;
			data[38762] <= 8'h10 ;
			data[38763] <= 8'h10 ;
			data[38764] <= 8'h10 ;
			data[38765] <= 8'h10 ;
			data[38766] <= 8'h10 ;
			data[38767] <= 8'h10 ;
			data[38768] <= 8'h10 ;
			data[38769] <= 8'h10 ;
			data[38770] <= 8'h10 ;
			data[38771] <= 8'h10 ;
			data[38772] <= 8'h10 ;
			data[38773] <= 8'h10 ;
			data[38774] <= 8'h10 ;
			data[38775] <= 8'h10 ;
			data[38776] <= 8'h10 ;
			data[38777] <= 8'h10 ;
			data[38778] <= 8'h10 ;
			data[38779] <= 8'h10 ;
			data[38780] <= 8'h10 ;
			data[38781] <= 8'h10 ;
			data[38782] <= 8'h10 ;
			data[38783] <= 8'h10 ;
			data[38784] <= 8'h10 ;
			data[38785] <= 8'h10 ;
			data[38786] <= 8'h10 ;
			data[38787] <= 8'h10 ;
			data[38788] <= 8'h10 ;
			data[38789] <= 8'h10 ;
			data[38790] <= 8'h10 ;
			data[38791] <= 8'h10 ;
			data[38792] <= 8'h10 ;
			data[38793] <= 8'h10 ;
			data[38794] <= 8'h10 ;
			data[38795] <= 8'h10 ;
			data[38796] <= 8'h10 ;
			data[38797] <= 8'h10 ;
			data[38798] <= 8'h10 ;
			data[38799] <= 8'h10 ;
			data[38800] <= 8'h10 ;
			data[38801] <= 8'h10 ;
			data[38802] <= 8'h10 ;
			data[38803] <= 8'h10 ;
			data[38804] <= 8'h10 ;
			data[38805] <= 8'h10 ;
			data[38806] <= 8'h10 ;
			data[38807] <= 8'h10 ;
			data[38808] <= 8'h10 ;
			data[38809] <= 8'h10 ;
			data[38810] <= 8'h10 ;
			data[38811] <= 8'h10 ;
			data[38812] <= 8'h10 ;
			data[38813] <= 8'h10 ;
			data[38814] <= 8'h10 ;
			data[38815] <= 8'h10 ;
			data[38816] <= 8'h10 ;
			data[38817] <= 8'h10 ;
			data[38818] <= 8'h10 ;
			data[38819] <= 8'h10 ;
			data[38820] <= 8'h10 ;
			data[38821] <= 8'h10 ;
			data[38822] <= 8'h10 ;
			data[38823] <= 8'h10 ;
			data[38824] <= 8'h10 ;
			data[38825] <= 8'h10 ;
			data[38826] <= 8'h10 ;
			data[38827] <= 8'h10 ;
			data[38828] <= 8'h10 ;
			data[38829] <= 8'h10 ;
			data[38830] <= 8'h10 ;
			data[38831] <= 8'h10 ;
			data[38832] <= 8'h10 ;
			data[38833] <= 8'h10 ;
			data[38834] <= 8'h10 ;
			data[38835] <= 8'h10 ;
			data[38836] <= 8'h10 ;
			data[38837] <= 8'h10 ;
			data[38838] <= 8'h10 ;
			data[38839] <= 8'h10 ;
			data[38840] <= 8'h10 ;
			data[38841] <= 8'h10 ;
			data[38842] <= 8'h10 ;
			data[38843] <= 8'h10 ;
			data[38844] <= 8'h10 ;
			data[38845] <= 8'h10 ;
			data[38846] <= 8'h10 ;
			data[38847] <= 8'h10 ;
			data[38848] <= 8'h10 ;
			data[38849] <= 8'h10 ;
			data[38850] <= 8'h10 ;
			data[38851] <= 8'h10 ;
			data[38852] <= 8'h10 ;
			data[38853] <= 8'h10 ;
			data[38854] <= 8'h10 ;
			data[38855] <= 8'h10 ;
			data[38856] <= 8'h10 ;
			data[38857] <= 8'h10 ;
			data[38858] <= 8'h10 ;
			data[38859] <= 8'h10 ;
			data[38860] <= 8'h10 ;
			data[38861] <= 8'h10 ;
			data[38862] <= 8'h10 ;
			data[38863] <= 8'h10 ;
			data[38864] <= 8'h10 ;
			data[38865] <= 8'h10 ;
			data[38866] <= 8'h10 ;
			data[38867] <= 8'h10 ;
			data[38868] <= 8'h10 ;
			data[38869] <= 8'h10 ;
			data[38870] <= 8'h10 ;
			data[38871] <= 8'h10 ;
			data[38872] <= 8'h10 ;
			data[38873] <= 8'h10 ;
			data[38874] <= 8'h10 ;
			data[38875] <= 8'h10 ;
			data[38876] <= 8'h10 ;
			data[38877] <= 8'h10 ;
			data[38878] <= 8'h10 ;
			data[38879] <= 8'h10 ;
			data[38880] <= 8'h10 ;
			data[38881] <= 8'h10 ;
			data[38882] <= 8'h10 ;
			data[38883] <= 8'h10 ;
			data[38884] <= 8'h10 ;
			data[38885] <= 8'h10 ;
			data[38886] <= 8'h10 ;
			data[38887] <= 8'h10 ;
			data[38888] <= 8'h10 ;
			data[38889] <= 8'h10 ;
			data[38890] <= 8'h10 ;
			data[38891] <= 8'h10 ;
			data[38892] <= 8'h10 ;
			data[38893] <= 8'h10 ;
			data[38894] <= 8'h10 ;
			data[38895] <= 8'h10 ;
			data[38896] <= 8'h10 ;
			data[38897] <= 8'h10 ;
			data[38898] <= 8'h10 ;
			data[38899] <= 8'h10 ;
			data[38900] <= 8'h10 ;
			data[38901] <= 8'h10 ;
			data[38902] <= 8'h10 ;
			data[38903] <= 8'h10 ;
			data[38904] <= 8'h10 ;
			data[38905] <= 8'h10 ;
			data[38906] <= 8'h10 ;
			data[38907] <= 8'h10 ;
			data[38908] <= 8'h10 ;
			data[38909] <= 8'h10 ;
			data[38910] <= 8'h10 ;
			data[38911] <= 8'h10 ;
			data[38912] <= 8'h10 ;
			data[38913] <= 8'h10 ;
			data[38914] <= 8'h10 ;
			data[38915] <= 8'h10 ;
			data[38916] <= 8'h10 ;
			data[38917] <= 8'h10 ;
			data[38918] <= 8'h10 ;
			data[38919] <= 8'h10 ;
			data[38920] <= 8'h10 ;
			data[38921] <= 8'h10 ;
			data[38922] <= 8'h10 ;
			data[38923] <= 8'h10 ;
			data[38924] <= 8'h10 ;
			data[38925] <= 8'h10 ;
			data[38926] <= 8'h10 ;
			data[38927] <= 8'h10 ;
			data[38928] <= 8'h10 ;
			data[38929] <= 8'h10 ;
			data[38930] <= 8'h10 ;
			data[38931] <= 8'h10 ;
			data[38932] <= 8'h10 ;
			data[38933] <= 8'h10 ;
			data[38934] <= 8'h10 ;
			data[38935] <= 8'h10 ;
			data[38936] <= 8'h10 ;
			data[38937] <= 8'h10 ;
			data[38938] <= 8'h10 ;
			data[38939] <= 8'h10 ;
			data[38940] <= 8'h10 ;
			data[38941] <= 8'h10 ;
			data[38942] <= 8'h10 ;
			data[38943] <= 8'h10 ;
			data[38944] <= 8'h10 ;
			data[38945] <= 8'h10 ;
			data[38946] <= 8'h10 ;
			data[38947] <= 8'h10 ;
			data[38948] <= 8'h10 ;
			data[38949] <= 8'h10 ;
			data[38950] <= 8'h10 ;
			data[38951] <= 8'h10 ;
			data[38952] <= 8'h10 ;
			data[38953] <= 8'h10 ;
			data[38954] <= 8'h10 ;
			data[38955] <= 8'h10 ;
			data[38956] <= 8'h10 ;
			data[38957] <= 8'h10 ;
			data[38958] <= 8'h10 ;
			data[38959] <= 8'h10 ;
			data[38960] <= 8'h10 ;
			data[38961] <= 8'h10 ;
			data[38962] <= 8'h10 ;
			data[38963] <= 8'h10 ;
			data[38964] <= 8'h10 ;
			data[38965] <= 8'h10 ;
			data[38966] <= 8'h10 ;
			data[38967] <= 8'h10 ;
			data[38968] <= 8'h10 ;
			data[38969] <= 8'h10 ;
			data[38970] <= 8'h10 ;
			data[38971] <= 8'h10 ;
			data[38972] <= 8'h10 ;
			data[38973] <= 8'h10 ;
			data[38974] <= 8'h10 ;
			data[38975] <= 8'h10 ;
			data[38976] <= 8'h10 ;
			data[38977] <= 8'h10 ;
			data[38978] <= 8'h10 ;
			data[38979] <= 8'h10 ;
			data[38980] <= 8'h10 ;
			data[38981] <= 8'h10 ;
			data[38982] <= 8'h10 ;
			data[38983] <= 8'h10 ;
			data[38984] <= 8'h10 ;
			data[38985] <= 8'h10 ;
			data[38986] <= 8'h10 ;
			data[38987] <= 8'h10 ;
			data[38988] <= 8'h10 ;
			data[38989] <= 8'h10 ;
			data[38990] <= 8'h10 ;
			data[38991] <= 8'h10 ;
			data[38992] <= 8'h10 ;
			data[38993] <= 8'h10 ;
			data[38994] <= 8'h10 ;
			data[38995] <= 8'h10 ;
			data[38996] <= 8'h10 ;
			data[38997] <= 8'h10 ;
			data[38998] <= 8'h10 ;
			data[38999] <= 8'h10 ;
			data[39000] <= 8'h10 ;
			data[39001] <= 8'h10 ;
			data[39002] <= 8'h10 ;
			data[39003] <= 8'h10 ;
			data[39004] <= 8'h10 ;
			data[39005] <= 8'h10 ;
			data[39006] <= 8'h10 ;
			data[39007] <= 8'h10 ;
			data[39008] <= 8'h10 ;
			data[39009] <= 8'h10 ;
			data[39010] <= 8'h10 ;
			data[39011] <= 8'h10 ;
			data[39012] <= 8'h10 ;
			data[39013] <= 8'h10 ;
			data[39014] <= 8'h10 ;
			data[39015] <= 8'h10 ;
			data[39016] <= 8'h10 ;
			data[39017] <= 8'h10 ;
			data[39018] <= 8'h10 ;
			data[39019] <= 8'h10 ;
			data[39020] <= 8'h10 ;
			data[39021] <= 8'h10 ;
			data[39022] <= 8'h10 ;
			data[39023] <= 8'h10 ;
			data[39024] <= 8'h10 ;
			data[39025] <= 8'h10 ;
			data[39026] <= 8'h10 ;
			data[39027] <= 8'h10 ;
			data[39028] <= 8'h10 ;
			data[39029] <= 8'h10 ;
			data[39030] <= 8'h10 ;
			data[39031] <= 8'h10 ;
			data[39032] <= 8'h10 ;
			data[39033] <= 8'h10 ;
			data[39034] <= 8'h10 ;
			data[39035] <= 8'h10 ;
			data[39036] <= 8'h10 ;
			data[39037] <= 8'h10 ;
			data[39038] <= 8'h10 ;
			data[39039] <= 8'h10 ;
			data[39040] <= 8'h10 ;
			data[39041] <= 8'h10 ;
			data[39042] <= 8'h10 ;
			data[39043] <= 8'h10 ;
			data[39044] <= 8'h10 ;
			data[39045] <= 8'h10 ;
			data[39046] <= 8'h10 ;
			data[39047] <= 8'h10 ;
			data[39048] <= 8'h10 ;
			data[39049] <= 8'h10 ;
			data[39050] <= 8'h10 ;
			data[39051] <= 8'h10 ;
			data[39052] <= 8'h10 ;
			data[39053] <= 8'h10 ;
			data[39054] <= 8'h10 ;
			data[39055] <= 8'h10 ;
			data[39056] <= 8'h10 ;
			data[39057] <= 8'h10 ;
			data[39058] <= 8'h10 ;
			data[39059] <= 8'h10 ;
			data[39060] <= 8'h10 ;
			data[39061] <= 8'h10 ;
			data[39062] <= 8'h10 ;
			data[39063] <= 8'h10 ;
			data[39064] <= 8'h10 ;
			data[39065] <= 8'h10 ;
			data[39066] <= 8'h10 ;
			data[39067] <= 8'h10 ;
			data[39068] <= 8'h10 ;
			data[39069] <= 8'h10 ;
			data[39070] <= 8'h10 ;
			data[39071] <= 8'h10 ;
			data[39072] <= 8'h10 ;
			data[39073] <= 8'h10 ;
			data[39074] <= 8'h10 ;
			data[39075] <= 8'h10 ;
			data[39076] <= 8'h10 ;
			data[39077] <= 8'h10 ;
			data[39078] <= 8'h10 ;
			data[39079] <= 8'h10 ;
			data[39080] <= 8'h10 ;
			data[39081] <= 8'h10 ;
			data[39082] <= 8'h10 ;
			data[39083] <= 8'h10 ;
			data[39084] <= 8'h10 ;
			data[39085] <= 8'h10 ;
			data[39086] <= 8'h10 ;
			data[39087] <= 8'h10 ;
			data[39088] <= 8'h10 ;
			data[39089] <= 8'h10 ;
			data[39090] <= 8'h10 ;
			data[39091] <= 8'h10 ;
			data[39092] <= 8'h10 ;
			data[39093] <= 8'h10 ;
			data[39094] <= 8'h10 ;
			data[39095] <= 8'h10 ;
			data[39096] <= 8'h10 ;
			data[39097] <= 8'h10 ;
			data[39098] <= 8'h10 ;
			data[39099] <= 8'h10 ;
			data[39100] <= 8'h10 ;
			data[39101] <= 8'h10 ;
			data[39102] <= 8'h10 ;
			data[39103] <= 8'h10 ;
			data[39104] <= 8'h10 ;
			data[39105] <= 8'h10 ;
			data[39106] <= 8'h10 ;
			data[39107] <= 8'h10 ;
			data[39108] <= 8'h10 ;
			data[39109] <= 8'h10 ;
			data[39110] <= 8'h10 ;
			data[39111] <= 8'h10 ;
			data[39112] <= 8'h10 ;
			data[39113] <= 8'h10 ;
			data[39114] <= 8'h10 ;
			data[39115] <= 8'h10 ;
			data[39116] <= 8'h10 ;
			data[39117] <= 8'h10 ;
			data[39118] <= 8'h10 ;
			data[39119] <= 8'h10 ;
			data[39120] <= 8'h10 ;
			data[39121] <= 8'h10 ;
			data[39122] <= 8'h10 ;
			data[39123] <= 8'h10 ;
			data[39124] <= 8'h10 ;
			data[39125] <= 8'h10 ;
			data[39126] <= 8'h10 ;
			data[39127] <= 8'h10 ;
			data[39128] <= 8'h10 ;
			data[39129] <= 8'h10 ;
			data[39130] <= 8'h10 ;
			data[39131] <= 8'h10 ;
			data[39132] <= 8'h10 ;
			data[39133] <= 8'h10 ;
			data[39134] <= 8'h10 ;
			data[39135] <= 8'h10 ;
			data[39136] <= 8'h10 ;
			data[39137] <= 8'h10 ;
			data[39138] <= 8'h10 ;
			data[39139] <= 8'h10 ;
			data[39140] <= 8'h10 ;
			data[39141] <= 8'h10 ;
			data[39142] <= 8'h10 ;
			data[39143] <= 8'h10 ;
			data[39144] <= 8'h10 ;
			data[39145] <= 8'h10 ;
			data[39146] <= 8'h10 ;
			data[39147] <= 8'h10 ;
			data[39148] <= 8'h10 ;
			data[39149] <= 8'h10 ;
			data[39150] <= 8'h10 ;
			data[39151] <= 8'h10 ;
			data[39152] <= 8'h10 ;
			data[39153] <= 8'h10 ;
			data[39154] <= 8'h10 ;
			data[39155] <= 8'h10 ;
			data[39156] <= 8'h10 ;
			data[39157] <= 8'h10 ;
			data[39158] <= 8'h10 ;
			data[39159] <= 8'h10 ;
			data[39160] <= 8'h10 ;
			data[39161] <= 8'h10 ;
			data[39162] <= 8'h10 ;
			data[39163] <= 8'h10 ;
			data[39164] <= 8'h10 ;
			data[39165] <= 8'h10 ;
			data[39166] <= 8'h10 ;
			data[39167] <= 8'h10 ;
			data[39168] <= 8'h10 ;
			data[39169] <= 8'h10 ;
			data[39170] <= 8'h10 ;
			data[39171] <= 8'h10 ;
			data[39172] <= 8'h10 ;
			data[39173] <= 8'h10 ;
			data[39174] <= 8'h10 ;
			data[39175] <= 8'h10 ;
			data[39176] <= 8'h10 ;
			data[39177] <= 8'h10 ;
			data[39178] <= 8'h10 ;
			data[39179] <= 8'h10 ;
			data[39180] <= 8'h10 ;
			data[39181] <= 8'h10 ;
			data[39182] <= 8'h10 ;
			data[39183] <= 8'h10 ;
			data[39184] <= 8'h10 ;
			data[39185] <= 8'h10 ;
			data[39186] <= 8'h10 ;
			data[39187] <= 8'h10 ;
			data[39188] <= 8'h10 ;
			data[39189] <= 8'h10 ;
			data[39190] <= 8'h10 ;
			data[39191] <= 8'h10 ;
			data[39192] <= 8'h10 ;
			data[39193] <= 8'h10 ;
			data[39194] <= 8'h10 ;
			data[39195] <= 8'h10 ;
			data[39196] <= 8'h10 ;
			data[39197] <= 8'h10 ;
			data[39198] <= 8'h10 ;
			data[39199] <= 8'h10 ;
			data[39200] <= 8'h10 ;
			data[39201] <= 8'h10 ;
			data[39202] <= 8'h10 ;
			data[39203] <= 8'h10 ;
			data[39204] <= 8'h10 ;
			data[39205] <= 8'h10 ;
			data[39206] <= 8'h10 ;
			data[39207] <= 8'h10 ;
			data[39208] <= 8'h10 ;
			data[39209] <= 8'h10 ;
			data[39210] <= 8'h10 ;
			data[39211] <= 8'h10 ;
			data[39212] <= 8'h10 ;
			data[39213] <= 8'h10 ;
			data[39214] <= 8'h10 ;
			data[39215] <= 8'h10 ;
			data[39216] <= 8'h10 ;
			data[39217] <= 8'h10 ;
			data[39218] <= 8'h10 ;
			data[39219] <= 8'h10 ;
			data[39220] <= 8'h10 ;
			data[39221] <= 8'h10 ;
			data[39222] <= 8'h10 ;
			data[39223] <= 8'h10 ;
			data[39224] <= 8'h10 ;
			data[39225] <= 8'h10 ;
			data[39226] <= 8'h10 ;
			data[39227] <= 8'h10 ;
			data[39228] <= 8'h10 ;
			data[39229] <= 8'h10 ;
			data[39230] <= 8'h10 ;
			data[39231] <= 8'h10 ;
			data[39232] <= 8'h10 ;
			data[39233] <= 8'h10 ;
			data[39234] <= 8'h10 ;
			data[39235] <= 8'h10 ;
			data[39236] <= 8'h10 ;
			data[39237] <= 8'h10 ;
			data[39238] <= 8'h10 ;
			data[39239] <= 8'h10 ;
			data[39240] <= 8'h10 ;
			data[39241] <= 8'h10 ;
			data[39242] <= 8'h10 ;
			data[39243] <= 8'h10 ;
			data[39244] <= 8'h10 ;
			data[39245] <= 8'h10 ;
			data[39246] <= 8'h10 ;
			data[39247] <= 8'h10 ;
			data[39248] <= 8'h10 ;
			data[39249] <= 8'h10 ;
			data[39250] <= 8'h10 ;
			data[39251] <= 8'h10 ;
			data[39252] <= 8'h10 ;
			data[39253] <= 8'h10 ;
			data[39254] <= 8'h10 ;
			data[39255] <= 8'h10 ;
			data[39256] <= 8'h10 ;
			data[39257] <= 8'h10 ;
			data[39258] <= 8'h10 ;
			data[39259] <= 8'h10 ;
			data[39260] <= 8'h10 ;
			data[39261] <= 8'h10 ;
			data[39262] <= 8'h10 ;
			data[39263] <= 8'h10 ;
			data[39264] <= 8'h10 ;
			data[39265] <= 8'h10 ;
			data[39266] <= 8'h10 ;
			data[39267] <= 8'h10 ;
			data[39268] <= 8'h10 ;
			data[39269] <= 8'h10 ;
			data[39270] <= 8'h10 ;
			data[39271] <= 8'h10 ;
			data[39272] <= 8'h10 ;
			data[39273] <= 8'h10 ;
			data[39274] <= 8'h10 ;
			data[39275] <= 8'h10 ;
			data[39276] <= 8'h10 ;
			data[39277] <= 8'h10 ;
			data[39278] <= 8'h10 ;
			data[39279] <= 8'h10 ;
			data[39280] <= 8'h10 ;
			data[39281] <= 8'h10 ;
			data[39282] <= 8'h10 ;
			data[39283] <= 8'h10 ;
			data[39284] <= 8'h10 ;
			data[39285] <= 8'h10 ;
			data[39286] <= 8'h10 ;
			data[39287] <= 8'h10 ;
			data[39288] <= 8'h10 ;
			data[39289] <= 8'h10 ;
			data[39290] <= 8'h10 ;
			data[39291] <= 8'h10 ;
			data[39292] <= 8'h10 ;
			data[39293] <= 8'h10 ;
			data[39294] <= 8'h10 ;
			data[39295] <= 8'h10 ;
			data[39296] <= 8'h10 ;
			data[39297] <= 8'h10 ;
			data[39298] <= 8'h10 ;
			data[39299] <= 8'h10 ;
			data[39300] <= 8'h10 ;
			data[39301] <= 8'h10 ;
			data[39302] <= 8'h10 ;
			data[39303] <= 8'h10 ;
			data[39304] <= 8'h10 ;
			data[39305] <= 8'h10 ;
			data[39306] <= 8'h10 ;
			data[39307] <= 8'h10 ;
			data[39308] <= 8'h10 ;
			data[39309] <= 8'h10 ;
			data[39310] <= 8'h10 ;
			data[39311] <= 8'h10 ;
			data[39312] <= 8'h10 ;
			data[39313] <= 8'h10 ;
			data[39314] <= 8'h10 ;
			data[39315] <= 8'h10 ;
			data[39316] <= 8'h10 ;
			data[39317] <= 8'h10 ;
			data[39318] <= 8'h10 ;
			data[39319] <= 8'h10 ;
			data[39320] <= 8'h10 ;
			data[39321] <= 8'h10 ;
			data[39322] <= 8'h10 ;
			data[39323] <= 8'h10 ;
			data[39324] <= 8'h10 ;
			data[39325] <= 8'h10 ;
			data[39326] <= 8'h10 ;
			data[39327] <= 8'h10 ;
			data[39328] <= 8'h10 ;
			data[39329] <= 8'h10 ;
			data[39330] <= 8'h10 ;
			data[39331] <= 8'h10 ;
			data[39332] <= 8'h10 ;
			data[39333] <= 8'h10 ;
			data[39334] <= 8'h10 ;
			data[39335] <= 8'h10 ;
			data[39336] <= 8'h10 ;
			data[39337] <= 8'h10 ;
			data[39338] <= 8'h10 ;
			data[39339] <= 8'h10 ;
			data[39340] <= 8'h10 ;
			data[39341] <= 8'h10 ;
			data[39342] <= 8'h10 ;
			data[39343] <= 8'h10 ;
			data[39344] <= 8'h10 ;
			data[39345] <= 8'h10 ;
			data[39346] <= 8'h10 ;
			data[39347] <= 8'h10 ;
			data[39348] <= 8'h10 ;
			data[39349] <= 8'h10 ;
			data[39350] <= 8'h10 ;
			data[39351] <= 8'h10 ;
			data[39352] <= 8'h10 ;
			data[39353] <= 8'h10 ;
			data[39354] <= 8'h10 ;
			data[39355] <= 8'h10 ;
			data[39356] <= 8'h10 ;
			data[39357] <= 8'h10 ;
			data[39358] <= 8'h10 ;
			data[39359] <= 8'h10 ;
			data[39360] <= 8'h10 ;
			data[39361] <= 8'h10 ;
			data[39362] <= 8'h10 ;
			data[39363] <= 8'h10 ;
			data[39364] <= 8'h10 ;
			data[39365] <= 8'h10 ;
			data[39366] <= 8'h10 ;
			data[39367] <= 8'h10 ;
			data[39368] <= 8'h10 ;
			data[39369] <= 8'h10 ;
			data[39370] <= 8'h10 ;
			data[39371] <= 8'h10 ;
			data[39372] <= 8'h10 ;
			data[39373] <= 8'h10 ;
			data[39374] <= 8'h10 ;
			data[39375] <= 8'h10 ;
			data[39376] <= 8'h10 ;
			data[39377] <= 8'h10 ;
			data[39378] <= 8'h10 ;
			data[39379] <= 8'h10 ;
			data[39380] <= 8'h10 ;
			data[39381] <= 8'h10 ;
			data[39382] <= 8'h10 ;
			data[39383] <= 8'h10 ;
			data[39384] <= 8'h10 ;
			data[39385] <= 8'h10 ;
			data[39386] <= 8'h10 ;
			data[39387] <= 8'h10 ;
			data[39388] <= 8'h10 ;
			data[39389] <= 8'h10 ;
			data[39390] <= 8'h10 ;
			data[39391] <= 8'h10 ;
			data[39392] <= 8'h10 ;
			data[39393] <= 8'h10 ;
			data[39394] <= 8'h10 ;
			data[39395] <= 8'h10 ;
			data[39396] <= 8'h10 ;
			data[39397] <= 8'h10 ;
			data[39398] <= 8'h10 ;
			data[39399] <= 8'h10 ;
			data[39400] <= 8'h10 ;
			data[39401] <= 8'h10 ;
			data[39402] <= 8'h10 ;
			data[39403] <= 8'h10 ;
			data[39404] <= 8'h10 ;
			data[39405] <= 8'h10 ;
			data[39406] <= 8'h10 ;
			data[39407] <= 8'h10 ;
			data[39408] <= 8'h10 ;
			data[39409] <= 8'h10 ;
			data[39410] <= 8'h10 ;
			data[39411] <= 8'h10 ;
			data[39412] <= 8'h10 ;
			data[39413] <= 8'h10 ;
			data[39414] <= 8'h10 ;
			data[39415] <= 8'h10 ;
			data[39416] <= 8'h10 ;
			data[39417] <= 8'h10 ;
			data[39418] <= 8'h10 ;
			data[39419] <= 8'h10 ;
			data[39420] <= 8'h10 ;
			data[39421] <= 8'h10 ;
			data[39422] <= 8'h10 ;
			data[39423] <= 8'h10 ;
			data[39424] <= 8'h10 ;
			data[39425] <= 8'h10 ;
			data[39426] <= 8'h10 ;
			data[39427] <= 8'h10 ;
			data[39428] <= 8'h10 ;
			data[39429] <= 8'h10 ;
			data[39430] <= 8'h10 ;
			data[39431] <= 8'h10 ;
			data[39432] <= 8'h10 ;
			data[39433] <= 8'h10 ;
			data[39434] <= 8'h10 ;
			data[39435] <= 8'h10 ;
			data[39436] <= 8'h10 ;
			data[39437] <= 8'h10 ;
			data[39438] <= 8'h10 ;
			data[39439] <= 8'h10 ;
			data[39440] <= 8'h10 ;
			data[39441] <= 8'h10 ;
			data[39442] <= 8'h10 ;
			data[39443] <= 8'h10 ;
			data[39444] <= 8'h10 ;
			data[39445] <= 8'h10 ;
			data[39446] <= 8'h10 ;
			data[39447] <= 8'h10 ;
			data[39448] <= 8'h10 ;
			data[39449] <= 8'h10 ;
			data[39450] <= 8'h10 ;
			data[39451] <= 8'h10 ;
			data[39452] <= 8'h10 ;
			data[39453] <= 8'h10 ;
			data[39454] <= 8'h10 ;
			data[39455] <= 8'h10 ;
			data[39456] <= 8'h10 ;
			data[39457] <= 8'h10 ;
			data[39458] <= 8'h10 ;
			data[39459] <= 8'h10 ;
			data[39460] <= 8'h10 ;
			data[39461] <= 8'h10 ;
			data[39462] <= 8'h10 ;
			data[39463] <= 8'h10 ;
			data[39464] <= 8'h10 ;
			data[39465] <= 8'h10 ;
			data[39466] <= 8'h10 ;
			data[39467] <= 8'h10 ;
			data[39468] <= 8'h10 ;
			data[39469] <= 8'h10 ;
			data[39470] <= 8'h10 ;
			data[39471] <= 8'h10 ;
			data[39472] <= 8'h10 ;
			data[39473] <= 8'h10 ;
			data[39474] <= 8'h10 ;
			data[39475] <= 8'h10 ;
			data[39476] <= 8'h10 ;
			data[39477] <= 8'h10 ;
			data[39478] <= 8'h10 ;
			data[39479] <= 8'h10 ;
			data[39480] <= 8'h10 ;
			data[39481] <= 8'h10 ;
			data[39482] <= 8'h10 ;
			data[39483] <= 8'h10 ;
			data[39484] <= 8'h10 ;
			data[39485] <= 8'h10 ;
			data[39486] <= 8'h10 ;
			data[39487] <= 8'h10 ;
			data[39488] <= 8'h10 ;
			data[39489] <= 8'h10 ;
			data[39490] <= 8'h10 ;
			data[39491] <= 8'h10 ;
			data[39492] <= 8'h10 ;
			data[39493] <= 8'h10 ;
			data[39494] <= 8'h10 ;
			data[39495] <= 8'h10 ;
			data[39496] <= 8'h10 ;
			data[39497] <= 8'h10 ;
			data[39498] <= 8'h10 ;
			data[39499] <= 8'h10 ;
			data[39500] <= 8'h10 ;
			data[39501] <= 8'h10 ;
			data[39502] <= 8'h10 ;
			data[39503] <= 8'h10 ;
			data[39504] <= 8'h10 ;
			data[39505] <= 8'h10 ;
			data[39506] <= 8'h10 ;
			data[39507] <= 8'h10 ;
			data[39508] <= 8'h10 ;
			data[39509] <= 8'h10 ;
			data[39510] <= 8'h10 ;
			data[39511] <= 8'h10 ;
			data[39512] <= 8'h10 ;
			data[39513] <= 8'h10 ;
			data[39514] <= 8'h10 ;
			data[39515] <= 8'h10 ;
			data[39516] <= 8'h10 ;
			data[39517] <= 8'h10 ;
			data[39518] <= 8'h10 ;
			data[39519] <= 8'h10 ;
			data[39520] <= 8'h10 ;
			data[39521] <= 8'h10 ;
			data[39522] <= 8'h10 ;
			data[39523] <= 8'h10 ;
			data[39524] <= 8'h10 ;
			data[39525] <= 8'h10 ;
			data[39526] <= 8'h10 ;
			data[39527] <= 8'h10 ;
			data[39528] <= 8'h10 ;
			data[39529] <= 8'h10 ;
			data[39530] <= 8'h10 ;
			data[39531] <= 8'h10 ;
			data[39532] <= 8'h10 ;
			data[39533] <= 8'h10 ;
			data[39534] <= 8'h10 ;
			data[39535] <= 8'h10 ;
			data[39536] <= 8'h10 ;
			data[39537] <= 8'h10 ;
			data[39538] <= 8'h10 ;
			data[39539] <= 8'h10 ;
			data[39540] <= 8'h10 ;
			data[39541] <= 8'h10 ;
			data[39542] <= 8'h10 ;
			data[39543] <= 8'h10 ;
			data[39544] <= 8'h10 ;
			data[39545] <= 8'h10 ;
			data[39546] <= 8'h10 ;
			data[39547] <= 8'h10 ;
			data[39548] <= 8'h10 ;
			data[39549] <= 8'h10 ;
			data[39550] <= 8'h10 ;
			data[39551] <= 8'h10 ;
			data[39552] <= 8'h10 ;
			data[39553] <= 8'h10 ;
			data[39554] <= 8'h10 ;
			data[39555] <= 8'h10 ;
			data[39556] <= 8'h10 ;
			data[39557] <= 8'h10 ;
			data[39558] <= 8'h10 ;
			data[39559] <= 8'h10 ;
			data[39560] <= 8'h10 ;
			data[39561] <= 8'h10 ;
			data[39562] <= 8'h10 ;
			data[39563] <= 8'h10 ;
			data[39564] <= 8'h10 ;
			data[39565] <= 8'h10 ;
			data[39566] <= 8'h10 ;
			data[39567] <= 8'h10 ;
			data[39568] <= 8'h10 ;
			data[39569] <= 8'h10 ;
			data[39570] <= 8'h10 ;
			data[39571] <= 8'h10 ;
			data[39572] <= 8'h10 ;
			data[39573] <= 8'h10 ;
			data[39574] <= 8'h10 ;
			data[39575] <= 8'h10 ;
			data[39576] <= 8'h10 ;
			data[39577] <= 8'h10 ;
			data[39578] <= 8'h10 ;
			data[39579] <= 8'h10 ;
			data[39580] <= 8'h10 ;
			data[39581] <= 8'h10 ;
			data[39582] <= 8'h10 ;
			data[39583] <= 8'h10 ;
			data[39584] <= 8'h10 ;
			data[39585] <= 8'h10 ;
			data[39586] <= 8'h10 ;
			data[39587] <= 8'h10 ;
			data[39588] <= 8'h10 ;
			data[39589] <= 8'h10 ;
			data[39590] <= 8'h10 ;
			data[39591] <= 8'h10 ;
			data[39592] <= 8'h10 ;
			data[39593] <= 8'h10 ;
			data[39594] <= 8'h10 ;
			data[39595] <= 8'h10 ;
			data[39596] <= 8'h10 ;
			data[39597] <= 8'h10 ;
			data[39598] <= 8'h10 ;
			data[39599] <= 8'h10 ;
			data[39600] <= 8'h10 ;
			data[39601] <= 8'h10 ;
			data[39602] <= 8'h10 ;
			data[39603] <= 8'h10 ;
			data[39604] <= 8'h10 ;
			data[39605] <= 8'h10 ;
			data[39606] <= 8'h10 ;
			data[39607] <= 8'h10 ;
			data[39608] <= 8'h10 ;
			data[39609] <= 8'h10 ;
			data[39610] <= 8'h10 ;
			data[39611] <= 8'h10 ;
			data[39612] <= 8'h10 ;
			data[39613] <= 8'h10 ;
			data[39614] <= 8'h10 ;
			data[39615] <= 8'h10 ;
			data[39616] <= 8'h10 ;
			data[39617] <= 8'h10 ;
			data[39618] <= 8'h10 ;
			data[39619] <= 8'h10 ;
			data[39620] <= 8'h10 ;
			data[39621] <= 8'h10 ;
			data[39622] <= 8'h10 ;
			data[39623] <= 8'h10 ;
			data[39624] <= 8'h10 ;
			data[39625] <= 8'h10 ;
			data[39626] <= 8'h10 ;
			data[39627] <= 8'h10 ;
			data[39628] <= 8'h10 ;
			data[39629] <= 8'h10 ;
			data[39630] <= 8'h10 ;
			data[39631] <= 8'h10 ;
			data[39632] <= 8'h10 ;
			data[39633] <= 8'h10 ;
			data[39634] <= 8'h10 ;
			data[39635] <= 8'h10 ;
			data[39636] <= 8'h10 ;
			data[39637] <= 8'h10 ;
			data[39638] <= 8'h10 ;
			data[39639] <= 8'h10 ;
			data[39640] <= 8'h10 ;
			data[39641] <= 8'h10 ;
			data[39642] <= 8'h10 ;
			data[39643] <= 8'h10 ;
			data[39644] <= 8'h10 ;
			data[39645] <= 8'h10 ;
			data[39646] <= 8'h10 ;
			data[39647] <= 8'h10 ;
			data[39648] <= 8'h10 ;
			data[39649] <= 8'h10 ;
			data[39650] <= 8'h10 ;
			data[39651] <= 8'h10 ;
			data[39652] <= 8'h10 ;
			data[39653] <= 8'h10 ;
			data[39654] <= 8'h10 ;
			data[39655] <= 8'h10 ;
			data[39656] <= 8'h10 ;
			data[39657] <= 8'h10 ;
			data[39658] <= 8'h10 ;
			data[39659] <= 8'h10 ;
			data[39660] <= 8'h10 ;
			data[39661] <= 8'h10 ;
			data[39662] <= 8'h10 ;
			data[39663] <= 8'h10 ;
			data[39664] <= 8'h10 ;
			data[39665] <= 8'h10 ;
			data[39666] <= 8'h10 ;
			data[39667] <= 8'h10 ;
			data[39668] <= 8'h10 ;
			data[39669] <= 8'h10 ;
			data[39670] <= 8'h10 ;
			data[39671] <= 8'h10 ;
			data[39672] <= 8'h10 ;
			data[39673] <= 8'h10 ;
			data[39674] <= 8'h10 ;
			data[39675] <= 8'h10 ;
			data[39676] <= 8'h10 ;
			data[39677] <= 8'h10 ;
			data[39678] <= 8'h10 ;
			data[39679] <= 8'h10 ;
			data[39680] <= 8'h10 ;
			data[39681] <= 8'h10 ;
			data[39682] <= 8'h10 ;
			data[39683] <= 8'h10 ;
			data[39684] <= 8'h10 ;
			data[39685] <= 8'h10 ;
			data[39686] <= 8'h10 ;
			data[39687] <= 8'h10 ;
			data[39688] <= 8'h10 ;
			data[39689] <= 8'h10 ;
			data[39690] <= 8'h10 ;
			data[39691] <= 8'h10 ;
			data[39692] <= 8'h10 ;
			data[39693] <= 8'h10 ;
			data[39694] <= 8'h10 ;
			data[39695] <= 8'h10 ;
			data[39696] <= 8'h10 ;
			data[39697] <= 8'h10 ;
			data[39698] <= 8'h10 ;
			data[39699] <= 8'h10 ;
			data[39700] <= 8'h10 ;
			data[39701] <= 8'h10 ;
			data[39702] <= 8'h10 ;
			data[39703] <= 8'h10 ;
			data[39704] <= 8'h10 ;
			data[39705] <= 8'h10 ;
			data[39706] <= 8'h10 ;
			data[39707] <= 8'h10 ;
			data[39708] <= 8'h10 ;
			data[39709] <= 8'h10 ;
			data[39710] <= 8'h10 ;
			data[39711] <= 8'h10 ;
			data[39712] <= 8'h10 ;
			data[39713] <= 8'h10 ;
			data[39714] <= 8'h10 ;
			data[39715] <= 8'h10 ;
			data[39716] <= 8'h10 ;
			data[39717] <= 8'h10 ;
			data[39718] <= 8'h10 ;
			data[39719] <= 8'h10 ;
			data[39720] <= 8'h10 ;
			data[39721] <= 8'h10 ;
			data[39722] <= 8'h10 ;
			data[39723] <= 8'h10 ;
			data[39724] <= 8'h10 ;
			data[39725] <= 8'h10 ;
			data[39726] <= 8'h10 ;
			data[39727] <= 8'h10 ;
			data[39728] <= 8'h10 ;
			data[39729] <= 8'h10 ;
			data[39730] <= 8'h10 ;
			data[39731] <= 8'h10 ;
			data[39732] <= 8'h10 ;
			data[39733] <= 8'h10 ;
			data[39734] <= 8'h10 ;
			data[39735] <= 8'h10 ;
			data[39736] <= 8'h10 ;
			data[39737] <= 8'h10 ;
			data[39738] <= 8'h10 ;
			data[39739] <= 8'h10 ;
			data[39740] <= 8'h10 ;
			data[39741] <= 8'h10 ;
			data[39742] <= 8'h10 ;
			data[39743] <= 8'h10 ;
			data[39744] <= 8'h10 ;
			data[39745] <= 8'h10 ;
			data[39746] <= 8'h10 ;
			data[39747] <= 8'h10 ;
			data[39748] <= 8'h10 ;
			data[39749] <= 8'h10 ;
			data[39750] <= 8'h10 ;
			data[39751] <= 8'h10 ;
			data[39752] <= 8'h10 ;
			data[39753] <= 8'h10 ;
			data[39754] <= 8'h10 ;
			data[39755] <= 8'h10 ;
			data[39756] <= 8'h10 ;
			data[39757] <= 8'h10 ;
			data[39758] <= 8'h10 ;
			data[39759] <= 8'h10 ;
			data[39760] <= 8'h10 ;
			data[39761] <= 8'h10 ;
			data[39762] <= 8'h10 ;
			data[39763] <= 8'h10 ;
			data[39764] <= 8'h10 ;
			data[39765] <= 8'h10 ;
			data[39766] <= 8'h10 ;
			data[39767] <= 8'h10 ;
			data[39768] <= 8'h10 ;
			data[39769] <= 8'h10 ;
			data[39770] <= 8'h10 ;
			data[39771] <= 8'h10 ;
			data[39772] <= 8'h10 ;
			data[39773] <= 8'h10 ;
			data[39774] <= 8'h10 ;
			data[39775] <= 8'h10 ;
			data[39776] <= 8'h10 ;
			data[39777] <= 8'h10 ;
			data[39778] <= 8'h10 ;
			data[39779] <= 8'h10 ;
			data[39780] <= 8'h10 ;
			data[39781] <= 8'h10 ;
			data[39782] <= 8'h10 ;
			data[39783] <= 8'h10 ;
			data[39784] <= 8'h10 ;
			data[39785] <= 8'h10 ;
			data[39786] <= 8'h10 ;
			data[39787] <= 8'h10 ;
			data[39788] <= 8'h10 ;
			data[39789] <= 8'h10 ;
			data[39790] <= 8'h10 ;
			data[39791] <= 8'h10 ;
			data[39792] <= 8'h10 ;
			data[39793] <= 8'h10 ;
			data[39794] <= 8'h10 ;
			data[39795] <= 8'h10 ;
			data[39796] <= 8'h10 ;
			data[39797] <= 8'h10 ;
			data[39798] <= 8'h10 ;
			data[39799] <= 8'h10 ;
			data[39800] <= 8'h10 ;
			data[39801] <= 8'h10 ;
			data[39802] <= 8'h10 ;
			data[39803] <= 8'h10 ;
			data[39804] <= 8'h10 ;
			data[39805] <= 8'h10 ;
			data[39806] <= 8'h10 ;
			data[39807] <= 8'h10 ;
			data[39808] <= 8'h10 ;
			data[39809] <= 8'h10 ;
			data[39810] <= 8'h10 ;
			data[39811] <= 8'h10 ;
			data[39812] <= 8'h10 ;
			data[39813] <= 8'h10 ;
			data[39814] <= 8'h10 ;
			data[39815] <= 8'h10 ;
			data[39816] <= 8'h10 ;
			data[39817] <= 8'h10 ;
			data[39818] <= 8'h10 ;
			data[39819] <= 8'h10 ;
			data[39820] <= 8'h10 ;
			data[39821] <= 8'h10 ;
			data[39822] <= 8'h10 ;
			data[39823] <= 8'h10 ;
			data[39824] <= 8'h10 ;
			data[39825] <= 8'h10 ;
			data[39826] <= 8'h10 ;
			data[39827] <= 8'h10 ;
			data[39828] <= 8'h10 ;
			data[39829] <= 8'h10 ;
			data[39830] <= 8'h10 ;
			data[39831] <= 8'h10 ;
			data[39832] <= 8'h10 ;
			data[39833] <= 8'h10 ;
			data[39834] <= 8'h10 ;
			data[39835] <= 8'h10 ;
			data[39836] <= 8'h10 ;
			data[39837] <= 8'h10 ;
			data[39838] <= 8'h10 ;
			data[39839] <= 8'h10 ;
			data[39840] <= 8'h10 ;
			data[39841] <= 8'h10 ;
			data[39842] <= 8'h10 ;
			data[39843] <= 8'h10 ;
			data[39844] <= 8'h10 ;
			data[39845] <= 8'h10 ;
			data[39846] <= 8'h10 ;
			data[39847] <= 8'h10 ;
			data[39848] <= 8'h10 ;
			data[39849] <= 8'h10 ;
			data[39850] <= 8'h10 ;
			data[39851] <= 8'h10 ;
			data[39852] <= 8'h10 ;
			data[39853] <= 8'h10 ;
			data[39854] <= 8'h10 ;
			data[39855] <= 8'h10 ;
			data[39856] <= 8'h10 ;
			data[39857] <= 8'h10 ;
			data[39858] <= 8'h10 ;
			data[39859] <= 8'h10 ;
			data[39860] <= 8'h10 ;
			data[39861] <= 8'h10 ;
			data[39862] <= 8'h10 ;
			data[39863] <= 8'h10 ;
			data[39864] <= 8'h10 ;
			data[39865] <= 8'h10 ;
			data[39866] <= 8'h10 ;
			data[39867] <= 8'h10 ;
			data[39868] <= 8'h10 ;
			data[39869] <= 8'h10 ;
			data[39870] <= 8'h10 ;
			data[39871] <= 8'h10 ;
			data[39872] <= 8'h10 ;
			data[39873] <= 8'h10 ;
			data[39874] <= 8'h10 ;
			data[39875] <= 8'h10 ;
			data[39876] <= 8'h10 ;
			data[39877] <= 8'h10 ;
			data[39878] <= 8'h10 ;
			data[39879] <= 8'h10 ;
			data[39880] <= 8'h10 ;
			data[39881] <= 8'h10 ;
			data[39882] <= 8'h10 ;
			data[39883] <= 8'h10 ;
			data[39884] <= 8'h10 ;
			data[39885] <= 8'h10 ;
			data[39886] <= 8'h10 ;
			data[39887] <= 8'h10 ;
			data[39888] <= 8'h10 ;
			data[39889] <= 8'h10 ;
			data[39890] <= 8'h10 ;
			data[39891] <= 8'h10 ;
			data[39892] <= 8'h10 ;
			data[39893] <= 8'h10 ;
			data[39894] <= 8'h10 ;
			data[39895] <= 8'h10 ;
			data[39896] <= 8'h10 ;
			data[39897] <= 8'h10 ;
			data[39898] <= 8'h10 ;
			data[39899] <= 8'h10 ;
			data[39900] <= 8'h10 ;
			data[39901] <= 8'h10 ;
			data[39902] <= 8'h10 ;
			data[39903] <= 8'h10 ;
			data[39904] <= 8'h10 ;
			data[39905] <= 8'h10 ;
			data[39906] <= 8'h10 ;
			data[39907] <= 8'h10 ;
			data[39908] <= 8'h10 ;
			data[39909] <= 8'h10 ;
			data[39910] <= 8'h10 ;
			data[39911] <= 8'h10 ;
			data[39912] <= 8'h10 ;
			data[39913] <= 8'h10 ;
			data[39914] <= 8'h10 ;
			data[39915] <= 8'h10 ;
			data[39916] <= 8'h10 ;
			data[39917] <= 8'h10 ;
			data[39918] <= 8'h10 ;
			data[39919] <= 8'h10 ;
			data[39920] <= 8'h10 ;
			data[39921] <= 8'h10 ;
			data[39922] <= 8'h10 ;
			data[39923] <= 8'h10 ;
			data[39924] <= 8'h10 ;
			data[39925] <= 8'h10 ;
			data[39926] <= 8'h10 ;
			data[39927] <= 8'h10 ;
			data[39928] <= 8'h10 ;
			data[39929] <= 8'h10 ;
			data[39930] <= 8'h10 ;
			data[39931] <= 8'h10 ;
			data[39932] <= 8'h10 ;
			data[39933] <= 8'h10 ;
			data[39934] <= 8'h10 ;
			data[39935] <= 8'h10 ;
			data[39936] <= 8'h10 ;
			data[39937] <= 8'h10 ;
			data[39938] <= 8'h10 ;
			data[39939] <= 8'h10 ;
			data[39940] <= 8'h10 ;
			data[39941] <= 8'h10 ;
			data[39942] <= 8'h10 ;
			data[39943] <= 8'h10 ;
			data[39944] <= 8'h10 ;
			data[39945] <= 8'h10 ;
			data[39946] <= 8'h10 ;
			data[39947] <= 8'h10 ;
			data[39948] <= 8'h10 ;
			data[39949] <= 8'h10 ;
			data[39950] <= 8'h10 ;
			data[39951] <= 8'h10 ;
			data[39952] <= 8'h10 ;
			data[39953] <= 8'h10 ;
			data[39954] <= 8'h10 ;
			data[39955] <= 8'h10 ;
			data[39956] <= 8'h10 ;
			data[39957] <= 8'h10 ;
			data[39958] <= 8'h10 ;
			data[39959] <= 8'h10 ;
			data[39960] <= 8'h10 ;
			data[39961] <= 8'h10 ;
			data[39962] <= 8'h10 ;
			data[39963] <= 8'h10 ;
			data[39964] <= 8'h10 ;
			data[39965] <= 8'h10 ;
			data[39966] <= 8'h10 ;
			data[39967] <= 8'h10 ;
			data[39968] <= 8'h10 ;
			data[39969] <= 8'h10 ;
			data[39970] <= 8'h10 ;
			data[39971] <= 8'h10 ;
			data[39972] <= 8'h10 ;
			data[39973] <= 8'h10 ;
			data[39974] <= 8'h10 ;
			data[39975] <= 8'h10 ;
			data[39976] <= 8'h10 ;
			data[39977] <= 8'h10 ;
			data[39978] <= 8'h10 ;
			data[39979] <= 8'h10 ;
			data[39980] <= 8'h10 ;
			data[39981] <= 8'h10 ;
			data[39982] <= 8'h10 ;
			data[39983] <= 8'h10 ;
			data[39984] <= 8'h10 ;
			data[39985] <= 8'h10 ;
			data[39986] <= 8'h10 ;
			data[39987] <= 8'h10 ;
			data[39988] <= 8'h10 ;
			data[39989] <= 8'h10 ;
			data[39990] <= 8'h10 ;
			data[39991] <= 8'h10 ;
			data[39992] <= 8'h10 ;
			data[39993] <= 8'h10 ;
			data[39994] <= 8'h10 ;
			data[39995] <= 8'h10 ;
			data[39996] <= 8'h10 ;
			data[39997] <= 8'h10 ;
			data[39998] <= 8'h10 ;
			data[39999] <= 8'h10 ;
			data[40000] <= 8'h10 ;
			data[40001] <= 8'h10 ;
			data[40002] <= 8'h10 ;
			data[40003] <= 8'h10 ;
			data[40004] <= 8'h10 ;
			data[40005] <= 8'h10 ;
			data[40006] <= 8'h10 ;
			data[40007] <= 8'h10 ;
			data[40008] <= 8'h10 ;
			data[40009] <= 8'h10 ;
			data[40010] <= 8'h10 ;
			data[40011] <= 8'h10 ;
			data[40012] <= 8'h10 ;
			data[40013] <= 8'h10 ;
			data[40014] <= 8'h10 ;
			data[40015] <= 8'h10 ;
			data[40016] <= 8'h10 ;
			data[40017] <= 8'h10 ;
			data[40018] <= 8'h10 ;
			data[40019] <= 8'h10 ;
			data[40020] <= 8'h10 ;
			data[40021] <= 8'h10 ;
			data[40022] <= 8'h10 ;
			data[40023] <= 8'h10 ;
			data[40024] <= 8'h10 ;
			data[40025] <= 8'h10 ;
			data[40026] <= 8'h10 ;
			data[40027] <= 8'h10 ;
			data[40028] <= 8'h10 ;
			data[40029] <= 8'h10 ;
			data[40030] <= 8'h10 ;
			data[40031] <= 8'h10 ;
			data[40032] <= 8'h10 ;
			data[40033] <= 8'h10 ;
			data[40034] <= 8'h10 ;
			data[40035] <= 8'h10 ;
			data[40036] <= 8'h10 ;
			data[40037] <= 8'h10 ;
			data[40038] <= 8'h10 ;
			data[40039] <= 8'h10 ;
			data[40040] <= 8'h10 ;
			data[40041] <= 8'h10 ;
			data[40042] <= 8'h10 ;
			data[40043] <= 8'h10 ;
			data[40044] <= 8'h10 ;
			data[40045] <= 8'h10 ;
			data[40046] <= 8'h10 ;
			data[40047] <= 8'h10 ;
			data[40048] <= 8'h10 ;
			data[40049] <= 8'h10 ;
			data[40050] <= 8'h10 ;
			data[40051] <= 8'h10 ;
			data[40052] <= 8'h10 ;
			data[40053] <= 8'h10 ;
			data[40054] <= 8'h10 ;
			data[40055] <= 8'h10 ;
			data[40056] <= 8'h10 ;
			data[40057] <= 8'h10 ;
			data[40058] <= 8'h10 ;
			data[40059] <= 8'h10 ;
			data[40060] <= 8'h10 ;
			data[40061] <= 8'h10 ;
			data[40062] <= 8'h10 ;
			data[40063] <= 8'h10 ;
			data[40064] <= 8'h10 ;
			data[40065] <= 8'h10 ;
			data[40066] <= 8'h10 ;
			data[40067] <= 8'h10 ;
			data[40068] <= 8'h10 ;
			data[40069] <= 8'h10 ;
			data[40070] <= 8'h10 ;
			data[40071] <= 8'h10 ;
			data[40072] <= 8'h10 ;
			data[40073] <= 8'h10 ;
			data[40074] <= 8'h10 ;
			data[40075] <= 8'h10 ;
			data[40076] <= 8'h10 ;
			data[40077] <= 8'h10 ;
			data[40078] <= 8'h10 ;
			data[40079] <= 8'h10 ;
			data[40080] <= 8'h10 ;
			data[40081] <= 8'h10 ;
			data[40082] <= 8'h10 ;
			data[40083] <= 8'h10 ;
			data[40084] <= 8'h10 ;
			data[40085] <= 8'h10 ;
			data[40086] <= 8'h10 ;
			data[40087] <= 8'h10 ;
			data[40088] <= 8'h10 ;
			data[40089] <= 8'h10 ;
			data[40090] <= 8'h10 ;
			data[40091] <= 8'h10 ;
			data[40092] <= 8'h10 ;
			data[40093] <= 8'h10 ;
			data[40094] <= 8'h10 ;
			data[40095] <= 8'h10 ;
			data[40096] <= 8'h10 ;
			data[40097] <= 8'h10 ;
			data[40098] <= 8'h10 ;
			data[40099] <= 8'h10 ;
			data[40100] <= 8'h10 ;
			data[40101] <= 8'h10 ;
			data[40102] <= 8'h10 ;
			data[40103] <= 8'h10 ;
			data[40104] <= 8'h10 ;
			data[40105] <= 8'h10 ;
			data[40106] <= 8'h10 ;
			data[40107] <= 8'h10 ;
			data[40108] <= 8'h10 ;
			data[40109] <= 8'h10 ;
			data[40110] <= 8'h10 ;
			data[40111] <= 8'h10 ;
			data[40112] <= 8'h10 ;
			data[40113] <= 8'h10 ;
			data[40114] <= 8'h10 ;
			data[40115] <= 8'h10 ;
			data[40116] <= 8'h10 ;
			data[40117] <= 8'h10 ;
			data[40118] <= 8'h10 ;
			data[40119] <= 8'h10 ;
			data[40120] <= 8'h10 ;
			data[40121] <= 8'h10 ;
			data[40122] <= 8'h10 ;
			data[40123] <= 8'h10 ;
			data[40124] <= 8'h10 ;
			data[40125] <= 8'h10 ;
			data[40126] <= 8'h10 ;
			data[40127] <= 8'h10 ;
			data[40128] <= 8'h10 ;
			data[40129] <= 8'h10 ;
			data[40130] <= 8'h10 ;
			data[40131] <= 8'h10 ;
			data[40132] <= 8'h10 ;
			data[40133] <= 8'h10 ;
			data[40134] <= 8'h10 ;
			data[40135] <= 8'h10 ;
			data[40136] <= 8'h10 ;
			data[40137] <= 8'h10 ;
			data[40138] <= 8'h10 ;
			data[40139] <= 8'h10 ;
			data[40140] <= 8'h10 ;
			data[40141] <= 8'h10 ;
			data[40142] <= 8'h10 ;
			data[40143] <= 8'h10 ;
			data[40144] <= 8'h10 ;
			data[40145] <= 8'h10 ;
			data[40146] <= 8'h10 ;
			data[40147] <= 8'h10 ;
			data[40148] <= 8'h10 ;
			data[40149] <= 8'h10 ;
			data[40150] <= 8'h10 ;
			data[40151] <= 8'h10 ;
			data[40152] <= 8'h10 ;
			data[40153] <= 8'h10 ;
			data[40154] <= 8'h10 ;
			data[40155] <= 8'h10 ;
			data[40156] <= 8'h10 ;
			data[40157] <= 8'h10 ;
			data[40158] <= 8'h10 ;
			data[40159] <= 8'h10 ;
			data[40160] <= 8'h10 ;
			data[40161] <= 8'h10 ;
			data[40162] <= 8'h10 ;
			data[40163] <= 8'h10 ;
			data[40164] <= 8'h10 ;
			data[40165] <= 8'h10 ;
			data[40166] <= 8'h10 ;
			data[40167] <= 8'h10 ;
			data[40168] <= 8'h10 ;
			data[40169] <= 8'h10 ;
			data[40170] <= 8'h10 ;
			data[40171] <= 8'h10 ;
			data[40172] <= 8'h10 ;
			data[40173] <= 8'h10 ;
			data[40174] <= 8'h10 ;
			data[40175] <= 8'h10 ;
			data[40176] <= 8'h10 ;
			data[40177] <= 8'h10 ;
			data[40178] <= 8'h10 ;
			data[40179] <= 8'h10 ;
			data[40180] <= 8'h10 ;
			data[40181] <= 8'h10 ;
			data[40182] <= 8'h10 ;
			data[40183] <= 8'h10 ;
			data[40184] <= 8'h10 ;
			data[40185] <= 8'h10 ;
			data[40186] <= 8'h10 ;
			data[40187] <= 8'h10 ;
			data[40188] <= 8'h10 ;
			data[40189] <= 8'h10 ;
			data[40190] <= 8'h10 ;
			data[40191] <= 8'h10 ;
			data[40192] <= 8'h10 ;
			data[40193] <= 8'h10 ;
			data[40194] <= 8'h10 ;
			data[40195] <= 8'h10 ;
			data[40196] <= 8'h10 ;
			data[40197] <= 8'h10 ;
			data[40198] <= 8'h10 ;
			data[40199] <= 8'h10 ;
			data[40200] <= 8'h10 ;
			data[40201] <= 8'h10 ;
			data[40202] <= 8'h10 ;
			data[40203] <= 8'h10 ;
			data[40204] <= 8'h10 ;
			data[40205] <= 8'h10 ;
			data[40206] <= 8'h10 ;
			data[40207] <= 8'h10 ;
			data[40208] <= 8'h10 ;
			data[40209] <= 8'h10 ;
			data[40210] <= 8'h10 ;
			data[40211] <= 8'h10 ;
			data[40212] <= 8'h10 ;
			data[40213] <= 8'h10 ;
			data[40214] <= 8'h10 ;
			data[40215] <= 8'h10 ;
			data[40216] <= 8'h10 ;
			data[40217] <= 8'h10 ;
			data[40218] <= 8'h10 ;
			data[40219] <= 8'h10 ;
			data[40220] <= 8'h10 ;
			data[40221] <= 8'h10 ;
			data[40222] <= 8'h10 ;
			data[40223] <= 8'h10 ;
			data[40224] <= 8'h10 ;
			data[40225] <= 8'h10 ;
			data[40226] <= 8'h10 ;
			data[40227] <= 8'h10 ;
			data[40228] <= 8'h10 ;
			data[40229] <= 8'h10 ;
			data[40230] <= 8'h10 ;
			data[40231] <= 8'h10 ;
			data[40232] <= 8'h10 ;
			data[40233] <= 8'h10 ;
			data[40234] <= 8'h10 ;
			data[40235] <= 8'h10 ;
			data[40236] <= 8'h10 ;
			data[40237] <= 8'h10 ;
			data[40238] <= 8'h10 ;
			data[40239] <= 8'h10 ;
			data[40240] <= 8'h10 ;
			data[40241] <= 8'h10 ;
			data[40242] <= 8'h10 ;
			data[40243] <= 8'h10 ;
			data[40244] <= 8'h10 ;
			data[40245] <= 8'h10 ;
			data[40246] <= 8'h10 ;
			data[40247] <= 8'h10 ;
			data[40248] <= 8'h10 ;
			data[40249] <= 8'h10 ;
			data[40250] <= 8'h10 ;
			data[40251] <= 8'h10 ;
			data[40252] <= 8'h10 ;
			data[40253] <= 8'h10 ;
			data[40254] <= 8'h10 ;
			data[40255] <= 8'h10 ;
			data[40256] <= 8'h10 ;
			data[40257] <= 8'h10 ;
			data[40258] <= 8'h10 ;
			data[40259] <= 8'h10 ;
			data[40260] <= 8'h10 ;
			data[40261] <= 8'h10 ;
			data[40262] <= 8'h10 ;
			data[40263] <= 8'h10 ;
			data[40264] <= 8'h10 ;
			data[40265] <= 8'h10 ;
			data[40266] <= 8'h10 ;
			data[40267] <= 8'h10 ;
			data[40268] <= 8'h10 ;
			data[40269] <= 8'h10 ;
			data[40270] <= 8'h10 ;
			data[40271] <= 8'h10 ;
			data[40272] <= 8'h10 ;
			data[40273] <= 8'h10 ;
			data[40274] <= 8'h10 ;
			data[40275] <= 8'h10 ;
			data[40276] <= 8'h10 ;
			data[40277] <= 8'h10 ;
			data[40278] <= 8'h10 ;
			data[40279] <= 8'h10 ;
			data[40280] <= 8'h10 ;
			data[40281] <= 8'h10 ;
			data[40282] <= 8'h10 ;
			data[40283] <= 8'h10 ;
			data[40284] <= 8'h10 ;
			data[40285] <= 8'h10 ;
			data[40286] <= 8'h10 ;
			data[40287] <= 8'h10 ;
			data[40288] <= 8'h10 ;
			data[40289] <= 8'h10 ;
			data[40290] <= 8'h10 ;
			data[40291] <= 8'h10 ;
			data[40292] <= 8'h10 ;
			data[40293] <= 8'h10 ;
			data[40294] <= 8'h10 ;
			data[40295] <= 8'h10 ;
			data[40296] <= 8'h10 ;
			data[40297] <= 8'h10 ;
			data[40298] <= 8'h10 ;
			data[40299] <= 8'h10 ;
			data[40300] <= 8'h10 ;
			data[40301] <= 8'h10 ;
			data[40302] <= 8'h10 ;
			data[40303] <= 8'h10 ;
			data[40304] <= 8'h10 ;
			data[40305] <= 8'h10 ;
			data[40306] <= 8'h10 ;
			data[40307] <= 8'h10 ;
			data[40308] <= 8'h10 ;
			data[40309] <= 8'h10 ;
			data[40310] <= 8'h10 ;
			data[40311] <= 8'h10 ;
			data[40312] <= 8'h10 ;
			data[40313] <= 8'h10 ;
			data[40314] <= 8'h10 ;
			data[40315] <= 8'h10 ;
			data[40316] <= 8'h10 ;
			data[40317] <= 8'h10 ;
			data[40318] <= 8'h10 ;
			data[40319] <= 8'h10 ;
			data[40320] <= 8'h10 ;
			data[40321] <= 8'h10 ;
			data[40322] <= 8'h10 ;
			data[40323] <= 8'h10 ;
			data[40324] <= 8'h10 ;
			data[40325] <= 8'h10 ;
			data[40326] <= 8'h10 ;
			data[40327] <= 8'h10 ;
			data[40328] <= 8'h10 ;
			data[40329] <= 8'h10 ;
			data[40330] <= 8'h10 ;
			data[40331] <= 8'h10 ;
			data[40332] <= 8'h10 ;
			data[40333] <= 8'h10 ;
			data[40334] <= 8'h10 ;
			data[40335] <= 8'h10 ;
			data[40336] <= 8'h10 ;
			data[40337] <= 8'h10 ;
			data[40338] <= 8'h10 ;
			data[40339] <= 8'h10 ;
			data[40340] <= 8'h10 ;
			data[40341] <= 8'h10 ;
			data[40342] <= 8'h10 ;
			data[40343] <= 8'h10 ;
			data[40344] <= 8'h10 ;
			data[40345] <= 8'h10 ;
			data[40346] <= 8'h10 ;
			data[40347] <= 8'h10 ;
			data[40348] <= 8'h10 ;
			data[40349] <= 8'h10 ;
			data[40350] <= 8'h10 ;
			data[40351] <= 8'h10 ;
			data[40352] <= 8'h10 ;
			data[40353] <= 8'h10 ;
			data[40354] <= 8'h10 ;
			data[40355] <= 8'h10 ;
			data[40356] <= 8'h10 ;
			data[40357] <= 8'h10 ;
			data[40358] <= 8'h10 ;
			data[40359] <= 8'h10 ;
			data[40360] <= 8'h10 ;
			data[40361] <= 8'h10 ;
			data[40362] <= 8'h10 ;
			data[40363] <= 8'h10 ;
			data[40364] <= 8'h10 ;
			data[40365] <= 8'h10 ;
			data[40366] <= 8'h10 ;
			data[40367] <= 8'h10 ;
			data[40368] <= 8'h10 ;
			data[40369] <= 8'h10 ;
			data[40370] <= 8'h10 ;
			data[40371] <= 8'h10 ;
			data[40372] <= 8'h10 ;
			data[40373] <= 8'h10 ;
			data[40374] <= 8'h10 ;
			data[40375] <= 8'h10 ;
			data[40376] <= 8'h10 ;
			data[40377] <= 8'h10 ;
			data[40378] <= 8'h10 ;
			data[40379] <= 8'h10 ;
			data[40380] <= 8'h10 ;
			data[40381] <= 8'h10 ;
			data[40382] <= 8'h10 ;
			data[40383] <= 8'h10 ;
			data[40384] <= 8'h10 ;
			data[40385] <= 8'h10 ;
			data[40386] <= 8'h10 ;
			data[40387] <= 8'h10 ;
			data[40388] <= 8'h10 ;
			data[40389] <= 8'h10 ;
			data[40390] <= 8'h10 ;
			data[40391] <= 8'h10 ;
			data[40392] <= 8'h10 ;
			data[40393] <= 8'h10 ;
			data[40394] <= 8'h10 ;
			data[40395] <= 8'h10 ;
			data[40396] <= 8'h10 ;
			data[40397] <= 8'h10 ;
			data[40398] <= 8'h10 ;
			data[40399] <= 8'h10 ;
			data[40400] <= 8'h10 ;
			data[40401] <= 8'h10 ;
			data[40402] <= 8'h10 ;
			data[40403] <= 8'h10 ;
			data[40404] <= 8'h10 ;
			data[40405] <= 8'h10 ;
			data[40406] <= 8'h10 ;
			data[40407] <= 8'h10 ;
			data[40408] <= 8'h10 ;
			data[40409] <= 8'h10 ;
			data[40410] <= 8'h10 ;
			data[40411] <= 8'h10 ;
			data[40412] <= 8'h10 ;
			data[40413] <= 8'h10 ;
			data[40414] <= 8'h10 ;
			data[40415] <= 8'h10 ;
			data[40416] <= 8'h10 ;
			data[40417] <= 8'h10 ;
			data[40418] <= 8'h10 ;
			data[40419] <= 8'h10 ;
			data[40420] <= 8'h10 ;
			data[40421] <= 8'h10 ;
			data[40422] <= 8'h10 ;
			data[40423] <= 8'h10 ;
			data[40424] <= 8'h10 ;
			data[40425] <= 8'h10 ;
			data[40426] <= 8'h10 ;
			data[40427] <= 8'h10 ;
			data[40428] <= 8'h10 ;
			data[40429] <= 8'h10 ;
			data[40430] <= 8'h10 ;
			data[40431] <= 8'h10 ;
			data[40432] <= 8'h10 ;
			data[40433] <= 8'h10 ;
			data[40434] <= 8'h10 ;
			data[40435] <= 8'h10 ;
			data[40436] <= 8'h10 ;
			data[40437] <= 8'h10 ;
			data[40438] <= 8'h10 ;
			data[40439] <= 8'h10 ;
			data[40440] <= 8'h10 ;
			data[40441] <= 8'h10 ;
			data[40442] <= 8'h10 ;
			data[40443] <= 8'h10 ;
			data[40444] <= 8'h10 ;
			data[40445] <= 8'h10 ;
			data[40446] <= 8'h10 ;
			data[40447] <= 8'h10 ;
			data[40448] <= 8'h10 ;
			data[40449] <= 8'h10 ;
			data[40450] <= 8'h10 ;
			data[40451] <= 8'h10 ;
			data[40452] <= 8'h10 ;
			data[40453] <= 8'h10 ;
			data[40454] <= 8'h10 ;
			data[40455] <= 8'h10 ;
			data[40456] <= 8'h10 ;
			data[40457] <= 8'h10 ;
			data[40458] <= 8'h10 ;
			data[40459] <= 8'h10 ;
			data[40460] <= 8'h10 ;
			data[40461] <= 8'h10 ;
			data[40462] <= 8'h10 ;
			data[40463] <= 8'h10 ;
			data[40464] <= 8'h10 ;
			data[40465] <= 8'h10 ;
			data[40466] <= 8'h10 ;
			data[40467] <= 8'h10 ;
			data[40468] <= 8'h10 ;
			data[40469] <= 8'h10 ;
			data[40470] <= 8'h10 ;
			data[40471] <= 8'h10 ;
			data[40472] <= 8'h10 ;
			data[40473] <= 8'h10 ;
			data[40474] <= 8'h10 ;
			data[40475] <= 8'h10 ;
			data[40476] <= 8'h10 ;
			data[40477] <= 8'h10 ;
			data[40478] <= 8'h10 ;
			data[40479] <= 8'h10 ;
			data[40480] <= 8'h10 ;
			data[40481] <= 8'h10 ;
			data[40482] <= 8'h10 ;
			data[40483] <= 8'h10 ;
			data[40484] <= 8'h10 ;
			data[40485] <= 8'h10 ;
			data[40486] <= 8'h10 ;
			data[40487] <= 8'h10 ;
			data[40488] <= 8'h10 ;
			data[40489] <= 8'h10 ;
			data[40490] <= 8'h10 ;
			data[40491] <= 8'h10 ;
			data[40492] <= 8'h10 ;
			data[40493] <= 8'h10 ;
			data[40494] <= 8'h10 ;
			data[40495] <= 8'h10 ;
			data[40496] <= 8'h10 ;
			data[40497] <= 8'h10 ;
			data[40498] <= 8'h10 ;
			data[40499] <= 8'h10 ;
			data[40500] <= 8'h10 ;
			data[40501] <= 8'h10 ;
			data[40502] <= 8'h10 ;
			data[40503] <= 8'h10 ;
			data[40504] <= 8'h10 ;
			data[40505] <= 8'h10 ;
			data[40506] <= 8'h10 ;
			data[40507] <= 8'h10 ;
			data[40508] <= 8'h10 ;
			data[40509] <= 8'h10 ;
			data[40510] <= 8'h10 ;
			data[40511] <= 8'h10 ;
			data[40512] <= 8'h10 ;
			data[40513] <= 8'h10 ;
			data[40514] <= 8'h10 ;
			data[40515] <= 8'h10 ;
			data[40516] <= 8'h10 ;
			data[40517] <= 8'h10 ;
			data[40518] <= 8'h10 ;
			data[40519] <= 8'h10 ;
			data[40520] <= 8'h10 ;
			data[40521] <= 8'h10 ;
			data[40522] <= 8'h10 ;
			data[40523] <= 8'h10 ;
			data[40524] <= 8'h10 ;
			data[40525] <= 8'h10 ;
			data[40526] <= 8'h10 ;
			data[40527] <= 8'h10 ;
			data[40528] <= 8'h10 ;
			data[40529] <= 8'h10 ;
			data[40530] <= 8'h10 ;
			data[40531] <= 8'h10 ;
			data[40532] <= 8'h10 ;
			data[40533] <= 8'h10 ;
			data[40534] <= 8'h10 ;
			data[40535] <= 8'h10 ;
			data[40536] <= 8'h10 ;
			data[40537] <= 8'h10 ;
			data[40538] <= 8'h10 ;
			data[40539] <= 8'h10 ;
			data[40540] <= 8'h10 ;
			data[40541] <= 8'h10 ;
			data[40542] <= 8'h10 ;
			data[40543] <= 8'h10 ;
			data[40544] <= 8'h10 ;
			data[40545] <= 8'h10 ;
			data[40546] <= 8'h10 ;
			data[40547] <= 8'h10 ;
			data[40548] <= 8'h10 ;
			data[40549] <= 8'h10 ;
			data[40550] <= 8'h10 ;
			data[40551] <= 8'h10 ;
			data[40552] <= 8'h10 ;
			data[40553] <= 8'h10 ;
			data[40554] <= 8'h10 ;
			data[40555] <= 8'h10 ;
			data[40556] <= 8'h10 ;
			data[40557] <= 8'h10 ;
			data[40558] <= 8'h10 ;
			data[40559] <= 8'h10 ;
			data[40560] <= 8'h10 ;
			data[40561] <= 8'h10 ;
			data[40562] <= 8'h10 ;
			data[40563] <= 8'h10 ;
			data[40564] <= 8'h10 ;
			data[40565] <= 8'h10 ;
			data[40566] <= 8'h10 ;
			data[40567] <= 8'h10 ;
			data[40568] <= 8'h10 ;
			data[40569] <= 8'h10 ;
			data[40570] <= 8'h10 ;
			data[40571] <= 8'h10 ;
			data[40572] <= 8'h10 ;
			data[40573] <= 8'h10 ;
			data[40574] <= 8'h10 ;
			data[40575] <= 8'h10 ;
			data[40576] <= 8'h10 ;
			data[40577] <= 8'h10 ;
			data[40578] <= 8'h10 ;
			data[40579] <= 8'h10 ;
			data[40580] <= 8'h10 ;
			data[40581] <= 8'h10 ;
			data[40582] <= 8'h10 ;
			data[40583] <= 8'h10 ;
			data[40584] <= 8'h10 ;
			data[40585] <= 8'h10 ;
			data[40586] <= 8'h10 ;
			data[40587] <= 8'h10 ;
			data[40588] <= 8'h10 ;
			data[40589] <= 8'h10 ;
			data[40590] <= 8'h10 ;
			data[40591] <= 8'h10 ;
			data[40592] <= 8'h10 ;
			data[40593] <= 8'h10 ;
			data[40594] <= 8'h10 ;
			data[40595] <= 8'h10 ;
			data[40596] <= 8'h10 ;
			data[40597] <= 8'h10 ;
			data[40598] <= 8'h10 ;
			data[40599] <= 8'h10 ;
			data[40600] <= 8'h10 ;
			data[40601] <= 8'h10 ;
			data[40602] <= 8'h10 ;
			data[40603] <= 8'h10 ;
			data[40604] <= 8'h10 ;
			data[40605] <= 8'h10 ;
			data[40606] <= 8'h10 ;
			data[40607] <= 8'h10 ;
			data[40608] <= 8'h10 ;
			data[40609] <= 8'h10 ;
			data[40610] <= 8'h10 ;
			data[40611] <= 8'h10 ;
			data[40612] <= 8'h10 ;
			data[40613] <= 8'h10 ;
			data[40614] <= 8'h10 ;
			data[40615] <= 8'h10 ;
			data[40616] <= 8'h10 ;
			data[40617] <= 8'h10 ;
			data[40618] <= 8'h10 ;
			data[40619] <= 8'h10 ;
			data[40620] <= 8'h10 ;
			data[40621] <= 8'h10 ;
			data[40622] <= 8'h10 ;
			data[40623] <= 8'h10 ;
			data[40624] <= 8'h10 ;
			data[40625] <= 8'h10 ;
			data[40626] <= 8'h10 ;
			data[40627] <= 8'h10 ;
			data[40628] <= 8'h10 ;
			data[40629] <= 8'h10 ;
			data[40630] <= 8'h10 ;
			data[40631] <= 8'h10 ;
			data[40632] <= 8'h10 ;
			data[40633] <= 8'h10 ;
			data[40634] <= 8'h10 ;
			data[40635] <= 8'h10 ;
			data[40636] <= 8'h10 ;
			data[40637] <= 8'h10 ;
			data[40638] <= 8'h10 ;
			data[40639] <= 8'h10 ;
			data[40640] <= 8'h10 ;
			data[40641] <= 8'h10 ;
			data[40642] <= 8'h10 ;
			data[40643] <= 8'h10 ;
			data[40644] <= 8'h10 ;
			data[40645] <= 8'h10 ;
			data[40646] <= 8'h10 ;
			data[40647] <= 8'h10 ;
			data[40648] <= 8'h10 ;
			data[40649] <= 8'h10 ;
			data[40650] <= 8'h10 ;
			data[40651] <= 8'h10 ;
			data[40652] <= 8'h10 ;
			data[40653] <= 8'h10 ;
			data[40654] <= 8'h10 ;
			data[40655] <= 8'h10 ;
			data[40656] <= 8'h10 ;
			data[40657] <= 8'h10 ;
			data[40658] <= 8'h10 ;
			data[40659] <= 8'h10 ;
			data[40660] <= 8'h10 ;
			data[40661] <= 8'h10 ;
			data[40662] <= 8'h10 ;
			data[40663] <= 8'h10 ;
			data[40664] <= 8'h10 ;
			data[40665] <= 8'h10 ;
			data[40666] <= 8'h10 ;
			data[40667] <= 8'h10 ;
			data[40668] <= 8'h10 ;
			data[40669] <= 8'h10 ;
			data[40670] <= 8'h10 ;
			data[40671] <= 8'h10 ;
			data[40672] <= 8'h10 ;
			data[40673] <= 8'h10 ;
			data[40674] <= 8'h10 ;
			data[40675] <= 8'h10 ;
			data[40676] <= 8'h10 ;
			data[40677] <= 8'h10 ;
			data[40678] <= 8'h10 ;
			data[40679] <= 8'h10 ;
			data[40680] <= 8'h10 ;
			data[40681] <= 8'h10 ;
			data[40682] <= 8'h10 ;
			data[40683] <= 8'h10 ;
			data[40684] <= 8'h10 ;
			data[40685] <= 8'h10 ;
			data[40686] <= 8'h10 ;
			data[40687] <= 8'h10 ;
			data[40688] <= 8'h10 ;
			data[40689] <= 8'h10 ;
			data[40690] <= 8'h10 ;
			data[40691] <= 8'h10 ;
			data[40692] <= 8'h10 ;
			data[40693] <= 8'h10 ;
			data[40694] <= 8'h10 ;
			data[40695] <= 8'h10 ;
			data[40696] <= 8'h10 ;
			data[40697] <= 8'h10 ;
			data[40698] <= 8'h10 ;
			data[40699] <= 8'h10 ;
			data[40700] <= 8'h10 ;
			data[40701] <= 8'h10 ;
			data[40702] <= 8'h10 ;
			data[40703] <= 8'h10 ;
			data[40704] <= 8'h10 ;
			data[40705] <= 8'h10 ;
			data[40706] <= 8'h10 ;
			data[40707] <= 8'h10 ;
			data[40708] <= 8'h10 ;
			data[40709] <= 8'h10 ;
			data[40710] <= 8'h10 ;
			data[40711] <= 8'h10 ;
			data[40712] <= 8'h10 ;
			data[40713] <= 8'h10 ;
			data[40714] <= 8'h10 ;
			data[40715] <= 8'h10 ;
			data[40716] <= 8'h10 ;
			data[40717] <= 8'h10 ;
			data[40718] <= 8'h10 ;
			data[40719] <= 8'h10 ;
			data[40720] <= 8'h10 ;
			data[40721] <= 8'h10 ;
			data[40722] <= 8'h10 ;
			data[40723] <= 8'h10 ;
			data[40724] <= 8'h10 ;
			data[40725] <= 8'h10 ;
			data[40726] <= 8'h10 ;
			data[40727] <= 8'h10 ;
			data[40728] <= 8'h10 ;
			data[40729] <= 8'h10 ;
			data[40730] <= 8'h10 ;
			data[40731] <= 8'h10 ;
			data[40732] <= 8'h10 ;
			data[40733] <= 8'h10 ;
			data[40734] <= 8'h10 ;
			data[40735] <= 8'h10 ;
			data[40736] <= 8'h10 ;
			data[40737] <= 8'h10 ;
			data[40738] <= 8'h10 ;
			data[40739] <= 8'h10 ;
			data[40740] <= 8'h10 ;
			data[40741] <= 8'h10 ;
			data[40742] <= 8'h10 ;
			data[40743] <= 8'h10 ;
			data[40744] <= 8'h10 ;
			data[40745] <= 8'h10 ;
			data[40746] <= 8'h10 ;
			data[40747] <= 8'h10 ;
			data[40748] <= 8'h10 ;
			data[40749] <= 8'h10 ;
			data[40750] <= 8'h10 ;
			data[40751] <= 8'h10 ;
			data[40752] <= 8'h10 ;
			data[40753] <= 8'h10 ;
			data[40754] <= 8'h10 ;
			data[40755] <= 8'h10 ;
			data[40756] <= 8'h10 ;
			data[40757] <= 8'h10 ;
			data[40758] <= 8'h10 ;
			data[40759] <= 8'h10 ;
			data[40760] <= 8'h10 ;
			data[40761] <= 8'h10 ;
			data[40762] <= 8'h10 ;
			data[40763] <= 8'h10 ;
			data[40764] <= 8'h10 ;
			data[40765] <= 8'h10 ;
			data[40766] <= 8'h10 ;
			data[40767] <= 8'h10 ;
			data[40768] <= 8'h10 ;
			data[40769] <= 8'h10 ;
			data[40770] <= 8'h10 ;
			data[40771] <= 8'h10 ;
			data[40772] <= 8'h10 ;
			data[40773] <= 8'h10 ;
			data[40774] <= 8'h10 ;
			data[40775] <= 8'h10 ;
			data[40776] <= 8'h10 ;
			data[40777] <= 8'h10 ;
			data[40778] <= 8'h10 ;
			data[40779] <= 8'h10 ;
			data[40780] <= 8'h10 ;
			data[40781] <= 8'h10 ;
			data[40782] <= 8'h10 ;
			data[40783] <= 8'h10 ;
			data[40784] <= 8'h10 ;
			data[40785] <= 8'h10 ;
			data[40786] <= 8'h10 ;
			data[40787] <= 8'h10 ;
			data[40788] <= 8'h10 ;
			data[40789] <= 8'h10 ;
			data[40790] <= 8'h10 ;
			data[40791] <= 8'h10 ;
			data[40792] <= 8'h10 ;
			data[40793] <= 8'h10 ;
			data[40794] <= 8'h10 ;
			data[40795] <= 8'h10 ;
			data[40796] <= 8'h10 ;
			data[40797] <= 8'h10 ;
			data[40798] <= 8'h10 ;
			data[40799] <= 8'h10 ;
			data[40800] <= 8'h10 ;
			data[40801] <= 8'h10 ;
			data[40802] <= 8'h10 ;
			data[40803] <= 8'h10 ;
			data[40804] <= 8'h10 ;
			data[40805] <= 8'h10 ;
			data[40806] <= 8'h10 ;
			data[40807] <= 8'h10 ;
			data[40808] <= 8'h10 ;
			data[40809] <= 8'h10 ;
			data[40810] <= 8'h10 ;
			data[40811] <= 8'h10 ;
			data[40812] <= 8'h10 ;
			data[40813] <= 8'h10 ;
			data[40814] <= 8'h10 ;
			data[40815] <= 8'h10 ;
			data[40816] <= 8'h10 ;
			data[40817] <= 8'h10 ;
			data[40818] <= 8'h10 ;
			data[40819] <= 8'h10 ;
			data[40820] <= 8'h10 ;
			data[40821] <= 8'h10 ;
			data[40822] <= 8'h10 ;
			data[40823] <= 8'h10 ;
			data[40824] <= 8'h10 ;
			data[40825] <= 8'h10 ;
			data[40826] <= 8'h10 ;
			data[40827] <= 8'h10 ;
			data[40828] <= 8'h10 ;
			data[40829] <= 8'h10 ;
			data[40830] <= 8'h10 ;
			data[40831] <= 8'h10 ;
			data[40832] <= 8'h10 ;
			data[40833] <= 8'h10 ;
			data[40834] <= 8'h10 ;
			data[40835] <= 8'h10 ;
			data[40836] <= 8'h10 ;
			data[40837] <= 8'h10 ;
			data[40838] <= 8'h10 ;
			data[40839] <= 8'h10 ;
			data[40840] <= 8'h10 ;
			data[40841] <= 8'h10 ;
			data[40842] <= 8'h10 ;
			data[40843] <= 8'h10 ;
			data[40844] <= 8'h10 ;
			data[40845] <= 8'h10 ;
			data[40846] <= 8'h10 ;
			data[40847] <= 8'h10 ;
			data[40848] <= 8'h10 ;
			data[40849] <= 8'h10 ;
			data[40850] <= 8'h10 ;
			data[40851] <= 8'h10 ;
			data[40852] <= 8'h10 ;
			data[40853] <= 8'h10 ;
			data[40854] <= 8'h10 ;
			data[40855] <= 8'h10 ;
			data[40856] <= 8'h10 ;
			data[40857] <= 8'h10 ;
			data[40858] <= 8'h10 ;
			data[40859] <= 8'h10 ;
			data[40860] <= 8'h10 ;
			data[40861] <= 8'h10 ;
			data[40862] <= 8'h10 ;
			data[40863] <= 8'h10 ;
			data[40864] <= 8'h10 ;
			data[40865] <= 8'h10 ;
			data[40866] <= 8'h10 ;
			data[40867] <= 8'h10 ;
			data[40868] <= 8'h10 ;
			data[40869] <= 8'h10 ;
			data[40870] <= 8'h10 ;
			data[40871] <= 8'h10 ;
			data[40872] <= 8'h10 ;
			data[40873] <= 8'h10 ;
			data[40874] <= 8'h10 ;
			data[40875] <= 8'h10 ;
			data[40876] <= 8'h10 ;
			data[40877] <= 8'h10 ;
			data[40878] <= 8'h10 ;
			data[40879] <= 8'h10 ;
			data[40880] <= 8'h10 ;
			data[40881] <= 8'h10 ;
			data[40882] <= 8'h10 ;
			data[40883] <= 8'h10 ;
			data[40884] <= 8'h10 ;
			data[40885] <= 8'h10 ;
			data[40886] <= 8'h10 ;
			data[40887] <= 8'h10 ;
			data[40888] <= 8'h10 ;
			data[40889] <= 8'h10 ;
			data[40890] <= 8'h10 ;
			data[40891] <= 8'h10 ;
			data[40892] <= 8'h10 ;
			data[40893] <= 8'h10 ;
			data[40894] <= 8'h10 ;
			data[40895] <= 8'h10 ;
			data[40896] <= 8'h10 ;
			data[40897] <= 8'h10 ;
			data[40898] <= 8'h10 ;
			data[40899] <= 8'h10 ;
			data[40900] <= 8'h10 ;
			data[40901] <= 8'h10 ;
			data[40902] <= 8'h10 ;
			data[40903] <= 8'h10 ;
			data[40904] <= 8'h10 ;
			data[40905] <= 8'h10 ;
			data[40906] <= 8'h10 ;
			data[40907] <= 8'h10 ;
			data[40908] <= 8'h10 ;
			data[40909] <= 8'h10 ;
			data[40910] <= 8'h10 ;
			data[40911] <= 8'h10 ;
			data[40912] <= 8'h10 ;
			data[40913] <= 8'h10 ;
			data[40914] <= 8'h10 ;
			data[40915] <= 8'h10 ;
			data[40916] <= 8'h10 ;
			data[40917] <= 8'h10 ;
			data[40918] <= 8'h10 ;
			data[40919] <= 8'h10 ;
			data[40920] <= 8'h10 ;
			data[40921] <= 8'h10 ;
			data[40922] <= 8'h10 ;
			data[40923] <= 8'h10 ;
			data[40924] <= 8'h10 ;
			data[40925] <= 8'h10 ;
			data[40926] <= 8'h10 ;
			data[40927] <= 8'h10 ;
			data[40928] <= 8'h10 ;
			data[40929] <= 8'h10 ;
			data[40930] <= 8'h10 ;
			data[40931] <= 8'h10 ;
			data[40932] <= 8'h10 ;
			data[40933] <= 8'h10 ;
			data[40934] <= 8'h10 ;
			data[40935] <= 8'h10 ;
			data[40936] <= 8'h10 ;
			data[40937] <= 8'h10 ;
			data[40938] <= 8'h10 ;
			data[40939] <= 8'h10 ;
			data[40940] <= 8'h10 ;
			data[40941] <= 8'h10 ;
			data[40942] <= 8'h10 ;
			data[40943] <= 8'h10 ;
			data[40944] <= 8'h10 ;
			data[40945] <= 8'h10 ;
			data[40946] <= 8'h10 ;
			data[40947] <= 8'h10 ;
			data[40948] <= 8'h10 ;
			data[40949] <= 8'h10 ;
			data[40950] <= 8'h10 ;
			data[40951] <= 8'h10 ;
			data[40952] <= 8'h10 ;
			data[40953] <= 8'h10 ;
			data[40954] <= 8'h10 ;
			data[40955] <= 8'h10 ;
			data[40956] <= 8'h10 ;
			data[40957] <= 8'h10 ;
			data[40958] <= 8'h10 ;
			data[40959] <= 8'h10 ;
			data[40960] <= 8'h10 ;
			data[40961] <= 8'h10 ;
			data[40962] <= 8'h10 ;
			data[40963] <= 8'h10 ;
			data[40964] <= 8'h10 ;
			data[40965] <= 8'h10 ;
			data[40966] <= 8'h10 ;
			data[40967] <= 8'h10 ;
			data[40968] <= 8'h10 ;
			data[40969] <= 8'h10 ;
			data[40970] <= 8'h10 ;
			data[40971] <= 8'h10 ;
			data[40972] <= 8'h10 ;
			data[40973] <= 8'h10 ;
			data[40974] <= 8'h10 ;
			data[40975] <= 8'h10 ;
			data[40976] <= 8'h10 ;
			data[40977] <= 8'h10 ;
			data[40978] <= 8'h10 ;
			data[40979] <= 8'h10 ;
			data[40980] <= 8'h10 ;
			data[40981] <= 8'h10 ;
			data[40982] <= 8'h10 ;
			data[40983] <= 8'h10 ;
			data[40984] <= 8'h10 ;
			data[40985] <= 8'h10 ;
			data[40986] <= 8'h10 ;
			data[40987] <= 8'h10 ;
			data[40988] <= 8'h10 ;
			data[40989] <= 8'h10 ;
			data[40990] <= 8'h10 ;
			data[40991] <= 8'h10 ;
			data[40992] <= 8'h10 ;
			data[40993] <= 8'h10 ;
			data[40994] <= 8'h10 ;
			data[40995] <= 8'h10 ;
			data[40996] <= 8'h10 ;
			data[40997] <= 8'h10 ;
			data[40998] <= 8'h10 ;
			data[40999] <= 8'h10 ;
			data[41000] <= 8'h10 ;
			data[41001] <= 8'h10 ;
			data[41002] <= 8'h10 ;
			data[41003] <= 8'h10 ;
			data[41004] <= 8'h10 ;
			data[41005] <= 8'h10 ;
			data[41006] <= 8'h10 ;
			data[41007] <= 8'h10 ;
			data[41008] <= 8'h10 ;
			data[41009] <= 8'h10 ;
			data[41010] <= 8'h10 ;
			data[41011] <= 8'h10 ;
			data[41012] <= 8'h10 ;
			data[41013] <= 8'h10 ;
			data[41014] <= 8'h10 ;
			data[41015] <= 8'h10 ;
			data[41016] <= 8'h10 ;
			data[41017] <= 8'h10 ;
			data[41018] <= 8'h10 ;
			data[41019] <= 8'h10 ;
			data[41020] <= 8'h10 ;
			data[41021] <= 8'h10 ;
			data[41022] <= 8'h10 ;
			data[41023] <= 8'h10 ;
			data[41024] <= 8'h10 ;
			data[41025] <= 8'h10 ;
			data[41026] <= 8'h10 ;
			data[41027] <= 8'h10 ;
			data[41028] <= 8'h10 ;
			data[41029] <= 8'h10 ;
			data[41030] <= 8'h10 ;
			data[41031] <= 8'h10 ;
			data[41032] <= 8'h10 ;
			data[41033] <= 8'h10 ;
			data[41034] <= 8'h10 ;
			data[41035] <= 8'h10 ;
			data[41036] <= 8'h10 ;
			data[41037] <= 8'h10 ;
			data[41038] <= 8'h10 ;
			data[41039] <= 8'h10 ;
			data[41040] <= 8'h10 ;
			data[41041] <= 8'h10 ;
			data[41042] <= 8'h10 ;
			data[41043] <= 8'h10 ;
			data[41044] <= 8'h10 ;
			data[41045] <= 8'h10 ;
			data[41046] <= 8'h10 ;
			data[41047] <= 8'h10 ;
			data[41048] <= 8'h10 ;
			data[41049] <= 8'h10 ;
			data[41050] <= 8'h10 ;
			data[41051] <= 8'h10 ;
			data[41052] <= 8'h10 ;
			data[41053] <= 8'h10 ;
			data[41054] <= 8'h10 ;
			data[41055] <= 8'h10 ;
			data[41056] <= 8'h10 ;
			data[41057] <= 8'h10 ;
			data[41058] <= 8'h10 ;
			data[41059] <= 8'h10 ;
			data[41060] <= 8'h10 ;
			data[41061] <= 8'h10 ;
			data[41062] <= 8'h10 ;
			data[41063] <= 8'h10 ;
			data[41064] <= 8'h10 ;
			data[41065] <= 8'h10 ;
			data[41066] <= 8'h10 ;
			data[41067] <= 8'h10 ;
			data[41068] <= 8'h10 ;
			data[41069] <= 8'h10 ;
			data[41070] <= 8'h10 ;
			data[41071] <= 8'h10 ;
			data[41072] <= 8'h10 ;
			data[41073] <= 8'h10 ;
			data[41074] <= 8'h10 ;
			data[41075] <= 8'h10 ;
			data[41076] <= 8'h10 ;
			data[41077] <= 8'h10 ;
			data[41078] <= 8'h10 ;
			data[41079] <= 8'h10 ;
			data[41080] <= 8'h10 ;
			data[41081] <= 8'h10 ;
			data[41082] <= 8'h10 ;
			data[41083] <= 8'h10 ;
			data[41084] <= 8'h10 ;
			data[41085] <= 8'h10 ;
			data[41086] <= 8'h10 ;
			data[41087] <= 8'h10 ;
			data[41088] <= 8'h10 ;
			data[41089] <= 8'h10 ;
			data[41090] <= 8'h10 ;
			data[41091] <= 8'h10 ;
			data[41092] <= 8'h10 ;
			data[41093] <= 8'h10 ;
			data[41094] <= 8'h10 ;
			data[41095] <= 8'h10 ;
			data[41096] <= 8'h10 ;
			data[41097] <= 8'h10 ;
			data[41098] <= 8'h10 ;
			data[41099] <= 8'h10 ;
			data[41100] <= 8'h10 ;
			data[41101] <= 8'h10 ;
			data[41102] <= 8'h10 ;
			data[41103] <= 8'h10 ;
			data[41104] <= 8'h10 ;
			data[41105] <= 8'h10 ;
			data[41106] <= 8'h10 ;
			data[41107] <= 8'h10 ;
			data[41108] <= 8'h10 ;
			data[41109] <= 8'h10 ;
			data[41110] <= 8'h10 ;
			data[41111] <= 8'h10 ;
			data[41112] <= 8'h10 ;
			data[41113] <= 8'h10 ;
			data[41114] <= 8'h10 ;
			data[41115] <= 8'h10 ;
			data[41116] <= 8'h10 ;
			data[41117] <= 8'h10 ;
			data[41118] <= 8'h10 ;
			data[41119] <= 8'h10 ;
			data[41120] <= 8'h10 ;
			data[41121] <= 8'h10 ;
			data[41122] <= 8'h10 ;
			data[41123] <= 8'h10 ;
			data[41124] <= 8'h10 ;
			data[41125] <= 8'h10 ;
			data[41126] <= 8'h10 ;
			data[41127] <= 8'h10 ;
			data[41128] <= 8'h10 ;
			data[41129] <= 8'h10 ;
			data[41130] <= 8'h10 ;
			data[41131] <= 8'h10 ;
			data[41132] <= 8'h10 ;
			data[41133] <= 8'h10 ;
			data[41134] <= 8'h10 ;
			data[41135] <= 8'h10 ;
			data[41136] <= 8'h10 ;
			data[41137] <= 8'h10 ;
			data[41138] <= 8'h10 ;
			data[41139] <= 8'h10 ;
			data[41140] <= 8'h10 ;
			data[41141] <= 8'h10 ;
			data[41142] <= 8'h10 ;
			data[41143] <= 8'h10 ;
			data[41144] <= 8'h10 ;
			data[41145] <= 8'h10 ;
			data[41146] <= 8'h10 ;
			data[41147] <= 8'h10 ;
			data[41148] <= 8'h10 ;
			data[41149] <= 8'h10 ;
			data[41150] <= 8'h10 ;
			data[41151] <= 8'h10 ;
			data[41152] <= 8'h10 ;
			data[41153] <= 8'h10 ;
			data[41154] <= 8'h10 ;
			data[41155] <= 8'h10 ;
			data[41156] <= 8'h10 ;
			data[41157] <= 8'h10 ;
			data[41158] <= 8'h10 ;
			data[41159] <= 8'h10 ;
			data[41160] <= 8'h10 ;
			data[41161] <= 8'h10 ;
			data[41162] <= 8'h10 ;
			data[41163] <= 8'h10 ;
			data[41164] <= 8'h10 ;
			data[41165] <= 8'h10 ;
			data[41166] <= 8'h10 ;
			data[41167] <= 8'h10 ;
			data[41168] <= 8'h10 ;
			data[41169] <= 8'h10 ;
			data[41170] <= 8'h10 ;
			data[41171] <= 8'h10 ;
			data[41172] <= 8'h10 ;
			data[41173] <= 8'h10 ;
			data[41174] <= 8'h10 ;
			data[41175] <= 8'h10 ;
			data[41176] <= 8'h10 ;
			data[41177] <= 8'h10 ;
			data[41178] <= 8'h10 ;
			data[41179] <= 8'h10 ;
			data[41180] <= 8'h10 ;
			data[41181] <= 8'h10 ;
			data[41182] <= 8'h10 ;
			data[41183] <= 8'h10 ;
			data[41184] <= 8'h10 ;
			data[41185] <= 8'h10 ;
			data[41186] <= 8'h10 ;
			data[41187] <= 8'h10 ;
			data[41188] <= 8'h10 ;
			data[41189] <= 8'h10 ;
			data[41190] <= 8'h10 ;
			data[41191] <= 8'h10 ;
			data[41192] <= 8'h10 ;
			data[41193] <= 8'h10 ;
			data[41194] <= 8'h10 ;
			data[41195] <= 8'h10 ;
			data[41196] <= 8'h10 ;
			data[41197] <= 8'h10 ;
			data[41198] <= 8'h10 ;
			data[41199] <= 8'h10 ;
			data[41200] <= 8'h10 ;
			data[41201] <= 8'h10 ;
			data[41202] <= 8'h10 ;
			data[41203] <= 8'h10 ;
			data[41204] <= 8'h10 ;
			data[41205] <= 8'h10 ;
			data[41206] <= 8'h10 ;
			data[41207] <= 8'h10 ;
			data[41208] <= 8'h10 ;
			data[41209] <= 8'h10 ;
			data[41210] <= 8'h10 ;
			data[41211] <= 8'h10 ;
			data[41212] <= 8'h10 ;
			data[41213] <= 8'h10 ;
			data[41214] <= 8'h10 ;
			data[41215] <= 8'h10 ;
			data[41216] <= 8'h10 ;
			data[41217] <= 8'h10 ;
			data[41218] <= 8'h10 ;
			data[41219] <= 8'h10 ;
			data[41220] <= 8'h10 ;
			data[41221] <= 8'h10 ;
			data[41222] <= 8'h10 ;
			data[41223] <= 8'h10 ;
			data[41224] <= 8'h10 ;
			data[41225] <= 8'h10 ;
			data[41226] <= 8'h10 ;
			data[41227] <= 8'h10 ;
			data[41228] <= 8'h10 ;
			data[41229] <= 8'h10 ;
			data[41230] <= 8'h10 ;
			data[41231] <= 8'h10 ;
			data[41232] <= 8'h10 ;
			data[41233] <= 8'h10 ;
			data[41234] <= 8'h10 ;
			data[41235] <= 8'h10 ;
			data[41236] <= 8'h10 ;
			data[41237] <= 8'h10 ;
			data[41238] <= 8'h10 ;
			data[41239] <= 8'h10 ;
			data[41240] <= 8'h10 ;
			data[41241] <= 8'h10 ;
			data[41242] <= 8'h10 ;
			data[41243] <= 8'h10 ;
			data[41244] <= 8'h10 ;
			data[41245] <= 8'h10 ;
			data[41246] <= 8'h10 ;
			data[41247] <= 8'h10 ;
			data[41248] <= 8'h10 ;
			data[41249] <= 8'h10 ;
			data[41250] <= 8'h10 ;
			data[41251] <= 8'h10 ;
			data[41252] <= 8'h10 ;
			data[41253] <= 8'h10 ;
			data[41254] <= 8'h10 ;
			data[41255] <= 8'h10 ;
			data[41256] <= 8'h10 ;
			data[41257] <= 8'h10 ;
			data[41258] <= 8'h10 ;
			data[41259] <= 8'h10 ;
			data[41260] <= 8'h10 ;
			data[41261] <= 8'h10 ;
			data[41262] <= 8'h10 ;
			data[41263] <= 8'h10 ;
			data[41264] <= 8'h10 ;
			data[41265] <= 8'h10 ;
			data[41266] <= 8'h10 ;
			data[41267] <= 8'h10 ;
			data[41268] <= 8'h10 ;
			data[41269] <= 8'h10 ;
			data[41270] <= 8'h10 ;
			data[41271] <= 8'h10 ;
			data[41272] <= 8'h10 ;
			data[41273] <= 8'h10 ;
			data[41274] <= 8'h10 ;
			data[41275] <= 8'h10 ;
			data[41276] <= 8'h10 ;
			data[41277] <= 8'h10 ;
			data[41278] <= 8'h10 ;
			data[41279] <= 8'h10 ;
			data[41280] <= 8'h10 ;
			data[41281] <= 8'h10 ;
			data[41282] <= 8'h10 ;
			data[41283] <= 8'h10 ;
			data[41284] <= 8'h10 ;
			data[41285] <= 8'h10 ;
			data[41286] <= 8'h10 ;
			data[41287] <= 8'h10 ;
			data[41288] <= 8'h10 ;
			data[41289] <= 8'h10 ;
			data[41290] <= 8'h10 ;
			data[41291] <= 8'h10 ;
			data[41292] <= 8'h10 ;
			data[41293] <= 8'h10 ;
			data[41294] <= 8'h10 ;
			data[41295] <= 8'h10 ;
			data[41296] <= 8'h10 ;
			data[41297] <= 8'h10 ;
			data[41298] <= 8'h10 ;
			data[41299] <= 8'h10 ;
			data[41300] <= 8'h10 ;
			data[41301] <= 8'h10 ;
			data[41302] <= 8'h10 ;
			data[41303] <= 8'h10 ;
			data[41304] <= 8'h10 ;
			data[41305] <= 8'h10 ;
			data[41306] <= 8'h10 ;
			data[41307] <= 8'h10 ;
			data[41308] <= 8'h10 ;
			data[41309] <= 8'h10 ;
			data[41310] <= 8'h10 ;
			data[41311] <= 8'h10 ;
			data[41312] <= 8'h10 ;
			data[41313] <= 8'h10 ;
			data[41314] <= 8'h10 ;
			data[41315] <= 8'h10 ;
			data[41316] <= 8'h10 ;
			data[41317] <= 8'h10 ;
			data[41318] <= 8'h10 ;
			data[41319] <= 8'h10 ;
			data[41320] <= 8'h10 ;
			data[41321] <= 8'h10 ;
			data[41322] <= 8'h10 ;
			data[41323] <= 8'h10 ;
			data[41324] <= 8'h10 ;
			data[41325] <= 8'h10 ;
			data[41326] <= 8'h10 ;
			data[41327] <= 8'h10 ;
			data[41328] <= 8'h10 ;
			data[41329] <= 8'h10 ;
			data[41330] <= 8'h10 ;
			data[41331] <= 8'h10 ;
			data[41332] <= 8'h10 ;
			data[41333] <= 8'h10 ;
			data[41334] <= 8'h10 ;
			data[41335] <= 8'h10 ;
			data[41336] <= 8'h10 ;
			data[41337] <= 8'h10 ;
			data[41338] <= 8'h10 ;
			data[41339] <= 8'h10 ;
			data[41340] <= 8'h10 ;
			data[41341] <= 8'h10 ;
			data[41342] <= 8'h10 ;
			data[41343] <= 8'h10 ;
			data[41344] <= 8'h10 ;
			data[41345] <= 8'h10 ;
			data[41346] <= 8'h10 ;
			data[41347] <= 8'h10 ;
			data[41348] <= 8'h10 ;
			data[41349] <= 8'h10 ;
			data[41350] <= 8'h10 ;
			data[41351] <= 8'h10 ;
			data[41352] <= 8'h10 ;
			data[41353] <= 8'h10 ;
			data[41354] <= 8'h10 ;
			data[41355] <= 8'h10 ;
			data[41356] <= 8'h10 ;
			data[41357] <= 8'h10 ;
			data[41358] <= 8'h10 ;
			data[41359] <= 8'h10 ;
			data[41360] <= 8'h10 ;
			data[41361] <= 8'h10 ;
			data[41362] <= 8'h10 ;
			data[41363] <= 8'h10 ;
			data[41364] <= 8'h10 ;
			data[41365] <= 8'h10 ;
			data[41366] <= 8'h10 ;
			data[41367] <= 8'h10 ;
			data[41368] <= 8'h10 ;
			data[41369] <= 8'h10 ;
			data[41370] <= 8'h10 ;
			data[41371] <= 8'h10 ;
			data[41372] <= 8'h10 ;
			data[41373] <= 8'h10 ;
			data[41374] <= 8'h10 ;
			data[41375] <= 8'h10 ;
			data[41376] <= 8'h10 ;
			data[41377] <= 8'h10 ;
			data[41378] <= 8'h10 ;
			data[41379] <= 8'h10 ;
			data[41380] <= 8'h10 ;
			data[41381] <= 8'h10 ;
			data[41382] <= 8'h10 ;
			data[41383] <= 8'h10 ;
			data[41384] <= 8'h10 ;
			data[41385] <= 8'h10 ;
			data[41386] <= 8'h10 ;
			data[41387] <= 8'h10 ;
			data[41388] <= 8'h10 ;
			data[41389] <= 8'h10 ;
			data[41390] <= 8'h10 ;
			data[41391] <= 8'h10 ;
			data[41392] <= 8'h10 ;
			data[41393] <= 8'h10 ;
			data[41394] <= 8'h10 ;
			data[41395] <= 8'h10 ;
			data[41396] <= 8'h10 ;
			data[41397] <= 8'h10 ;
			data[41398] <= 8'h10 ;
			data[41399] <= 8'h10 ;
			data[41400] <= 8'h10 ;
			data[41401] <= 8'h10 ;
			data[41402] <= 8'h10 ;
			data[41403] <= 8'h10 ;
			data[41404] <= 8'h10 ;
			data[41405] <= 8'h10 ;
			data[41406] <= 8'h10 ;
			data[41407] <= 8'h10 ;
			data[41408] <= 8'h10 ;
			data[41409] <= 8'h10 ;
			data[41410] <= 8'h10 ;
			data[41411] <= 8'h10 ;
			data[41412] <= 8'h10 ;
			data[41413] <= 8'h10 ;
			data[41414] <= 8'h10 ;
			data[41415] <= 8'h10 ;
			data[41416] <= 8'h10 ;
			data[41417] <= 8'h10 ;
			data[41418] <= 8'h10 ;
			data[41419] <= 8'h10 ;
			data[41420] <= 8'h10 ;
			data[41421] <= 8'h10 ;
			data[41422] <= 8'h10 ;
			data[41423] <= 8'h10 ;
			data[41424] <= 8'h10 ;
			data[41425] <= 8'h10 ;
			data[41426] <= 8'h10 ;
			data[41427] <= 8'h10 ;
			data[41428] <= 8'h10 ;
			data[41429] <= 8'h10 ;
			data[41430] <= 8'h10 ;
			data[41431] <= 8'h10 ;
			data[41432] <= 8'h10 ;
			data[41433] <= 8'h10 ;
			data[41434] <= 8'h10 ;
			data[41435] <= 8'h10 ;
			data[41436] <= 8'h10 ;
			data[41437] <= 8'h10 ;
			data[41438] <= 8'h10 ;
			data[41439] <= 8'h10 ;
			data[41440] <= 8'h10 ;
			data[41441] <= 8'h10 ;
			data[41442] <= 8'h10 ;
			data[41443] <= 8'h10 ;
			data[41444] <= 8'h10 ;
			data[41445] <= 8'h10 ;
			data[41446] <= 8'h10 ;
			data[41447] <= 8'h10 ;
			data[41448] <= 8'h10 ;
			data[41449] <= 8'h10 ;
			data[41450] <= 8'h10 ;
			data[41451] <= 8'h10 ;
			data[41452] <= 8'h10 ;
			data[41453] <= 8'h10 ;
			data[41454] <= 8'h10 ;
			data[41455] <= 8'h10 ;
			data[41456] <= 8'h10 ;
			data[41457] <= 8'h10 ;
			data[41458] <= 8'h10 ;
			data[41459] <= 8'h10 ;
			data[41460] <= 8'h10 ;
			data[41461] <= 8'h10 ;
			data[41462] <= 8'h10 ;
			data[41463] <= 8'h10 ;
			data[41464] <= 8'h10 ;
			data[41465] <= 8'h10 ;
			data[41466] <= 8'h10 ;
			data[41467] <= 8'h10 ;
			data[41468] <= 8'h10 ;
			data[41469] <= 8'h10 ;
			data[41470] <= 8'h10 ;
			data[41471] <= 8'h10 ;
			data[41472] <= 8'h10 ;
			data[41473] <= 8'h10 ;
			data[41474] <= 8'h10 ;
			data[41475] <= 8'h10 ;
			data[41476] <= 8'h10 ;
			data[41477] <= 8'h10 ;
			data[41478] <= 8'h10 ;
			data[41479] <= 8'h10 ;
			data[41480] <= 8'h10 ;
			data[41481] <= 8'h10 ;
			data[41482] <= 8'h10 ;
			data[41483] <= 8'h10 ;
			data[41484] <= 8'h10 ;
			data[41485] <= 8'h10 ;
			data[41486] <= 8'h10 ;
			data[41487] <= 8'h10 ;
			data[41488] <= 8'h10 ;
			data[41489] <= 8'h10 ;
			data[41490] <= 8'h10 ;
			data[41491] <= 8'h10 ;
			data[41492] <= 8'h10 ;
			data[41493] <= 8'h10 ;
			data[41494] <= 8'h10 ;
			data[41495] <= 8'h10 ;
			data[41496] <= 8'h10 ;
			data[41497] <= 8'h10 ;
			data[41498] <= 8'h10 ;
			data[41499] <= 8'h10 ;
			data[41500] <= 8'h10 ;
			data[41501] <= 8'h10 ;
			data[41502] <= 8'h10 ;
			data[41503] <= 8'h10 ;
			data[41504] <= 8'h10 ;
			data[41505] <= 8'h10 ;
			data[41506] <= 8'h10 ;
			data[41507] <= 8'h10 ;
			data[41508] <= 8'h10 ;
			data[41509] <= 8'h10 ;
			data[41510] <= 8'h10 ;
			data[41511] <= 8'h10 ;
			data[41512] <= 8'h10 ;
			data[41513] <= 8'h10 ;
			data[41514] <= 8'h10 ;
			data[41515] <= 8'h10 ;
			data[41516] <= 8'h10 ;
			data[41517] <= 8'h10 ;
			data[41518] <= 8'h10 ;
			data[41519] <= 8'h10 ;
			data[41520] <= 8'h10 ;
			data[41521] <= 8'h10 ;
			data[41522] <= 8'h10 ;
			data[41523] <= 8'h10 ;
			data[41524] <= 8'h10 ;
			data[41525] <= 8'h10 ;
			data[41526] <= 8'h10 ;
			data[41527] <= 8'h10 ;
			data[41528] <= 8'h10 ;
			data[41529] <= 8'h10 ;
			data[41530] <= 8'h10 ;
			data[41531] <= 8'h10 ;
			data[41532] <= 8'h10 ;
			data[41533] <= 8'h10 ;
			data[41534] <= 8'h10 ;
			data[41535] <= 8'h10 ;
			data[41536] <= 8'h10 ;
			data[41537] <= 8'h10 ;
			data[41538] <= 8'h10 ;
			data[41539] <= 8'h10 ;
			data[41540] <= 8'h10 ;
			data[41541] <= 8'h10 ;
			data[41542] <= 8'h10 ;
			data[41543] <= 8'h10 ;
			data[41544] <= 8'h10 ;
			data[41545] <= 8'h10 ;
			data[41546] <= 8'h10 ;
			data[41547] <= 8'h10 ;
			data[41548] <= 8'h10 ;
			data[41549] <= 8'h10 ;
			data[41550] <= 8'h10 ;
			data[41551] <= 8'h10 ;
			data[41552] <= 8'h10 ;
			data[41553] <= 8'h10 ;
			data[41554] <= 8'h10 ;
			data[41555] <= 8'h10 ;
			data[41556] <= 8'h10 ;
			data[41557] <= 8'h10 ;
			data[41558] <= 8'h10 ;
			data[41559] <= 8'h10 ;
			data[41560] <= 8'h10 ;
			data[41561] <= 8'h10 ;
			data[41562] <= 8'h10 ;
			data[41563] <= 8'h10 ;
			data[41564] <= 8'h10 ;
			data[41565] <= 8'h10 ;
			data[41566] <= 8'h10 ;
			data[41567] <= 8'h10 ;
			data[41568] <= 8'h10 ;
			data[41569] <= 8'h10 ;
			data[41570] <= 8'h10 ;
			data[41571] <= 8'h10 ;
			data[41572] <= 8'h10 ;
			data[41573] <= 8'h10 ;
			data[41574] <= 8'h10 ;
			data[41575] <= 8'h10 ;
			data[41576] <= 8'h10 ;
			data[41577] <= 8'h10 ;
			data[41578] <= 8'h10 ;
			data[41579] <= 8'h10 ;
			data[41580] <= 8'h10 ;
			data[41581] <= 8'h10 ;
			data[41582] <= 8'h10 ;
			data[41583] <= 8'h10 ;
			data[41584] <= 8'h10 ;
			data[41585] <= 8'h10 ;
			data[41586] <= 8'h10 ;
			data[41587] <= 8'h10 ;
			data[41588] <= 8'h10 ;
			data[41589] <= 8'h10 ;
			data[41590] <= 8'h10 ;
			data[41591] <= 8'h10 ;
			data[41592] <= 8'h10 ;
			data[41593] <= 8'h10 ;
			data[41594] <= 8'h10 ;
			data[41595] <= 8'h10 ;
			data[41596] <= 8'h10 ;
			data[41597] <= 8'h10 ;
			data[41598] <= 8'h10 ;
			data[41599] <= 8'h10 ;
			data[41600] <= 8'h10 ;
			data[41601] <= 8'h10 ;
			data[41602] <= 8'h10 ;
			data[41603] <= 8'h10 ;
			data[41604] <= 8'h10 ;
			data[41605] <= 8'h10 ;
			data[41606] <= 8'h10 ;
			data[41607] <= 8'h10 ;
			data[41608] <= 8'h10 ;
			data[41609] <= 8'h10 ;
			data[41610] <= 8'h10 ;
			data[41611] <= 8'h10 ;
			data[41612] <= 8'h10 ;
			data[41613] <= 8'h10 ;
			data[41614] <= 8'h10 ;
			data[41615] <= 8'h10 ;
			data[41616] <= 8'h10 ;
			data[41617] <= 8'h10 ;
			data[41618] <= 8'h10 ;
			data[41619] <= 8'h10 ;
			data[41620] <= 8'h10 ;
			data[41621] <= 8'h10 ;
			data[41622] <= 8'h10 ;
			data[41623] <= 8'h10 ;
			data[41624] <= 8'h10 ;
			data[41625] <= 8'h10 ;
			data[41626] <= 8'h10 ;
			data[41627] <= 8'h10 ;
			data[41628] <= 8'h10 ;
			data[41629] <= 8'h10 ;
			data[41630] <= 8'h10 ;
			data[41631] <= 8'h10 ;
			data[41632] <= 8'h10 ;
			data[41633] <= 8'h10 ;
			data[41634] <= 8'h10 ;
			data[41635] <= 8'h10 ;
			data[41636] <= 8'h10 ;
			data[41637] <= 8'h10 ;
			data[41638] <= 8'h10 ;
			data[41639] <= 8'h10 ;
			data[41640] <= 8'h10 ;
			data[41641] <= 8'h10 ;
			data[41642] <= 8'h10 ;
			data[41643] <= 8'h10 ;
			data[41644] <= 8'h10 ;
			data[41645] <= 8'h10 ;
			data[41646] <= 8'h10 ;
			data[41647] <= 8'h10 ;
			data[41648] <= 8'h10 ;
			data[41649] <= 8'h10 ;
			data[41650] <= 8'h10 ;
			data[41651] <= 8'h10 ;
			data[41652] <= 8'h10 ;
			data[41653] <= 8'h10 ;
			data[41654] <= 8'h10 ;
			data[41655] <= 8'h10 ;
			data[41656] <= 8'h10 ;
			data[41657] <= 8'h10 ;
			data[41658] <= 8'h10 ;
			data[41659] <= 8'h10 ;
			data[41660] <= 8'h10 ;
			data[41661] <= 8'h10 ;
			data[41662] <= 8'h10 ;
			data[41663] <= 8'h10 ;
			data[41664] <= 8'h10 ;
			data[41665] <= 8'h10 ;
			data[41666] <= 8'h10 ;
			data[41667] <= 8'h10 ;
			data[41668] <= 8'h10 ;
			data[41669] <= 8'h10 ;
			data[41670] <= 8'h10 ;
			data[41671] <= 8'h10 ;
			data[41672] <= 8'h10 ;
			data[41673] <= 8'h10 ;
			data[41674] <= 8'h10 ;
			data[41675] <= 8'h10 ;
			data[41676] <= 8'h10 ;
			data[41677] <= 8'h10 ;
			data[41678] <= 8'h10 ;
			data[41679] <= 8'h10 ;
			data[41680] <= 8'h10 ;
			data[41681] <= 8'h10 ;
			data[41682] <= 8'h10 ;
			data[41683] <= 8'h10 ;
			data[41684] <= 8'h10 ;
			data[41685] <= 8'h10 ;
			data[41686] <= 8'h10 ;
			data[41687] <= 8'h10 ;
			data[41688] <= 8'h10 ;
			data[41689] <= 8'h10 ;
			data[41690] <= 8'h10 ;
			data[41691] <= 8'h10 ;
			data[41692] <= 8'h10 ;
			data[41693] <= 8'h10 ;
			data[41694] <= 8'h10 ;
			data[41695] <= 8'h10 ;
			data[41696] <= 8'h10 ;
			data[41697] <= 8'h10 ;
			data[41698] <= 8'h10 ;
			data[41699] <= 8'h10 ;
			data[41700] <= 8'h10 ;
			data[41701] <= 8'h10 ;
			data[41702] <= 8'h10 ;
			data[41703] <= 8'h10 ;
			data[41704] <= 8'h10 ;
			data[41705] <= 8'h10 ;
			data[41706] <= 8'h10 ;
			data[41707] <= 8'h10 ;
			data[41708] <= 8'h10 ;
			data[41709] <= 8'h10 ;
			data[41710] <= 8'h10 ;
			data[41711] <= 8'h10 ;
			data[41712] <= 8'h10 ;
			data[41713] <= 8'h10 ;
			data[41714] <= 8'h10 ;
			data[41715] <= 8'h10 ;
			data[41716] <= 8'h10 ;
			data[41717] <= 8'h10 ;
			data[41718] <= 8'h10 ;
			data[41719] <= 8'h10 ;
			data[41720] <= 8'h10 ;
			data[41721] <= 8'h10 ;
			data[41722] <= 8'h10 ;
			data[41723] <= 8'h10 ;
			data[41724] <= 8'h10 ;
			data[41725] <= 8'h10 ;
			data[41726] <= 8'h10 ;
			data[41727] <= 8'h10 ;
			data[41728] <= 8'h10 ;
			data[41729] <= 8'h10 ;
			data[41730] <= 8'h10 ;
			data[41731] <= 8'h10 ;
			data[41732] <= 8'h10 ;
			data[41733] <= 8'h10 ;
			data[41734] <= 8'h10 ;
			data[41735] <= 8'h10 ;
			data[41736] <= 8'h10 ;
			data[41737] <= 8'h10 ;
			data[41738] <= 8'h10 ;
			data[41739] <= 8'h10 ;
			data[41740] <= 8'h10 ;
			data[41741] <= 8'h10 ;
			data[41742] <= 8'h10 ;
			data[41743] <= 8'h10 ;
			data[41744] <= 8'h10 ;
			data[41745] <= 8'h10 ;
			data[41746] <= 8'h10 ;
			data[41747] <= 8'h10 ;
			data[41748] <= 8'h10 ;
			data[41749] <= 8'h10 ;
			data[41750] <= 8'h10 ;
			data[41751] <= 8'h10 ;
			data[41752] <= 8'h10 ;
			data[41753] <= 8'h10 ;
			data[41754] <= 8'h10 ;
			data[41755] <= 8'h10 ;
			data[41756] <= 8'h10 ;
			data[41757] <= 8'h10 ;
			data[41758] <= 8'h10 ;
			data[41759] <= 8'h10 ;
			data[41760] <= 8'h10 ;
			data[41761] <= 8'h10 ;
			data[41762] <= 8'h10 ;
			data[41763] <= 8'h10 ;
			data[41764] <= 8'h10 ;
			data[41765] <= 8'h10 ;
			data[41766] <= 8'h10 ;
			data[41767] <= 8'h10 ;
			data[41768] <= 8'h10 ;
			data[41769] <= 8'h10 ;
			data[41770] <= 8'h10 ;
			data[41771] <= 8'h10 ;
			data[41772] <= 8'h10 ;
			data[41773] <= 8'h10 ;
			data[41774] <= 8'h10 ;
			data[41775] <= 8'h10 ;
			data[41776] <= 8'h10 ;
			data[41777] <= 8'h10 ;
			data[41778] <= 8'h10 ;
			data[41779] <= 8'h10 ;
			data[41780] <= 8'h10 ;
			data[41781] <= 8'h10 ;
			data[41782] <= 8'h10 ;
			data[41783] <= 8'h10 ;
			data[41784] <= 8'h10 ;
			data[41785] <= 8'h10 ;
			data[41786] <= 8'h10 ;
			data[41787] <= 8'h10 ;
			data[41788] <= 8'h10 ;
			data[41789] <= 8'h10 ;
			data[41790] <= 8'h10 ;
			data[41791] <= 8'h10 ;
			data[41792] <= 8'h10 ;
			data[41793] <= 8'h10 ;
			data[41794] <= 8'h10 ;
			data[41795] <= 8'h10 ;
			data[41796] <= 8'h10 ;
			data[41797] <= 8'h10 ;
			data[41798] <= 8'h10 ;
			data[41799] <= 8'h10 ;
			data[41800] <= 8'h10 ;
			data[41801] <= 8'h10 ;
			data[41802] <= 8'h10 ;
			data[41803] <= 8'h10 ;
			data[41804] <= 8'h10 ;
			data[41805] <= 8'h10 ;
			data[41806] <= 8'h10 ;
			data[41807] <= 8'h10 ;
			data[41808] <= 8'h10 ;
			data[41809] <= 8'h10 ;
			data[41810] <= 8'h10 ;
			data[41811] <= 8'h10 ;
			data[41812] <= 8'h10 ;
			data[41813] <= 8'h10 ;
			data[41814] <= 8'h10 ;
			data[41815] <= 8'h10 ;
			data[41816] <= 8'h10 ;
			data[41817] <= 8'h10 ;
			data[41818] <= 8'h10 ;
			data[41819] <= 8'h10 ;
			data[41820] <= 8'h10 ;
			data[41821] <= 8'h10 ;
			data[41822] <= 8'h10 ;
			data[41823] <= 8'h10 ;
			data[41824] <= 8'h10 ;
			data[41825] <= 8'h10 ;
			data[41826] <= 8'h10 ;
			data[41827] <= 8'h10 ;
			data[41828] <= 8'h10 ;
			data[41829] <= 8'h10 ;
			data[41830] <= 8'h10 ;
			data[41831] <= 8'h10 ;
			data[41832] <= 8'h10 ;
			data[41833] <= 8'h10 ;
			data[41834] <= 8'h10 ;
			data[41835] <= 8'h10 ;
			data[41836] <= 8'h10 ;
			data[41837] <= 8'h10 ;
			data[41838] <= 8'h10 ;
			data[41839] <= 8'h10 ;
			data[41840] <= 8'h10 ;
			data[41841] <= 8'h10 ;
			data[41842] <= 8'h10 ;
			data[41843] <= 8'h10 ;
			data[41844] <= 8'h10 ;
			data[41845] <= 8'h10 ;
			data[41846] <= 8'h10 ;
			data[41847] <= 8'h10 ;
			data[41848] <= 8'h10 ;
			data[41849] <= 8'h10 ;
			data[41850] <= 8'h10 ;
			data[41851] <= 8'h10 ;
			data[41852] <= 8'h10 ;
			data[41853] <= 8'h10 ;
			data[41854] <= 8'h10 ;
			data[41855] <= 8'h10 ;
			data[41856] <= 8'h10 ;
			data[41857] <= 8'h10 ;
			data[41858] <= 8'h10 ;
			data[41859] <= 8'h10 ;
			data[41860] <= 8'h10 ;
			data[41861] <= 8'h10 ;
			data[41862] <= 8'h10 ;
			data[41863] <= 8'h10 ;
			data[41864] <= 8'h10 ;
			data[41865] <= 8'h10 ;
			data[41866] <= 8'h10 ;
			data[41867] <= 8'h10 ;
			data[41868] <= 8'h10 ;
			data[41869] <= 8'h10 ;
			data[41870] <= 8'h10 ;
			data[41871] <= 8'h10 ;
			data[41872] <= 8'h10 ;
			data[41873] <= 8'h10 ;
			data[41874] <= 8'h10 ;
			data[41875] <= 8'h10 ;
			data[41876] <= 8'h10 ;
			data[41877] <= 8'h10 ;
			data[41878] <= 8'h10 ;
			data[41879] <= 8'h10 ;
			data[41880] <= 8'h10 ;
			data[41881] <= 8'h10 ;
			data[41882] <= 8'h10 ;
			data[41883] <= 8'h10 ;
			data[41884] <= 8'h10 ;
			data[41885] <= 8'h10 ;
			data[41886] <= 8'h10 ;
			data[41887] <= 8'h10 ;
			data[41888] <= 8'h10 ;
			data[41889] <= 8'h10 ;
			data[41890] <= 8'h10 ;
			data[41891] <= 8'h10 ;
			data[41892] <= 8'h10 ;
			data[41893] <= 8'h10 ;
			data[41894] <= 8'h10 ;
			data[41895] <= 8'h10 ;
			data[41896] <= 8'h10 ;
			data[41897] <= 8'h10 ;
			data[41898] <= 8'h10 ;
			data[41899] <= 8'h10 ;
			data[41900] <= 8'h10 ;
			data[41901] <= 8'h10 ;
			data[41902] <= 8'h10 ;
			data[41903] <= 8'h10 ;
			data[41904] <= 8'h10 ;
			data[41905] <= 8'h10 ;
			data[41906] <= 8'h10 ;
			data[41907] <= 8'h10 ;
			data[41908] <= 8'h10 ;
			data[41909] <= 8'h10 ;
			data[41910] <= 8'h10 ;
			data[41911] <= 8'h10 ;
			data[41912] <= 8'h10 ;
			data[41913] <= 8'h10 ;
			data[41914] <= 8'h10 ;
			data[41915] <= 8'h10 ;
			data[41916] <= 8'h10 ;
			data[41917] <= 8'h10 ;
			data[41918] <= 8'h10 ;
			data[41919] <= 8'h10 ;
			data[41920] <= 8'h10 ;
			data[41921] <= 8'h10 ;
			data[41922] <= 8'h10 ;
			data[41923] <= 8'h10 ;
			data[41924] <= 8'h10 ;
			data[41925] <= 8'h10 ;
			data[41926] <= 8'h10 ;
			data[41927] <= 8'h10 ;
			data[41928] <= 8'h10 ;
			data[41929] <= 8'h10 ;
			data[41930] <= 8'h10 ;
			data[41931] <= 8'h10 ;
			data[41932] <= 8'h10 ;
			data[41933] <= 8'h10 ;
			data[41934] <= 8'h10 ;
			data[41935] <= 8'h10 ;
			data[41936] <= 8'h10 ;
			data[41937] <= 8'h10 ;
			data[41938] <= 8'h10 ;
			data[41939] <= 8'h10 ;
			data[41940] <= 8'h10 ;
			data[41941] <= 8'h10 ;
			data[41942] <= 8'h10 ;
			data[41943] <= 8'h10 ;
			data[41944] <= 8'h10 ;
			data[41945] <= 8'h10 ;
			data[41946] <= 8'h10 ;
			data[41947] <= 8'h10 ;
			data[41948] <= 8'h10 ;
			data[41949] <= 8'h10 ;
			data[41950] <= 8'h10 ;
			data[41951] <= 8'h10 ;
			data[41952] <= 8'h10 ;
			data[41953] <= 8'h10 ;
			data[41954] <= 8'h10 ;
			data[41955] <= 8'h10 ;
			data[41956] <= 8'h10 ;
			data[41957] <= 8'h10 ;
			data[41958] <= 8'h10 ;
			data[41959] <= 8'h10 ;
			data[41960] <= 8'h10 ;
			data[41961] <= 8'h10 ;
			data[41962] <= 8'h10 ;
			data[41963] <= 8'h10 ;
			data[41964] <= 8'h10 ;
			data[41965] <= 8'h10 ;
			data[41966] <= 8'h10 ;
			data[41967] <= 8'h10 ;
			data[41968] <= 8'h10 ;
			data[41969] <= 8'h10 ;
			data[41970] <= 8'h10 ;
			data[41971] <= 8'h10 ;
			data[41972] <= 8'h10 ;
			data[41973] <= 8'h10 ;
			data[41974] <= 8'h10 ;
			data[41975] <= 8'h10 ;
			data[41976] <= 8'h10 ;
			data[41977] <= 8'h10 ;
			data[41978] <= 8'h10 ;
			data[41979] <= 8'h10 ;
			data[41980] <= 8'h10 ;
			data[41981] <= 8'h10 ;
			data[41982] <= 8'h10 ;
			data[41983] <= 8'h10 ;
			data[41984] <= 8'h10 ;
			data[41985] <= 8'h10 ;
			data[41986] <= 8'h10 ;
			data[41987] <= 8'h10 ;
			data[41988] <= 8'h10 ;
			data[41989] <= 8'h10 ;
			data[41990] <= 8'h10 ;
			data[41991] <= 8'h10 ;
			data[41992] <= 8'h10 ;
			data[41993] <= 8'h10 ;
			data[41994] <= 8'h10 ;
			data[41995] <= 8'h10 ;
			data[41996] <= 8'h10 ;
			data[41997] <= 8'h10 ;
			data[41998] <= 8'h10 ;
			data[41999] <= 8'h10 ;
			data[42000] <= 8'h10 ;
			data[42001] <= 8'h10 ;
			data[42002] <= 8'h10 ;
			data[42003] <= 8'h10 ;
			data[42004] <= 8'h10 ;
			data[42005] <= 8'h10 ;
			data[42006] <= 8'h10 ;
			data[42007] <= 8'h10 ;
			data[42008] <= 8'h10 ;
			data[42009] <= 8'h10 ;
			data[42010] <= 8'h10 ;
			data[42011] <= 8'h10 ;
			data[42012] <= 8'h10 ;
			data[42013] <= 8'h10 ;
			data[42014] <= 8'h10 ;
			data[42015] <= 8'h10 ;
			data[42016] <= 8'h10 ;
			data[42017] <= 8'h10 ;
			data[42018] <= 8'h10 ;
			data[42019] <= 8'h10 ;
			data[42020] <= 8'h10 ;
			data[42021] <= 8'h10 ;
			data[42022] <= 8'h10 ;
			data[42023] <= 8'h10 ;
			data[42024] <= 8'h10 ;
			data[42025] <= 8'h10 ;
			data[42026] <= 8'h10 ;
			data[42027] <= 8'h10 ;
			data[42028] <= 8'h10 ;
			data[42029] <= 8'h10 ;
			data[42030] <= 8'h10 ;
			data[42031] <= 8'h10 ;
			data[42032] <= 8'h10 ;
			data[42033] <= 8'h10 ;
			data[42034] <= 8'h10 ;
			data[42035] <= 8'h10 ;
			data[42036] <= 8'h10 ;
			data[42037] <= 8'h10 ;
			data[42038] <= 8'h10 ;
			data[42039] <= 8'h10 ;
			data[42040] <= 8'h10 ;
			data[42041] <= 8'h10 ;
			data[42042] <= 8'h10 ;
			data[42043] <= 8'h10 ;
			data[42044] <= 8'h10 ;
			data[42045] <= 8'h10 ;
			data[42046] <= 8'h10 ;
			data[42047] <= 8'h10 ;
			data[42048] <= 8'h10 ;
			data[42049] <= 8'h10 ;
			data[42050] <= 8'h10 ;
			data[42051] <= 8'h10 ;
			data[42052] <= 8'h10 ;
			data[42053] <= 8'h10 ;
			data[42054] <= 8'h10 ;
			data[42055] <= 8'h10 ;
			data[42056] <= 8'h10 ;
			data[42057] <= 8'h10 ;
			data[42058] <= 8'h10 ;
			data[42059] <= 8'h10 ;
			data[42060] <= 8'h10 ;
			data[42061] <= 8'h10 ;
			data[42062] <= 8'h10 ;
			data[42063] <= 8'h10 ;
			data[42064] <= 8'h10 ;
			data[42065] <= 8'h10 ;
			data[42066] <= 8'h10 ;
			data[42067] <= 8'h10 ;
			data[42068] <= 8'h10 ;
			data[42069] <= 8'h10 ;
			data[42070] <= 8'h10 ;
			data[42071] <= 8'h10 ;
			data[42072] <= 8'h10 ;
			data[42073] <= 8'h10 ;
			data[42074] <= 8'h10 ;
			data[42075] <= 8'h10 ;
			data[42076] <= 8'h10 ;
			data[42077] <= 8'h10 ;
			data[42078] <= 8'h10 ;
			data[42079] <= 8'h10 ;
			data[42080] <= 8'h10 ;
			data[42081] <= 8'h10 ;
			data[42082] <= 8'h10 ;
			data[42083] <= 8'h10 ;
			data[42084] <= 8'h10 ;
			data[42085] <= 8'h10 ;
			data[42086] <= 8'h10 ;
			data[42087] <= 8'h10 ;
			data[42088] <= 8'h10 ;
			data[42089] <= 8'h10 ;
			data[42090] <= 8'h10 ;
			data[42091] <= 8'h10 ;
			data[42092] <= 8'h10 ;
			data[42093] <= 8'h10 ;
			data[42094] <= 8'h10 ;
			data[42095] <= 8'h10 ;
			data[42096] <= 8'h10 ;
			data[42097] <= 8'h10 ;
			data[42098] <= 8'h10 ;
			data[42099] <= 8'h10 ;
			data[42100] <= 8'h10 ;
			data[42101] <= 8'h10 ;
			data[42102] <= 8'h10 ;
			data[42103] <= 8'h10 ;
			data[42104] <= 8'h10 ;
			data[42105] <= 8'h10 ;
			data[42106] <= 8'h10 ;
			data[42107] <= 8'h10 ;
			data[42108] <= 8'h10 ;
			data[42109] <= 8'h10 ;
			data[42110] <= 8'h10 ;
			data[42111] <= 8'h10 ;
			data[42112] <= 8'h10 ;
			data[42113] <= 8'h10 ;
			data[42114] <= 8'h10 ;
			data[42115] <= 8'h10 ;
			data[42116] <= 8'h10 ;
			data[42117] <= 8'h10 ;
			data[42118] <= 8'h10 ;
			data[42119] <= 8'h10 ;
			data[42120] <= 8'h10 ;
			data[42121] <= 8'h10 ;
			data[42122] <= 8'h10 ;
			data[42123] <= 8'h10 ;
			data[42124] <= 8'h10 ;
			data[42125] <= 8'h10 ;
			data[42126] <= 8'h10 ;
			data[42127] <= 8'h10 ;
			data[42128] <= 8'h10 ;
			data[42129] <= 8'h10 ;
			data[42130] <= 8'h10 ;
			data[42131] <= 8'h10 ;
			data[42132] <= 8'h10 ;
			data[42133] <= 8'h10 ;
			data[42134] <= 8'h10 ;
			data[42135] <= 8'h10 ;
			data[42136] <= 8'h10 ;
			data[42137] <= 8'h10 ;
			data[42138] <= 8'h10 ;
			data[42139] <= 8'h10 ;
			data[42140] <= 8'h10 ;
			data[42141] <= 8'h10 ;
			data[42142] <= 8'h10 ;
			data[42143] <= 8'h10 ;
			data[42144] <= 8'h10 ;
			data[42145] <= 8'h10 ;
			data[42146] <= 8'h10 ;
			data[42147] <= 8'h10 ;
			data[42148] <= 8'h10 ;
			data[42149] <= 8'h10 ;
			data[42150] <= 8'h10 ;
			data[42151] <= 8'h10 ;
			data[42152] <= 8'h10 ;
			data[42153] <= 8'h10 ;
			data[42154] <= 8'h10 ;
			data[42155] <= 8'h10 ;
			data[42156] <= 8'h10 ;
			data[42157] <= 8'h10 ;
			data[42158] <= 8'h10 ;
			data[42159] <= 8'h10 ;
			data[42160] <= 8'h10 ;
			data[42161] <= 8'h10 ;
			data[42162] <= 8'h10 ;
			data[42163] <= 8'h10 ;
			data[42164] <= 8'h10 ;
			data[42165] <= 8'h10 ;
			data[42166] <= 8'h10 ;
			data[42167] <= 8'h10 ;
			data[42168] <= 8'h10 ;
			data[42169] <= 8'h10 ;
			data[42170] <= 8'h10 ;
			data[42171] <= 8'h10 ;
			data[42172] <= 8'h10 ;
			data[42173] <= 8'h10 ;
			data[42174] <= 8'h10 ;
			data[42175] <= 8'h10 ;
			data[42176] <= 8'h10 ;
			data[42177] <= 8'h10 ;
			data[42178] <= 8'h10 ;
			data[42179] <= 8'h10 ;
			data[42180] <= 8'h10 ;
			data[42181] <= 8'h10 ;
			data[42182] <= 8'h10 ;
			data[42183] <= 8'h10 ;
			data[42184] <= 8'h10 ;
			data[42185] <= 8'h10 ;
			data[42186] <= 8'h10 ;
			data[42187] <= 8'h10 ;
			data[42188] <= 8'h10 ;
			data[42189] <= 8'h10 ;
			data[42190] <= 8'h10 ;
			data[42191] <= 8'h10 ;
			data[42192] <= 8'h10 ;
			data[42193] <= 8'h10 ;
			data[42194] <= 8'h10 ;
			data[42195] <= 8'h10 ;
			data[42196] <= 8'h10 ;
			data[42197] <= 8'h10 ;
			data[42198] <= 8'h10 ;
			data[42199] <= 8'h10 ;
			data[42200] <= 8'h10 ;
			data[42201] <= 8'h10 ;
			data[42202] <= 8'h10 ;
			data[42203] <= 8'h10 ;
			data[42204] <= 8'h10 ;
			data[42205] <= 8'h10 ;
			data[42206] <= 8'h10 ;
			data[42207] <= 8'h10 ;
			data[42208] <= 8'h10 ;
			data[42209] <= 8'h10 ;
			data[42210] <= 8'h10 ;
			data[42211] <= 8'h10 ;
			data[42212] <= 8'h10 ;
			data[42213] <= 8'h10 ;
			data[42214] <= 8'h10 ;
			data[42215] <= 8'h10 ;
			data[42216] <= 8'h10 ;
			data[42217] <= 8'h10 ;
			data[42218] <= 8'h10 ;
			data[42219] <= 8'h10 ;
			data[42220] <= 8'h10 ;
			data[42221] <= 8'h10 ;
			data[42222] <= 8'h10 ;
			data[42223] <= 8'h10 ;
			data[42224] <= 8'h10 ;
			data[42225] <= 8'h10 ;
			data[42226] <= 8'h10 ;
			data[42227] <= 8'h10 ;
			data[42228] <= 8'h10 ;
			data[42229] <= 8'h10 ;
			data[42230] <= 8'h10 ;
			data[42231] <= 8'h10 ;
			data[42232] <= 8'h10 ;
			data[42233] <= 8'h10 ;
			data[42234] <= 8'h10 ;
			data[42235] <= 8'h10 ;
			data[42236] <= 8'h10 ;
			data[42237] <= 8'h10 ;
			data[42238] <= 8'h10 ;
			data[42239] <= 8'h10 ;
			data[42240] <= 8'h10 ;
			data[42241] <= 8'h10 ;
			data[42242] <= 8'h10 ;
			data[42243] <= 8'h10 ;
			data[42244] <= 8'h10 ;
			data[42245] <= 8'h10 ;
			data[42246] <= 8'h10 ;
			data[42247] <= 8'h10 ;
			data[42248] <= 8'h10 ;
			data[42249] <= 8'h10 ;
			data[42250] <= 8'h10 ;
			data[42251] <= 8'h10 ;
			data[42252] <= 8'h10 ;
			data[42253] <= 8'h10 ;
			data[42254] <= 8'h10 ;
			data[42255] <= 8'h10 ;
			data[42256] <= 8'h10 ;
			data[42257] <= 8'h10 ;
			data[42258] <= 8'h10 ;
			data[42259] <= 8'h10 ;
			data[42260] <= 8'h10 ;
			data[42261] <= 8'h10 ;
			data[42262] <= 8'h10 ;
			data[42263] <= 8'h10 ;
			data[42264] <= 8'h10 ;
			data[42265] <= 8'h10 ;
			data[42266] <= 8'h10 ;
			data[42267] <= 8'h10 ;
			data[42268] <= 8'h10 ;
			data[42269] <= 8'h10 ;
			data[42270] <= 8'h10 ;
			data[42271] <= 8'h10 ;
			data[42272] <= 8'h10 ;
			data[42273] <= 8'h10 ;
			data[42274] <= 8'h10 ;
			data[42275] <= 8'h10 ;
			data[42276] <= 8'h10 ;
			data[42277] <= 8'h10 ;
			data[42278] <= 8'h10 ;
			data[42279] <= 8'h10 ;
			data[42280] <= 8'h10 ;
			data[42281] <= 8'h10 ;
			data[42282] <= 8'h10 ;
			data[42283] <= 8'h10 ;
			data[42284] <= 8'h10 ;
			data[42285] <= 8'h10 ;
			data[42286] <= 8'h10 ;
			data[42287] <= 8'h10 ;
			data[42288] <= 8'h10 ;
			data[42289] <= 8'h10 ;
			data[42290] <= 8'h10 ;
			data[42291] <= 8'h10 ;
			data[42292] <= 8'h10 ;
			data[42293] <= 8'h10 ;
			data[42294] <= 8'h10 ;
			data[42295] <= 8'h10 ;
			data[42296] <= 8'h10 ;
			data[42297] <= 8'h10 ;
			data[42298] <= 8'h10 ;
			data[42299] <= 8'h10 ;
			data[42300] <= 8'h10 ;
			data[42301] <= 8'h10 ;
			data[42302] <= 8'h10 ;
			data[42303] <= 8'h10 ;
			data[42304] <= 8'h10 ;
			data[42305] <= 8'h10 ;
			data[42306] <= 8'h10 ;
			data[42307] <= 8'h10 ;
			data[42308] <= 8'h10 ;
			data[42309] <= 8'h10 ;
			data[42310] <= 8'h10 ;
			data[42311] <= 8'h10 ;
			data[42312] <= 8'h10 ;
			data[42313] <= 8'h10 ;
			data[42314] <= 8'h10 ;
			data[42315] <= 8'h10 ;
			data[42316] <= 8'h10 ;
			data[42317] <= 8'h10 ;
			data[42318] <= 8'h10 ;
			data[42319] <= 8'h10 ;
			data[42320] <= 8'h10 ;
			data[42321] <= 8'h10 ;
			data[42322] <= 8'h10 ;
			data[42323] <= 8'h10 ;
			data[42324] <= 8'h10 ;
			data[42325] <= 8'h10 ;
			data[42326] <= 8'h10 ;
			data[42327] <= 8'h10 ;
			data[42328] <= 8'h10 ;
			data[42329] <= 8'h10 ;
			data[42330] <= 8'h10 ;
			data[42331] <= 8'h10 ;
			data[42332] <= 8'h10 ;
			data[42333] <= 8'h10 ;
			data[42334] <= 8'h10 ;
			data[42335] <= 8'h10 ;
			data[42336] <= 8'h10 ;
			data[42337] <= 8'h10 ;
			data[42338] <= 8'h10 ;
			data[42339] <= 8'h10 ;
			data[42340] <= 8'h10 ;
			data[42341] <= 8'h10 ;
			data[42342] <= 8'h10 ;
			data[42343] <= 8'h10 ;
			data[42344] <= 8'h10 ;
			data[42345] <= 8'h10 ;
			data[42346] <= 8'h10 ;
			data[42347] <= 8'h10 ;
			data[42348] <= 8'h10 ;
			data[42349] <= 8'h10 ;
			data[42350] <= 8'h10 ;
			data[42351] <= 8'h10 ;
			data[42352] <= 8'h10 ;
			data[42353] <= 8'h10 ;
			data[42354] <= 8'h10 ;
			data[42355] <= 8'h10 ;
			data[42356] <= 8'h10 ;
			data[42357] <= 8'h10 ;
			data[42358] <= 8'h10 ;
			data[42359] <= 8'h10 ;
			data[42360] <= 8'h10 ;
			data[42361] <= 8'h10 ;
			data[42362] <= 8'h10 ;
			data[42363] <= 8'h10 ;
			data[42364] <= 8'h10 ;
			data[42365] <= 8'h10 ;
			data[42366] <= 8'h10 ;
			data[42367] <= 8'h10 ;
			data[42368] <= 8'h10 ;
			data[42369] <= 8'h10 ;
			data[42370] <= 8'h10 ;
			data[42371] <= 8'h10 ;
			data[42372] <= 8'h10 ;
			data[42373] <= 8'h10 ;
			data[42374] <= 8'h10 ;
			data[42375] <= 8'h10 ;
			data[42376] <= 8'h10 ;
			data[42377] <= 8'h10 ;
			data[42378] <= 8'h10 ;
			data[42379] <= 8'h10 ;
			data[42380] <= 8'h10 ;
			data[42381] <= 8'h10 ;
			data[42382] <= 8'h10 ;
			data[42383] <= 8'h10 ;
			data[42384] <= 8'h10 ;
			data[42385] <= 8'h10 ;
			data[42386] <= 8'h10 ;
			data[42387] <= 8'h10 ;
			data[42388] <= 8'h10 ;
			data[42389] <= 8'h10 ;
			data[42390] <= 8'h10 ;
			data[42391] <= 8'h10 ;
			data[42392] <= 8'h10 ;
			data[42393] <= 8'h10 ;
			data[42394] <= 8'h10 ;
			data[42395] <= 8'h10 ;
			data[42396] <= 8'h10 ;
			data[42397] <= 8'h10 ;
			data[42398] <= 8'h10 ;
			data[42399] <= 8'h10 ;
			data[42400] <= 8'h10 ;
			data[42401] <= 8'h10 ;
			data[42402] <= 8'h10 ;
			data[42403] <= 8'h10 ;
			data[42404] <= 8'h10 ;
			data[42405] <= 8'h10 ;
			data[42406] <= 8'h10 ;
			data[42407] <= 8'h10 ;
			data[42408] <= 8'h10 ;
			data[42409] <= 8'h10 ;
			data[42410] <= 8'h10 ;
			data[42411] <= 8'h10 ;
			data[42412] <= 8'h10 ;
			data[42413] <= 8'h10 ;
			data[42414] <= 8'h10 ;
			data[42415] <= 8'h10 ;
			data[42416] <= 8'h10 ;
			data[42417] <= 8'h10 ;
			data[42418] <= 8'h10 ;
			data[42419] <= 8'h10 ;
			data[42420] <= 8'h10 ;
			data[42421] <= 8'h10 ;
			data[42422] <= 8'h10 ;
			data[42423] <= 8'h10 ;
			data[42424] <= 8'h10 ;
			data[42425] <= 8'h10 ;
			data[42426] <= 8'h10 ;
			data[42427] <= 8'h10 ;
			data[42428] <= 8'h10 ;
			data[42429] <= 8'h10 ;
			data[42430] <= 8'h10 ;
			data[42431] <= 8'h10 ;
			data[42432] <= 8'h10 ;
			data[42433] <= 8'h10 ;
			data[42434] <= 8'h10 ;
			data[42435] <= 8'h10 ;
			data[42436] <= 8'h10 ;
			data[42437] <= 8'h10 ;
			data[42438] <= 8'h10 ;
			data[42439] <= 8'h10 ;
			data[42440] <= 8'h10 ;
			data[42441] <= 8'h10 ;
			data[42442] <= 8'h10 ;
			data[42443] <= 8'h10 ;
			data[42444] <= 8'h10 ;
			data[42445] <= 8'h10 ;
			data[42446] <= 8'h10 ;
			data[42447] <= 8'h10 ;
			data[42448] <= 8'h10 ;
			data[42449] <= 8'h10 ;
			data[42450] <= 8'h10 ;
			data[42451] <= 8'h10 ;
			data[42452] <= 8'h10 ;
			data[42453] <= 8'h10 ;
			data[42454] <= 8'h10 ;
			data[42455] <= 8'h10 ;
			data[42456] <= 8'h10 ;
			data[42457] <= 8'h10 ;
			data[42458] <= 8'h10 ;
			data[42459] <= 8'h10 ;
			data[42460] <= 8'h10 ;
			data[42461] <= 8'h10 ;
			data[42462] <= 8'h10 ;
			data[42463] <= 8'h10 ;
			data[42464] <= 8'h10 ;
			data[42465] <= 8'h10 ;
			data[42466] <= 8'h10 ;
			data[42467] <= 8'h10 ;
			data[42468] <= 8'h10 ;
			data[42469] <= 8'h10 ;
			data[42470] <= 8'h10 ;
			data[42471] <= 8'h10 ;
			data[42472] <= 8'h10 ;
			data[42473] <= 8'h10 ;
			data[42474] <= 8'h10 ;
			data[42475] <= 8'h10 ;
			data[42476] <= 8'h10 ;
			data[42477] <= 8'h10 ;
			data[42478] <= 8'h10 ;
			data[42479] <= 8'h10 ;
			data[42480] <= 8'h10 ;
			data[42481] <= 8'h10 ;
			data[42482] <= 8'h10 ;
			data[42483] <= 8'h10 ;
			data[42484] <= 8'h10 ;
			data[42485] <= 8'h10 ;
			data[42486] <= 8'h10 ;
			data[42487] <= 8'h10 ;
			data[42488] <= 8'h10 ;
			data[42489] <= 8'h10 ;
			data[42490] <= 8'h10 ;
			data[42491] <= 8'h10 ;
			data[42492] <= 8'h10 ;
			data[42493] <= 8'h10 ;
			data[42494] <= 8'h10 ;
			data[42495] <= 8'h10 ;
			data[42496] <= 8'h10 ;
			data[42497] <= 8'h10 ;
			data[42498] <= 8'h10 ;
			data[42499] <= 8'h10 ;
			data[42500] <= 8'h10 ;
			data[42501] <= 8'h10 ;
			data[42502] <= 8'h10 ;
			data[42503] <= 8'h10 ;
			data[42504] <= 8'h10 ;
			data[42505] <= 8'h10 ;
			data[42506] <= 8'h10 ;
			data[42507] <= 8'h10 ;
			data[42508] <= 8'h10 ;
			data[42509] <= 8'h10 ;
			data[42510] <= 8'h10 ;
			data[42511] <= 8'h10 ;
			data[42512] <= 8'h10 ;
			data[42513] <= 8'h10 ;
			data[42514] <= 8'h10 ;
			data[42515] <= 8'h10 ;
			data[42516] <= 8'h10 ;
			data[42517] <= 8'h10 ;
			data[42518] <= 8'h10 ;
			data[42519] <= 8'h10 ;
			data[42520] <= 8'h10 ;
			data[42521] <= 8'h10 ;
			data[42522] <= 8'h10 ;
			data[42523] <= 8'h10 ;
			data[42524] <= 8'h10 ;
			data[42525] <= 8'h10 ;
			data[42526] <= 8'h10 ;
			data[42527] <= 8'h10 ;
			data[42528] <= 8'h10 ;
			data[42529] <= 8'h10 ;
			data[42530] <= 8'h10 ;
			data[42531] <= 8'h10 ;
			data[42532] <= 8'h10 ;
			data[42533] <= 8'h10 ;
			data[42534] <= 8'h10 ;
			data[42535] <= 8'h10 ;
			data[42536] <= 8'h10 ;
			data[42537] <= 8'h10 ;
			data[42538] <= 8'h10 ;
			data[42539] <= 8'h10 ;
			data[42540] <= 8'h10 ;
			data[42541] <= 8'h10 ;
			data[42542] <= 8'h10 ;
			data[42543] <= 8'h10 ;
			data[42544] <= 8'h10 ;
			data[42545] <= 8'h10 ;
			data[42546] <= 8'h10 ;
			data[42547] <= 8'h10 ;
			data[42548] <= 8'h10 ;
			data[42549] <= 8'h10 ;
			data[42550] <= 8'h10 ;
			data[42551] <= 8'h10 ;
			data[42552] <= 8'h10 ;
			data[42553] <= 8'h10 ;
			data[42554] <= 8'h10 ;
			data[42555] <= 8'h10 ;
			data[42556] <= 8'h10 ;
			data[42557] <= 8'h10 ;
			data[42558] <= 8'h10 ;
			data[42559] <= 8'h10 ;
			data[42560] <= 8'h10 ;
			data[42561] <= 8'h10 ;
			data[42562] <= 8'h10 ;
			data[42563] <= 8'h10 ;
			data[42564] <= 8'h10 ;
			data[42565] <= 8'h10 ;
			data[42566] <= 8'h10 ;
			data[42567] <= 8'h10 ;
			data[42568] <= 8'h10 ;
			data[42569] <= 8'h10 ;
			data[42570] <= 8'h10 ;
			data[42571] <= 8'h10 ;
			data[42572] <= 8'h10 ;
			data[42573] <= 8'h10 ;
			data[42574] <= 8'h10 ;
			data[42575] <= 8'h10 ;
			data[42576] <= 8'h10 ;
			data[42577] <= 8'h10 ;
			data[42578] <= 8'h10 ;
			data[42579] <= 8'h10 ;
			data[42580] <= 8'h10 ;
			data[42581] <= 8'h10 ;
			data[42582] <= 8'h10 ;
			data[42583] <= 8'h10 ;
			data[42584] <= 8'h10 ;
			data[42585] <= 8'h10 ;
			data[42586] <= 8'h10 ;
			data[42587] <= 8'h10 ;
			data[42588] <= 8'h10 ;
			data[42589] <= 8'h10 ;
			data[42590] <= 8'h10 ;
			data[42591] <= 8'h10 ;
			data[42592] <= 8'h10 ;
			data[42593] <= 8'h10 ;
			data[42594] <= 8'h10 ;
			data[42595] <= 8'h10 ;
			data[42596] <= 8'h10 ;
			data[42597] <= 8'h10 ;
			data[42598] <= 8'h10 ;
			data[42599] <= 8'h10 ;
			data[42600] <= 8'h10 ;
			data[42601] <= 8'h10 ;
			data[42602] <= 8'h10 ;
			data[42603] <= 8'h10 ;
			data[42604] <= 8'h10 ;
			data[42605] <= 8'h10 ;
			data[42606] <= 8'h10 ;
			data[42607] <= 8'h10 ;
			data[42608] <= 8'h10 ;
			data[42609] <= 8'h10 ;
			data[42610] <= 8'h10 ;
			data[42611] <= 8'h10 ;
			data[42612] <= 8'h10 ;
			data[42613] <= 8'h10 ;
			data[42614] <= 8'h10 ;
			data[42615] <= 8'h10 ;
			data[42616] <= 8'h10 ;
			data[42617] <= 8'h10 ;
			data[42618] <= 8'h10 ;
			data[42619] <= 8'h10 ;
			data[42620] <= 8'h10 ;
			data[42621] <= 8'h10 ;
			data[42622] <= 8'h10 ;
			data[42623] <= 8'h10 ;
			data[42624] <= 8'h10 ;
			data[42625] <= 8'h10 ;
			data[42626] <= 8'h10 ;
			data[42627] <= 8'h10 ;
			data[42628] <= 8'h10 ;
			data[42629] <= 8'h10 ;
			data[42630] <= 8'h10 ;
			data[42631] <= 8'h10 ;
			data[42632] <= 8'h10 ;
			data[42633] <= 8'h10 ;
			data[42634] <= 8'h10 ;
			data[42635] <= 8'h10 ;
			data[42636] <= 8'h10 ;
			data[42637] <= 8'h10 ;
			data[42638] <= 8'h10 ;
			data[42639] <= 8'h10 ;
			data[42640] <= 8'h10 ;
			data[42641] <= 8'h10 ;
			data[42642] <= 8'h10 ;
			data[42643] <= 8'h10 ;
			data[42644] <= 8'h10 ;
			data[42645] <= 8'h10 ;
			data[42646] <= 8'h10 ;
			data[42647] <= 8'h10 ;
			data[42648] <= 8'h10 ;
			data[42649] <= 8'h10 ;
			data[42650] <= 8'h10 ;
			data[42651] <= 8'h10 ;
			data[42652] <= 8'h10 ;
			data[42653] <= 8'h10 ;
			data[42654] <= 8'h10 ;
			data[42655] <= 8'h10 ;
			data[42656] <= 8'h10 ;
			data[42657] <= 8'h10 ;
			data[42658] <= 8'h10 ;
			data[42659] <= 8'h10 ;
			data[42660] <= 8'h10 ;
			data[42661] <= 8'h10 ;
			data[42662] <= 8'h10 ;
			data[42663] <= 8'h10 ;
			data[42664] <= 8'h10 ;
			data[42665] <= 8'h10 ;
			data[42666] <= 8'h10 ;
			data[42667] <= 8'h10 ;
			data[42668] <= 8'h10 ;
			data[42669] <= 8'h10 ;
			data[42670] <= 8'h10 ;
			data[42671] <= 8'h10 ;
			data[42672] <= 8'h10 ;
			data[42673] <= 8'h10 ;
			data[42674] <= 8'h10 ;
			data[42675] <= 8'h10 ;
			data[42676] <= 8'h10 ;
			data[42677] <= 8'h10 ;
			data[42678] <= 8'h10 ;
			data[42679] <= 8'h10 ;
			data[42680] <= 8'h10 ;
			data[42681] <= 8'h10 ;
			data[42682] <= 8'h10 ;
			data[42683] <= 8'h10 ;
			data[42684] <= 8'h10 ;
			data[42685] <= 8'h10 ;
			data[42686] <= 8'h10 ;
			data[42687] <= 8'h10 ;
			data[42688] <= 8'h10 ;
			data[42689] <= 8'h10 ;
			data[42690] <= 8'h10 ;
			data[42691] <= 8'h10 ;
			data[42692] <= 8'h10 ;
			data[42693] <= 8'h10 ;
			data[42694] <= 8'h10 ;
			data[42695] <= 8'h10 ;
			data[42696] <= 8'h10 ;
			data[42697] <= 8'h10 ;
			data[42698] <= 8'h10 ;
			data[42699] <= 8'h10 ;
			data[42700] <= 8'h10 ;
			data[42701] <= 8'h10 ;
			data[42702] <= 8'h10 ;
			data[42703] <= 8'h10 ;
			data[42704] <= 8'h10 ;
			data[42705] <= 8'h10 ;
			data[42706] <= 8'h10 ;
			data[42707] <= 8'h10 ;
			data[42708] <= 8'h10 ;
			data[42709] <= 8'h10 ;
			data[42710] <= 8'h10 ;
			data[42711] <= 8'h10 ;
			data[42712] <= 8'h10 ;
			data[42713] <= 8'h10 ;
			data[42714] <= 8'h10 ;
			data[42715] <= 8'h10 ;
			data[42716] <= 8'h10 ;
			data[42717] <= 8'h10 ;
			data[42718] <= 8'h10 ;
			data[42719] <= 8'h10 ;
			data[42720] <= 8'h10 ;
			data[42721] <= 8'h10 ;
			data[42722] <= 8'h10 ;
			data[42723] <= 8'h10 ;
			data[42724] <= 8'h10 ;
			data[42725] <= 8'h10 ;
			data[42726] <= 8'h10 ;
			data[42727] <= 8'h10 ;
			data[42728] <= 8'h10 ;
			data[42729] <= 8'h10 ;
			data[42730] <= 8'h10 ;
			data[42731] <= 8'h10 ;
			data[42732] <= 8'h10 ;
			data[42733] <= 8'h10 ;
			data[42734] <= 8'h10 ;
			data[42735] <= 8'h10 ;
			data[42736] <= 8'h10 ;
			data[42737] <= 8'h10 ;
			data[42738] <= 8'h10 ;
			data[42739] <= 8'h10 ;
			data[42740] <= 8'h10 ;
			data[42741] <= 8'h10 ;
			data[42742] <= 8'h10 ;
			data[42743] <= 8'h10 ;
			data[42744] <= 8'h10 ;
			data[42745] <= 8'h10 ;
			data[42746] <= 8'h10 ;
			data[42747] <= 8'h10 ;
			data[42748] <= 8'h10 ;
			data[42749] <= 8'h10 ;
			data[42750] <= 8'h10 ;
			data[42751] <= 8'h10 ;
			data[42752] <= 8'h10 ;
			data[42753] <= 8'h10 ;
			data[42754] <= 8'h10 ;
			data[42755] <= 8'h10 ;
			data[42756] <= 8'h10 ;
			data[42757] <= 8'h10 ;
			data[42758] <= 8'h10 ;
			data[42759] <= 8'h10 ;
			data[42760] <= 8'h10 ;
			data[42761] <= 8'h10 ;
			data[42762] <= 8'h10 ;
			data[42763] <= 8'h10 ;
			data[42764] <= 8'h10 ;
			data[42765] <= 8'h10 ;
			data[42766] <= 8'h10 ;
			data[42767] <= 8'h10 ;
			data[42768] <= 8'h10 ;
			data[42769] <= 8'h10 ;
			data[42770] <= 8'h10 ;
			data[42771] <= 8'h10 ;
			data[42772] <= 8'h10 ;
			data[42773] <= 8'h10 ;
			data[42774] <= 8'h10 ;
			data[42775] <= 8'h10 ;
			data[42776] <= 8'h10 ;
			data[42777] <= 8'h10 ;
			data[42778] <= 8'h10 ;
			data[42779] <= 8'h10 ;
			data[42780] <= 8'h10 ;
			data[42781] <= 8'h10 ;
			data[42782] <= 8'h10 ;
			data[42783] <= 8'h10 ;
			data[42784] <= 8'h10 ;
			data[42785] <= 8'h10 ;
			data[42786] <= 8'h10 ;
			data[42787] <= 8'h10 ;
			data[42788] <= 8'h10 ;
			data[42789] <= 8'h10 ;
			data[42790] <= 8'h10 ;
			data[42791] <= 8'h10 ;
			data[42792] <= 8'h10 ;
			data[42793] <= 8'h10 ;
			data[42794] <= 8'h10 ;
			data[42795] <= 8'h10 ;
			data[42796] <= 8'h10 ;
			data[42797] <= 8'h10 ;
			data[42798] <= 8'h10 ;
			data[42799] <= 8'h10 ;
			data[42800] <= 8'h10 ;
			data[42801] <= 8'h10 ;
			data[42802] <= 8'h10 ;
			data[42803] <= 8'h10 ;
			data[42804] <= 8'h10 ;
			data[42805] <= 8'h10 ;
			data[42806] <= 8'h10 ;
			data[42807] <= 8'h10 ;
			data[42808] <= 8'h10 ;
			data[42809] <= 8'h10 ;
			data[42810] <= 8'h10 ;
			data[42811] <= 8'h10 ;
			data[42812] <= 8'h10 ;
			data[42813] <= 8'h10 ;
			data[42814] <= 8'h10 ;
			data[42815] <= 8'h10 ;
			data[42816] <= 8'h10 ;
			data[42817] <= 8'h10 ;
			data[42818] <= 8'h10 ;
			data[42819] <= 8'h10 ;
			data[42820] <= 8'h10 ;
			data[42821] <= 8'h10 ;
			data[42822] <= 8'h10 ;
			data[42823] <= 8'h10 ;
			data[42824] <= 8'h10 ;
			data[42825] <= 8'h10 ;
			data[42826] <= 8'h10 ;
			data[42827] <= 8'h10 ;
			data[42828] <= 8'h10 ;
			data[42829] <= 8'h10 ;
			data[42830] <= 8'h10 ;
			data[42831] <= 8'h10 ;
			data[42832] <= 8'h10 ;
			data[42833] <= 8'h10 ;
			data[42834] <= 8'h10 ;
			data[42835] <= 8'h10 ;
			data[42836] <= 8'h10 ;
			data[42837] <= 8'h10 ;
			data[42838] <= 8'h10 ;
			data[42839] <= 8'h10 ;
			data[42840] <= 8'h10 ;
			data[42841] <= 8'h10 ;
			data[42842] <= 8'h10 ;
			data[42843] <= 8'h10 ;
			data[42844] <= 8'h10 ;
			data[42845] <= 8'h10 ;
			data[42846] <= 8'h10 ;
			data[42847] <= 8'h10 ;
			data[42848] <= 8'h10 ;
			data[42849] <= 8'h10 ;
			data[42850] <= 8'h10 ;
			data[42851] <= 8'h10 ;
			data[42852] <= 8'h10 ;
			data[42853] <= 8'h10 ;
			data[42854] <= 8'h10 ;
			data[42855] <= 8'h10 ;
			data[42856] <= 8'h10 ;
			data[42857] <= 8'h10 ;
			data[42858] <= 8'h10 ;
			data[42859] <= 8'h10 ;
			data[42860] <= 8'h10 ;
			data[42861] <= 8'h10 ;
			data[42862] <= 8'h10 ;
			data[42863] <= 8'h10 ;
			data[42864] <= 8'h10 ;
			data[42865] <= 8'h10 ;
			data[42866] <= 8'h10 ;
			data[42867] <= 8'h10 ;
			data[42868] <= 8'h10 ;
			data[42869] <= 8'h10 ;
			data[42870] <= 8'h10 ;
			data[42871] <= 8'h10 ;
			data[42872] <= 8'h10 ;
			data[42873] <= 8'h10 ;
			data[42874] <= 8'h10 ;
			data[42875] <= 8'h10 ;
			data[42876] <= 8'h10 ;
			data[42877] <= 8'h10 ;
			data[42878] <= 8'h10 ;
			data[42879] <= 8'h10 ;
			data[42880] <= 8'h10 ;
			data[42881] <= 8'h10 ;
			data[42882] <= 8'h10 ;
			data[42883] <= 8'h10 ;
			data[42884] <= 8'h10 ;
			data[42885] <= 8'h10 ;
			data[42886] <= 8'h10 ;
			data[42887] <= 8'h10 ;
			data[42888] <= 8'h10 ;
			data[42889] <= 8'h10 ;
			data[42890] <= 8'h10 ;
			data[42891] <= 8'h10 ;
			data[42892] <= 8'h10 ;
			data[42893] <= 8'h10 ;
			data[42894] <= 8'h10 ;
			data[42895] <= 8'h10 ;
			data[42896] <= 8'h10 ;
			data[42897] <= 8'h10 ;
			data[42898] <= 8'h10 ;
			data[42899] <= 8'h10 ;
			data[42900] <= 8'h10 ;
			data[42901] <= 8'h10 ;
			data[42902] <= 8'h10 ;
			data[42903] <= 8'h10 ;
			data[42904] <= 8'h10 ;
			data[42905] <= 8'h10 ;
			data[42906] <= 8'h10 ;
			data[42907] <= 8'h10 ;
			data[42908] <= 8'h10 ;
			data[42909] <= 8'h10 ;
			data[42910] <= 8'h10 ;
			data[42911] <= 8'h10 ;
			data[42912] <= 8'h10 ;
			data[42913] <= 8'h10 ;
			data[42914] <= 8'h10 ;
			data[42915] <= 8'h10 ;
			data[42916] <= 8'h10 ;
			data[42917] <= 8'h10 ;
			data[42918] <= 8'h10 ;
			data[42919] <= 8'h10 ;
			data[42920] <= 8'h10 ;
			data[42921] <= 8'h10 ;
			data[42922] <= 8'h10 ;
			data[42923] <= 8'h10 ;
			data[42924] <= 8'h10 ;
			data[42925] <= 8'h10 ;
			data[42926] <= 8'h10 ;
			data[42927] <= 8'h10 ;
			data[42928] <= 8'h10 ;
			data[42929] <= 8'h10 ;
			data[42930] <= 8'h10 ;
			data[42931] <= 8'h10 ;
			data[42932] <= 8'h10 ;
			data[42933] <= 8'h10 ;
			data[42934] <= 8'h10 ;
			data[42935] <= 8'h10 ;
			data[42936] <= 8'h10 ;
			data[42937] <= 8'h10 ;
			data[42938] <= 8'h10 ;
			data[42939] <= 8'h10 ;
			data[42940] <= 8'h10 ;
			data[42941] <= 8'h10 ;
			data[42942] <= 8'h10 ;
			data[42943] <= 8'h10 ;
			data[42944] <= 8'h10 ;
			data[42945] <= 8'h10 ;
			data[42946] <= 8'h10 ;
			data[42947] <= 8'h10 ;
			data[42948] <= 8'h10 ;
			data[42949] <= 8'h10 ;
			data[42950] <= 8'h10 ;
			data[42951] <= 8'h10 ;
			data[42952] <= 8'h10 ;
			data[42953] <= 8'h10 ;
			data[42954] <= 8'h10 ;
			data[42955] <= 8'h10 ;
			data[42956] <= 8'h10 ;
			data[42957] <= 8'h10 ;
			data[42958] <= 8'h10 ;
			data[42959] <= 8'h10 ;
			data[42960] <= 8'h10 ;
			data[42961] <= 8'h10 ;
			data[42962] <= 8'h10 ;
			data[42963] <= 8'h10 ;
			data[42964] <= 8'h10 ;
			data[42965] <= 8'h10 ;
			data[42966] <= 8'h10 ;
			data[42967] <= 8'h10 ;
			data[42968] <= 8'h10 ;
			data[42969] <= 8'h10 ;
			data[42970] <= 8'h10 ;
			data[42971] <= 8'h10 ;
			data[42972] <= 8'h10 ;
			data[42973] <= 8'h10 ;
			data[42974] <= 8'h10 ;
			data[42975] <= 8'h10 ;
			data[42976] <= 8'h10 ;
			data[42977] <= 8'h10 ;
			data[42978] <= 8'h10 ;
			data[42979] <= 8'h10 ;
			data[42980] <= 8'h10 ;
			data[42981] <= 8'h10 ;
			data[42982] <= 8'h10 ;
			data[42983] <= 8'h10 ;
			data[42984] <= 8'h10 ;
			data[42985] <= 8'h10 ;
			data[42986] <= 8'h10 ;
			data[42987] <= 8'h10 ;
			data[42988] <= 8'h10 ;
			data[42989] <= 8'h10 ;
			data[42990] <= 8'h10 ;
			data[42991] <= 8'h10 ;
			data[42992] <= 8'h10 ;
			data[42993] <= 8'h10 ;
			data[42994] <= 8'h10 ;
			data[42995] <= 8'h10 ;
			data[42996] <= 8'h10 ;
			data[42997] <= 8'h10 ;
			data[42998] <= 8'h10 ;
			data[42999] <= 8'h10 ;
			data[43000] <= 8'h10 ;
			data[43001] <= 8'h10 ;
			data[43002] <= 8'h10 ;
			data[43003] <= 8'h10 ;
			data[43004] <= 8'h10 ;
			data[43005] <= 8'h10 ;
			data[43006] <= 8'h10 ;
			data[43007] <= 8'h10 ;
			data[43008] <= 8'h10 ;
			data[43009] <= 8'h10 ;
			data[43010] <= 8'h10 ;
			data[43011] <= 8'h10 ;
			data[43012] <= 8'h10 ;
			data[43013] <= 8'h10 ;
			data[43014] <= 8'h10 ;
			data[43015] <= 8'h10 ;
			data[43016] <= 8'h10 ;
			data[43017] <= 8'h10 ;
			data[43018] <= 8'h10 ;
			data[43019] <= 8'h10 ;
			data[43020] <= 8'h10 ;
			data[43021] <= 8'h10 ;
			data[43022] <= 8'h10 ;
			data[43023] <= 8'h10 ;
			data[43024] <= 8'h10 ;
			data[43025] <= 8'h10 ;
			data[43026] <= 8'h10 ;
			data[43027] <= 8'h10 ;
			data[43028] <= 8'h10 ;
			data[43029] <= 8'h10 ;
			data[43030] <= 8'h10 ;
			data[43031] <= 8'h10 ;
			data[43032] <= 8'h10 ;
			data[43033] <= 8'h10 ;
			data[43034] <= 8'h10 ;
			data[43035] <= 8'h10 ;
			data[43036] <= 8'h10 ;
			data[43037] <= 8'h10 ;
			data[43038] <= 8'h10 ;
			data[43039] <= 8'h10 ;
			data[43040] <= 8'h10 ;
			data[43041] <= 8'h10 ;
			data[43042] <= 8'h10 ;
			data[43043] <= 8'h10 ;
			data[43044] <= 8'h10 ;
			data[43045] <= 8'h10 ;
			data[43046] <= 8'h10 ;
			data[43047] <= 8'h10 ;
			data[43048] <= 8'h10 ;
			data[43049] <= 8'h10 ;
			data[43050] <= 8'h10 ;
			data[43051] <= 8'h10 ;
			data[43052] <= 8'h10 ;
			data[43053] <= 8'h10 ;
			data[43054] <= 8'h10 ;
			data[43055] <= 8'h10 ;
			data[43056] <= 8'h10 ;
			data[43057] <= 8'h10 ;
			data[43058] <= 8'h10 ;
			data[43059] <= 8'h10 ;
			data[43060] <= 8'h10 ;
			data[43061] <= 8'h10 ;
			data[43062] <= 8'h10 ;
			data[43063] <= 8'h10 ;
			data[43064] <= 8'h10 ;
			data[43065] <= 8'h10 ;
			data[43066] <= 8'h10 ;
			data[43067] <= 8'h10 ;
			data[43068] <= 8'h10 ;
			data[43069] <= 8'h10 ;
			data[43070] <= 8'h10 ;
			data[43071] <= 8'h10 ;
			data[43072] <= 8'h10 ;
			data[43073] <= 8'h10 ;
			data[43074] <= 8'h10 ;
			data[43075] <= 8'h10 ;
			data[43076] <= 8'h10 ;
			data[43077] <= 8'h10 ;
			data[43078] <= 8'h10 ;
			data[43079] <= 8'h10 ;
			data[43080] <= 8'h10 ;
			data[43081] <= 8'h10 ;
			data[43082] <= 8'h10 ;
			data[43083] <= 8'h10 ;
			data[43084] <= 8'h10 ;
			data[43085] <= 8'h10 ;
			data[43086] <= 8'h10 ;
			data[43087] <= 8'h10 ;
			data[43088] <= 8'h10 ;
			data[43089] <= 8'h10 ;
			data[43090] <= 8'h10 ;
			data[43091] <= 8'h10 ;
			data[43092] <= 8'h10 ;
			data[43093] <= 8'h10 ;
			data[43094] <= 8'h10 ;
			data[43095] <= 8'h10 ;
			data[43096] <= 8'h10 ;
			data[43097] <= 8'h10 ;
			data[43098] <= 8'h10 ;
			data[43099] <= 8'h10 ;
			data[43100] <= 8'h10 ;
			data[43101] <= 8'h10 ;
			data[43102] <= 8'h10 ;
			data[43103] <= 8'h10 ;
			data[43104] <= 8'h10 ;
			data[43105] <= 8'h10 ;
			data[43106] <= 8'h10 ;
			data[43107] <= 8'h10 ;
			data[43108] <= 8'h10 ;
			data[43109] <= 8'h10 ;
			data[43110] <= 8'h10 ;
			data[43111] <= 8'h10 ;
			data[43112] <= 8'h10 ;
			data[43113] <= 8'h10 ;
			data[43114] <= 8'h10 ;
			data[43115] <= 8'h10 ;
			data[43116] <= 8'h10 ;
			data[43117] <= 8'h10 ;
			data[43118] <= 8'h10 ;
			data[43119] <= 8'h10 ;
			data[43120] <= 8'h10 ;
			data[43121] <= 8'h10 ;
			data[43122] <= 8'h10 ;
			data[43123] <= 8'h10 ;
			data[43124] <= 8'h10 ;
			data[43125] <= 8'h10 ;
			data[43126] <= 8'h10 ;
			data[43127] <= 8'h10 ;
			data[43128] <= 8'h10 ;
			data[43129] <= 8'h10 ;
			data[43130] <= 8'h10 ;
			data[43131] <= 8'h10 ;
			data[43132] <= 8'h10 ;
			data[43133] <= 8'h10 ;
			data[43134] <= 8'h10 ;
			data[43135] <= 8'h10 ;
			data[43136] <= 8'h10 ;
			data[43137] <= 8'h10 ;
			data[43138] <= 8'h10 ;
			data[43139] <= 8'h10 ;
			data[43140] <= 8'h10 ;
			data[43141] <= 8'h10 ;
			data[43142] <= 8'h10 ;
			data[43143] <= 8'h10 ;
			data[43144] <= 8'h10 ;
			data[43145] <= 8'h10 ;
			data[43146] <= 8'h10 ;
			data[43147] <= 8'h10 ;
			data[43148] <= 8'h10 ;
			data[43149] <= 8'h10 ;
			data[43150] <= 8'h10 ;
			data[43151] <= 8'h10 ;
			data[43152] <= 8'h10 ;
			data[43153] <= 8'h10 ;
			data[43154] <= 8'h10 ;
			data[43155] <= 8'h10 ;
			data[43156] <= 8'h10 ;
			data[43157] <= 8'h10 ;
			data[43158] <= 8'h10 ;
			data[43159] <= 8'h10 ;
			data[43160] <= 8'h10 ;
			data[43161] <= 8'h10 ;
			data[43162] <= 8'h10 ;
			data[43163] <= 8'h10 ;
			data[43164] <= 8'h10 ;
			data[43165] <= 8'h10 ;
			data[43166] <= 8'h10 ;
			data[43167] <= 8'h10 ;
			data[43168] <= 8'h10 ;
			data[43169] <= 8'h10 ;
			data[43170] <= 8'h10 ;
			data[43171] <= 8'h10 ;
			data[43172] <= 8'h10 ;
			data[43173] <= 8'h10 ;
			data[43174] <= 8'h10 ;
			data[43175] <= 8'h10 ;
			data[43176] <= 8'h10 ;
			data[43177] <= 8'h10 ;
			data[43178] <= 8'h10 ;
			data[43179] <= 8'h10 ;
			data[43180] <= 8'h10 ;
			data[43181] <= 8'h10 ;
			data[43182] <= 8'h10 ;
			data[43183] <= 8'h10 ;
			data[43184] <= 8'h10 ;
			data[43185] <= 8'h10 ;
			data[43186] <= 8'h10 ;
			data[43187] <= 8'h10 ;
			data[43188] <= 8'h10 ;
			data[43189] <= 8'h10 ;
			data[43190] <= 8'h10 ;
			data[43191] <= 8'h10 ;
			data[43192] <= 8'h10 ;
			data[43193] <= 8'h10 ;
			data[43194] <= 8'h10 ;
			data[43195] <= 8'h10 ;
			data[43196] <= 8'h10 ;
			data[43197] <= 8'h10 ;
			data[43198] <= 8'h10 ;
			data[43199] <= 8'h10 ;
			data[43200] <= 8'h10 ;
			data[43201] <= 8'h10 ;
			data[43202] <= 8'h10 ;
			data[43203] <= 8'h10 ;
			data[43204] <= 8'h10 ;
			data[43205] <= 8'h10 ;
			data[43206] <= 8'h10 ;
			data[43207] <= 8'h10 ;
			data[43208] <= 8'h10 ;
			data[43209] <= 8'h10 ;
			data[43210] <= 8'h10 ;
			data[43211] <= 8'h10 ;
			data[43212] <= 8'h10 ;
			data[43213] <= 8'h10 ;
			data[43214] <= 8'h10 ;
			data[43215] <= 8'h10 ;
			data[43216] <= 8'h10 ;
			data[43217] <= 8'h10 ;
			data[43218] <= 8'h10 ;
			data[43219] <= 8'h10 ;
			data[43220] <= 8'h10 ;
			data[43221] <= 8'h10 ;
			data[43222] <= 8'h10 ;
			data[43223] <= 8'h10 ;
			data[43224] <= 8'h10 ;
			data[43225] <= 8'h10 ;
			data[43226] <= 8'h10 ;
			data[43227] <= 8'h10 ;
			data[43228] <= 8'h10 ;
			data[43229] <= 8'h10 ;
			data[43230] <= 8'h10 ;
			data[43231] <= 8'h10 ;
			data[43232] <= 8'h10 ;
			data[43233] <= 8'h10 ;
			data[43234] <= 8'h10 ;
			data[43235] <= 8'h10 ;
			data[43236] <= 8'h10 ;
			data[43237] <= 8'h10 ;
			data[43238] <= 8'h10 ;
			data[43239] <= 8'h10 ;
			data[43240] <= 8'h10 ;
			data[43241] <= 8'h10 ;
			data[43242] <= 8'h10 ;
			data[43243] <= 8'h10 ;
			data[43244] <= 8'h10 ;
			data[43245] <= 8'h10 ;
			data[43246] <= 8'h10 ;
			data[43247] <= 8'h10 ;
			data[43248] <= 8'h10 ;
			data[43249] <= 8'h10 ;
			data[43250] <= 8'h10 ;
			data[43251] <= 8'h10 ;
			data[43252] <= 8'h10 ;
			data[43253] <= 8'h10 ;
			data[43254] <= 8'h10 ;
			data[43255] <= 8'h10 ;
			data[43256] <= 8'h10 ;
			data[43257] <= 8'h10 ;
			data[43258] <= 8'h10 ;
			data[43259] <= 8'h10 ;
			data[43260] <= 8'h10 ;
			data[43261] <= 8'h10 ;
			data[43262] <= 8'h10 ;
			data[43263] <= 8'h10 ;
			data[43264] <= 8'h10 ;
			data[43265] <= 8'h10 ;
			data[43266] <= 8'h10 ;
			data[43267] <= 8'h10 ;
			data[43268] <= 8'h10 ;
			data[43269] <= 8'h10 ;
			data[43270] <= 8'h10 ;
			data[43271] <= 8'h10 ;
			data[43272] <= 8'h10 ;
			data[43273] <= 8'h10 ;
			data[43274] <= 8'h10 ;
			data[43275] <= 8'h10 ;
			data[43276] <= 8'h10 ;
			data[43277] <= 8'h10 ;
			data[43278] <= 8'h10 ;
			data[43279] <= 8'h10 ;
			data[43280] <= 8'h10 ;
			data[43281] <= 8'h10 ;
			data[43282] <= 8'h10 ;
			data[43283] <= 8'h10 ;
			data[43284] <= 8'h10 ;
			data[43285] <= 8'h10 ;
			data[43286] <= 8'h10 ;
			data[43287] <= 8'h10 ;
			data[43288] <= 8'h10 ;
			data[43289] <= 8'h10 ;
			data[43290] <= 8'h10 ;
			data[43291] <= 8'h10 ;
			data[43292] <= 8'h10 ;
			data[43293] <= 8'h10 ;
			data[43294] <= 8'h10 ;
			data[43295] <= 8'h10 ;
			data[43296] <= 8'h10 ;
			data[43297] <= 8'h10 ;
			data[43298] <= 8'h10 ;
			data[43299] <= 8'h10 ;
			data[43300] <= 8'h10 ;
			data[43301] <= 8'h10 ;
			data[43302] <= 8'h10 ;
			data[43303] <= 8'h10 ;
			data[43304] <= 8'h10 ;
			data[43305] <= 8'h10 ;
			data[43306] <= 8'h10 ;
			data[43307] <= 8'h10 ;
			data[43308] <= 8'h10 ;
			data[43309] <= 8'h10 ;
			data[43310] <= 8'h10 ;
			data[43311] <= 8'h10 ;
			data[43312] <= 8'h10 ;
			data[43313] <= 8'h10 ;
			data[43314] <= 8'h10 ;
			data[43315] <= 8'h10 ;
			data[43316] <= 8'h10 ;
			data[43317] <= 8'h10 ;
			data[43318] <= 8'h10 ;
			data[43319] <= 8'h10 ;
			data[43320] <= 8'h10 ;
			data[43321] <= 8'h10 ;
			data[43322] <= 8'h10 ;
			data[43323] <= 8'h10 ;
			data[43324] <= 8'h10 ;
			data[43325] <= 8'h10 ;
			data[43326] <= 8'h10 ;
			data[43327] <= 8'h10 ;
			data[43328] <= 8'h10 ;
			data[43329] <= 8'h10 ;
			data[43330] <= 8'h10 ;
			data[43331] <= 8'h10 ;
			data[43332] <= 8'h10 ;
			data[43333] <= 8'h10 ;
			data[43334] <= 8'h10 ;
			data[43335] <= 8'h10 ;
			data[43336] <= 8'h10 ;
			data[43337] <= 8'h10 ;
			data[43338] <= 8'h10 ;
			data[43339] <= 8'h10 ;
			data[43340] <= 8'h10 ;
			data[43341] <= 8'h10 ;
			data[43342] <= 8'h10 ;
			data[43343] <= 8'h10 ;
			data[43344] <= 8'h10 ;
			data[43345] <= 8'h10 ;
			data[43346] <= 8'h10 ;
			data[43347] <= 8'h10 ;
			data[43348] <= 8'h10 ;
			data[43349] <= 8'h10 ;
			data[43350] <= 8'h10 ;
			data[43351] <= 8'h10 ;
			data[43352] <= 8'h10 ;
			data[43353] <= 8'h10 ;
			data[43354] <= 8'h10 ;
			data[43355] <= 8'h10 ;
			data[43356] <= 8'h10 ;
			data[43357] <= 8'h10 ;
			data[43358] <= 8'h10 ;
			data[43359] <= 8'h10 ;
			data[43360] <= 8'h10 ;
			data[43361] <= 8'h10 ;
			data[43362] <= 8'h10 ;
			data[43363] <= 8'h10 ;
			data[43364] <= 8'h10 ;
			data[43365] <= 8'h10 ;
			data[43366] <= 8'h10 ;
			data[43367] <= 8'h10 ;
			data[43368] <= 8'h10 ;
			data[43369] <= 8'h10 ;
			data[43370] <= 8'h10 ;
			data[43371] <= 8'h10 ;
			data[43372] <= 8'h10 ;
			data[43373] <= 8'h10 ;
			data[43374] <= 8'h10 ;
			data[43375] <= 8'h10 ;
			data[43376] <= 8'h10 ;
			data[43377] <= 8'h10 ;
			data[43378] <= 8'h10 ;
			data[43379] <= 8'h10 ;
			data[43380] <= 8'h10 ;
			data[43381] <= 8'h10 ;
			data[43382] <= 8'h10 ;
			data[43383] <= 8'h10 ;
			data[43384] <= 8'h10 ;
			data[43385] <= 8'h10 ;
			data[43386] <= 8'h10 ;
			data[43387] <= 8'h10 ;
			data[43388] <= 8'h10 ;
			data[43389] <= 8'h10 ;
			data[43390] <= 8'h10 ;
			data[43391] <= 8'h10 ;
			data[43392] <= 8'h10 ;
			data[43393] <= 8'h10 ;
			data[43394] <= 8'h10 ;
			data[43395] <= 8'h10 ;
			data[43396] <= 8'h10 ;
			data[43397] <= 8'h10 ;
			data[43398] <= 8'h10 ;
			data[43399] <= 8'h10 ;
			data[43400] <= 8'h10 ;
			data[43401] <= 8'h10 ;
			data[43402] <= 8'h10 ;
			data[43403] <= 8'h10 ;
			data[43404] <= 8'h10 ;
			data[43405] <= 8'h10 ;
			data[43406] <= 8'h10 ;
			data[43407] <= 8'h10 ;
			data[43408] <= 8'h10 ;
			data[43409] <= 8'h10 ;
			data[43410] <= 8'h10 ;
			data[43411] <= 8'h10 ;
			data[43412] <= 8'h10 ;
			data[43413] <= 8'h10 ;
			data[43414] <= 8'h10 ;
			data[43415] <= 8'h10 ;
			data[43416] <= 8'h10 ;
			data[43417] <= 8'h10 ;
			data[43418] <= 8'h10 ;
			data[43419] <= 8'h10 ;
			data[43420] <= 8'h10 ;
			data[43421] <= 8'h10 ;
			data[43422] <= 8'h10 ;
			data[43423] <= 8'h10 ;
			data[43424] <= 8'h10 ;
			data[43425] <= 8'h10 ;
			data[43426] <= 8'h10 ;
			data[43427] <= 8'h10 ;
			data[43428] <= 8'h10 ;
			data[43429] <= 8'h10 ;
			data[43430] <= 8'h10 ;
			data[43431] <= 8'h10 ;
			data[43432] <= 8'h10 ;
			data[43433] <= 8'h10 ;
			data[43434] <= 8'h10 ;
			data[43435] <= 8'h10 ;
			data[43436] <= 8'h10 ;
			data[43437] <= 8'h10 ;
			data[43438] <= 8'h10 ;
			data[43439] <= 8'h10 ;
			data[43440] <= 8'h10 ;
			data[43441] <= 8'h10 ;
			data[43442] <= 8'h10 ;
			data[43443] <= 8'h10 ;
			data[43444] <= 8'h10 ;
			data[43445] <= 8'h10 ;
			data[43446] <= 8'h10 ;
			data[43447] <= 8'h10 ;
			data[43448] <= 8'h10 ;
			data[43449] <= 8'h10 ;
			data[43450] <= 8'h10 ;
			data[43451] <= 8'h10 ;
			data[43452] <= 8'h10 ;
			data[43453] <= 8'h10 ;
			data[43454] <= 8'h10 ;
			data[43455] <= 8'h10 ;
			data[43456] <= 8'h10 ;
			data[43457] <= 8'h10 ;
			data[43458] <= 8'h10 ;
			data[43459] <= 8'h10 ;
			data[43460] <= 8'h10 ;
			data[43461] <= 8'h10 ;
			data[43462] <= 8'h10 ;
			data[43463] <= 8'h10 ;
			data[43464] <= 8'h10 ;
			data[43465] <= 8'h10 ;
			data[43466] <= 8'h10 ;
			data[43467] <= 8'h10 ;
			data[43468] <= 8'h10 ;
			data[43469] <= 8'h10 ;
			data[43470] <= 8'h10 ;
			data[43471] <= 8'h10 ;
			data[43472] <= 8'h10 ;
			data[43473] <= 8'h10 ;
			data[43474] <= 8'h10 ;
			data[43475] <= 8'h10 ;
			data[43476] <= 8'h10 ;
			data[43477] <= 8'h10 ;
			data[43478] <= 8'h10 ;
			data[43479] <= 8'h10 ;
			data[43480] <= 8'h10 ;
			data[43481] <= 8'h10 ;
			data[43482] <= 8'h10 ;
			data[43483] <= 8'h10 ;
			data[43484] <= 8'h10 ;
			data[43485] <= 8'h10 ;
			data[43486] <= 8'h10 ;
			data[43487] <= 8'h10 ;
			data[43488] <= 8'h10 ;
			data[43489] <= 8'h10 ;
			data[43490] <= 8'h10 ;
			data[43491] <= 8'h10 ;
			data[43492] <= 8'h10 ;
			data[43493] <= 8'h10 ;
			data[43494] <= 8'h10 ;
			data[43495] <= 8'h10 ;
			data[43496] <= 8'h10 ;
			data[43497] <= 8'h10 ;
			data[43498] <= 8'h10 ;
			data[43499] <= 8'h10 ;
			data[43500] <= 8'h10 ;
			data[43501] <= 8'h10 ;
			data[43502] <= 8'h10 ;
			data[43503] <= 8'h10 ;
			data[43504] <= 8'h10 ;
			data[43505] <= 8'h10 ;
			data[43506] <= 8'h10 ;
			data[43507] <= 8'h10 ;
			data[43508] <= 8'h10 ;
			data[43509] <= 8'h10 ;
			data[43510] <= 8'h10 ;
			data[43511] <= 8'h10 ;
			data[43512] <= 8'h10 ;
			data[43513] <= 8'h10 ;
			data[43514] <= 8'h10 ;
			data[43515] <= 8'h10 ;
			data[43516] <= 8'h10 ;
			data[43517] <= 8'h10 ;
			data[43518] <= 8'h10 ;
			data[43519] <= 8'h10 ;
			data[43520] <= 8'h10 ;
			data[43521] <= 8'h10 ;
			data[43522] <= 8'h10 ;
			data[43523] <= 8'h10 ;
			data[43524] <= 8'h10 ;
			data[43525] <= 8'h10 ;
			data[43526] <= 8'h10 ;
			data[43527] <= 8'h10 ;
			data[43528] <= 8'h10 ;
			data[43529] <= 8'h10 ;
			data[43530] <= 8'h10 ;
			data[43531] <= 8'h10 ;
			data[43532] <= 8'h10 ;
			data[43533] <= 8'h10 ;
			data[43534] <= 8'h10 ;
			data[43535] <= 8'h10 ;
			data[43536] <= 8'h10 ;
			data[43537] <= 8'h10 ;
			data[43538] <= 8'h10 ;
			data[43539] <= 8'h10 ;
			data[43540] <= 8'h10 ;
			data[43541] <= 8'h10 ;
			data[43542] <= 8'h10 ;
			data[43543] <= 8'h10 ;
			data[43544] <= 8'h10 ;
			data[43545] <= 8'h10 ;
			data[43546] <= 8'h10 ;
			data[43547] <= 8'h10 ;
			data[43548] <= 8'h10 ;
			data[43549] <= 8'h10 ;
			data[43550] <= 8'h10 ;
			data[43551] <= 8'h10 ;
			data[43552] <= 8'h10 ;
			data[43553] <= 8'h10 ;
			data[43554] <= 8'h10 ;
			data[43555] <= 8'h10 ;
			data[43556] <= 8'h10 ;
			data[43557] <= 8'h10 ;
			data[43558] <= 8'h10 ;
			data[43559] <= 8'h10 ;
			data[43560] <= 8'h10 ;
			data[43561] <= 8'h10 ;
			data[43562] <= 8'h10 ;
			data[43563] <= 8'h10 ;
			data[43564] <= 8'h10 ;
			data[43565] <= 8'h10 ;
			data[43566] <= 8'h10 ;
			data[43567] <= 8'h10 ;
			data[43568] <= 8'h10 ;
			data[43569] <= 8'h10 ;
			data[43570] <= 8'h10 ;
			data[43571] <= 8'h10 ;
			data[43572] <= 8'h10 ;
			data[43573] <= 8'h10 ;
			data[43574] <= 8'h10 ;
			data[43575] <= 8'h10 ;
			data[43576] <= 8'h10 ;
			data[43577] <= 8'h10 ;
			data[43578] <= 8'h10 ;
			data[43579] <= 8'h10 ;
			data[43580] <= 8'h10 ;
			data[43581] <= 8'h10 ;
			data[43582] <= 8'h10 ;
			data[43583] <= 8'h10 ;
			data[43584] <= 8'h10 ;
			data[43585] <= 8'h10 ;
			data[43586] <= 8'h10 ;
			data[43587] <= 8'h10 ;
			data[43588] <= 8'h10 ;
			data[43589] <= 8'h10 ;
			data[43590] <= 8'h10 ;
			data[43591] <= 8'h10 ;
			data[43592] <= 8'h10 ;
			data[43593] <= 8'h10 ;
			data[43594] <= 8'h10 ;
			data[43595] <= 8'h10 ;
			data[43596] <= 8'h10 ;
			data[43597] <= 8'h10 ;
			data[43598] <= 8'h10 ;
			data[43599] <= 8'h10 ;
			data[43600] <= 8'h10 ;
			data[43601] <= 8'h10 ;
			data[43602] <= 8'h10 ;
			data[43603] <= 8'h10 ;
			data[43604] <= 8'h10 ;
			data[43605] <= 8'h10 ;
			data[43606] <= 8'h10 ;
			data[43607] <= 8'h10 ;
			data[43608] <= 8'h10 ;
			data[43609] <= 8'h10 ;
			data[43610] <= 8'h10 ;
			data[43611] <= 8'h10 ;
			data[43612] <= 8'h10 ;
			data[43613] <= 8'h10 ;
			data[43614] <= 8'h10 ;
			data[43615] <= 8'h10 ;
			data[43616] <= 8'h10 ;
			data[43617] <= 8'h10 ;
			data[43618] <= 8'h10 ;
			data[43619] <= 8'h10 ;
			data[43620] <= 8'h10 ;
			data[43621] <= 8'h10 ;
			data[43622] <= 8'h10 ;
			data[43623] <= 8'h10 ;
			data[43624] <= 8'h10 ;
			data[43625] <= 8'h10 ;
			data[43626] <= 8'h10 ;
			data[43627] <= 8'h10 ;
			data[43628] <= 8'h10 ;
			data[43629] <= 8'h10 ;
			data[43630] <= 8'h10 ;
			data[43631] <= 8'h10 ;
			data[43632] <= 8'h10 ;
			data[43633] <= 8'h10 ;
			data[43634] <= 8'h10 ;
			data[43635] <= 8'h10 ;
			data[43636] <= 8'h10 ;
			data[43637] <= 8'h10 ;
			data[43638] <= 8'h10 ;
			data[43639] <= 8'h10 ;
			data[43640] <= 8'h10 ;
			data[43641] <= 8'h10 ;
			data[43642] <= 8'h10 ;
			data[43643] <= 8'h10 ;
			data[43644] <= 8'h10 ;
			data[43645] <= 8'h10 ;
			data[43646] <= 8'h10 ;
			data[43647] <= 8'h10 ;
			data[43648] <= 8'h10 ;
			data[43649] <= 8'h10 ;
			data[43650] <= 8'h10 ;
			data[43651] <= 8'h10 ;
			data[43652] <= 8'h10 ;
			data[43653] <= 8'h10 ;
			data[43654] <= 8'h10 ;
			data[43655] <= 8'h10 ;
			data[43656] <= 8'h10 ;
			data[43657] <= 8'h10 ;
			data[43658] <= 8'h10 ;
			data[43659] <= 8'h10 ;
			data[43660] <= 8'h10 ;
			data[43661] <= 8'h10 ;
			data[43662] <= 8'h10 ;
			data[43663] <= 8'h10 ;
			data[43664] <= 8'h10 ;
			data[43665] <= 8'h10 ;
			data[43666] <= 8'h10 ;
			data[43667] <= 8'h10 ;
			data[43668] <= 8'h10 ;
			data[43669] <= 8'h10 ;
			data[43670] <= 8'h10 ;
			data[43671] <= 8'h10 ;
			data[43672] <= 8'h10 ;
			data[43673] <= 8'h10 ;
			data[43674] <= 8'h10 ;
			data[43675] <= 8'h10 ;
			data[43676] <= 8'h10 ;
			data[43677] <= 8'h10 ;
			data[43678] <= 8'h10 ;
			data[43679] <= 8'h10 ;
			data[43680] <= 8'h10 ;
			data[43681] <= 8'h10 ;
			data[43682] <= 8'h10 ;
			data[43683] <= 8'h10 ;
			data[43684] <= 8'h10 ;
			data[43685] <= 8'h10 ;
			data[43686] <= 8'h10 ;
			data[43687] <= 8'h10 ;
			data[43688] <= 8'h10 ;
			data[43689] <= 8'h10 ;
			data[43690] <= 8'h10 ;
			data[43691] <= 8'h10 ;
			data[43692] <= 8'h10 ;
			data[43693] <= 8'h10 ;
			data[43694] <= 8'h10 ;
			data[43695] <= 8'h10 ;
			data[43696] <= 8'h10 ;
			data[43697] <= 8'h10 ;
			data[43698] <= 8'h10 ;
			data[43699] <= 8'h10 ;
			data[43700] <= 8'h10 ;
			data[43701] <= 8'h10 ;
			data[43702] <= 8'h10 ;
			data[43703] <= 8'h10 ;
			data[43704] <= 8'h10 ;
			data[43705] <= 8'h10 ;
			data[43706] <= 8'h10 ;
			data[43707] <= 8'h10 ;
			data[43708] <= 8'h10 ;
			data[43709] <= 8'h10 ;
			data[43710] <= 8'h10 ;
			data[43711] <= 8'h10 ;
			data[43712] <= 8'h10 ;
			data[43713] <= 8'h10 ;
			data[43714] <= 8'h10 ;
			data[43715] <= 8'h10 ;
			data[43716] <= 8'h10 ;
			data[43717] <= 8'h10 ;
			data[43718] <= 8'h10 ;
			data[43719] <= 8'h10 ;
			data[43720] <= 8'h10 ;
			data[43721] <= 8'h10 ;
			data[43722] <= 8'h10 ;
			data[43723] <= 8'h10 ;
			data[43724] <= 8'h10 ;
			data[43725] <= 8'h10 ;
			data[43726] <= 8'h10 ;
			data[43727] <= 8'h10 ;
			data[43728] <= 8'h10 ;
			data[43729] <= 8'h10 ;
			data[43730] <= 8'h10 ;
			data[43731] <= 8'h10 ;
			data[43732] <= 8'h10 ;
			data[43733] <= 8'h10 ;
			data[43734] <= 8'h10 ;
			data[43735] <= 8'h10 ;
			data[43736] <= 8'h10 ;
			data[43737] <= 8'h10 ;
			data[43738] <= 8'h10 ;
			data[43739] <= 8'h10 ;
			data[43740] <= 8'h10 ;
			data[43741] <= 8'h10 ;
			data[43742] <= 8'h10 ;
			data[43743] <= 8'h10 ;
			data[43744] <= 8'h10 ;
			data[43745] <= 8'h10 ;
			data[43746] <= 8'h10 ;
			data[43747] <= 8'h10 ;
			data[43748] <= 8'h10 ;
			data[43749] <= 8'h10 ;
			data[43750] <= 8'h10 ;
			data[43751] <= 8'h10 ;
			data[43752] <= 8'h10 ;
			data[43753] <= 8'h10 ;
			data[43754] <= 8'h10 ;
			data[43755] <= 8'h10 ;
			data[43756] <= 8'h10 ;
			data[43757] <= 8'h10 ;
			data[43758] <= 8'h10 ;
			data[43759] <= 8'h10 ;
			data[43760] <= 8'h10 ;
			data[43761] <= 8'h10 ;
			data[43762] <= 8'h10 ;
			data[43763] <= 8'h10 ;
			data[43764] <= 8'h10 ;
			data[43765] <= 8'h10 ;
			data[43766] <= 8'h10 ;
			data[43767] <= 8'h10 ;
			data[43768] <= 8'h10 ;
			data[43769] <= 8'h10 ;
			data[43770] <= 8'h10 ;
			data[43771] <= 8'h10 ;
			data[43772] <= 8'h10 ;
			data[43773] <= 8'h10 ;
			data[43774] <= 8'h10 ;
			data[43775] <= 8'h10 ;
			data[43776] <= 8'h10 ;
			data[43777] <= 8'h10 ;
			data[43778] <= 8'h10 ;
			data[43779] <= 8'h10 ;
			data[43780] <= 8'h10 ;
			data[43781] <= 8'h10 ;
			data[43782] <= 8'h10 ;
			data[43783] <= 8'h10 ;
			data[43784] <= 8'h10 ;
			data[43785] <= 8'h10 ;
			data[43786] <= 8'h10 ;
			data[43787] <= 8'h10 ;
			data[43788] <= 8'h10 ;
			data[43789] <= 8'h10 ;
			data[43790] <= 8'h10 ;
			data[43791] <= 8'h10 ;
			data[43792] <= 8'h10 ;
			data[43793] <= 8'h10 ;
			data[43794] <= 8'h10 ;
			data[43795] <= 8'h10 ;
			data[43796] <= 8'h10 ;
			data[43797] <= 8'h10 ;
			data[43798] <= 8'h10 ;
			data[43799] <= 8'h10 ;
			data[43800] <= 8'h10 ;
			data[43801] <= 8'h10 ;
			data[43802] <= 8'h10 ;
			data[43803] <= 8'h10 ;
			data[43804] <= 8'h10 ;
			data[43805] <= 8'h10 ;
			data[43806] <= 8'h10 ;
			data[43807] <= 8'h10 ;
			data[43808] <= 8'h10 ;
			data[43809] <= 8'h10 ;
			data[43810] <= 8'h10 ;
			data[43811] <= 8'h10 ;
			data[43812] <= 8'h10 ;
			data[43813] <= 8'h10 ;
			data[43814] <= 8'h10 ;
			data[43815] <= 8'h10 ;
			data[43816] <= 8'h10 ;
			data[43817] <= 8'h10 ;
			data[43818] <= 8'h10 ;
			data[43819] <= 8'h10 ;
			data[43820] <= 8'h10 ;
			data[43821] <= 8'h10 ;
			data[43822] <= 8'h10 ;
			data[43823] <= 8'h10 ;
			data[43824] <= 8'h10 ;
			data[43825] <= 8'h10 ;
			data[43826] <= 8'h10 ;
			data[43827] <= 8'h10 ;
			data[43828] <= 8'h10 ;
			data[43829] <= 8'h10 ;
			data[43830] <= 8'h10 ;
			data[43831] <= 8'h10 ;
			data[43832] <= 8'h10 ;
			data[43833] <= 8'h10 ;
			data[43834] <= 8'h10 ;
			data[43835] <= 8'h10 ;
			data[43836] <= 8'h10 ;
			data[43837] <= 8'h10 ;
			data[43838] <= 8'h10 ;
			data[43839] <= 8'h10 ;
			data[43840] <= 8'h10 ;
			data[43841] <= 8'h10 ;
			data[43842] <= 8'h10 ;
			data[43843] <= 8'h10 ;
			data[43844] <= 8'h10 ;
			data[43845] <= 8'h10 ;
			data[43846] <= 8'h10 ;
			data[43847] <= 8'h10 ;
			data[43848] <= 8'h10 ;
			data[43849] <= 8'h10 ;
			data[43850] <= 8'h10 ;
			data[43851] <= 8'h10 ;
			data[43852] <= 8'h10 ;
			data[43853] <= 8'h10 ;
			data[43854] <= 8'h10 ;
			data[43855] <= 8'h10 ;
			data[43856] <= 8'h10 ;
			data[43857] <= 8'h10 ;
			data[43858] <= 8'h10 ;
			data[43859] <= 8'h10 ;
			data[43860] <= 8'h10 ;
			data[43861] <= 8'h10 ;
			data[43862] <= 8'h10 ;
			data[43863] <= 8'h10 ;
			data[43864] <= 8'h10 ;
			data[43865] <= 8'h10 ;
			data[43866] <= 8'h10 ;
			data[43867] <= 8'h10 ;
			data[43868] <= 8'h10 ;
			data[43869] <= 8'h10 ;
			data[43870] <= 8'h10 ;
			data[43871] <= 8'h10 ;
			data[43872] <= 8'h10 ;
			data[43873] <= 8'h10 ;
			data[43874] <= 8'h10 ;
			data[43875] <= 8'h10 ;
			data[43876] <= 8'h10 ;
			data[43877] <= 8'h10 ;
			data[43878] <= 8'h10 ;
			data[43879] <= 8'h10 ;
			data[43880] <= 8'h10 ;
			data[43881] <= 8'h10 ;
			data[43882] <= 8'h10 ;
			data[43883] <= 8'h10 ;
			data[43884] <= 8'h10 ;
			data[43885] <= 8'h10 ;
			data[43886] <= 8'h10 ;
			data[43887] <= 8'h10 ;
			data[43888] <= 8'h10 ;
			data[43889] <= 8'h10 ;
			data[43890] <= 8'h10 ;
			data[43891] <= 8'h10 ;
			data[43892] <= 8'h10 ;
			data[43893] <= 8'h10 ;
			data[43894] <= 8'h10 ;
			data[43895] <= 8'h10 ;
			data[43896] <= 8'h10 ;
			data[43897] <= 8'h10 ;
			data[43898] <= 8'h10 ;
			data[43899] <= 8'h10 ;
			data[43900] <= 8'h10 ;
			data[43901] <= 8'h10 ;
			data[43902] <= 8'h10 ;
			data[43903] <= 8'h10 ;
			data[43904] <= 8'h10 ;
			data[43905] <= 8'h10 ;
			data[43906] <= 8'h10 ;
			data[43907] <= 8'h10 ;
			data[43908] <= 8'h10 ;
			data[43909] <= 8'h10 ;
			data[43910] <= 8'h10 ;
			data[43911] <= 8'h10 ;
			data[43912] <= 8'h10 ;
			data[43913] <= 8'h10 ;
			data[43914] <= 8'h10 ;
			data[43915] <= 8'h10 ;
			data[43916] <= 8'h10 ;
			data[43917] <= 8'h10 ;
			data[43918] <= 8'h10 ;
			data[43919] <= 8'h10 ;
			data[43920] <= 8'h10 ;
			data[43921] <= 8'h10 ;
			data[43922] <= 8'h10 ;
			data[43923] <= 8'h10 ;
			data[43924] <= 8'h10 ;
			data[43925] <= 8'h10 ;
			data[43926] <= 8'h10 ;
			data[43927] <= 8'h10 ;
			data[43928] <= 8'h10 ;
			data[43929] <= 8'h10 ;
			data[43930] <= 8'h10 ;
			data[43931] <= 8'h10 ;
			data[43932] <= 8'h10 ;
			data[43933] <= 8'h10 ;
			data[43934] <= 8'h10 ;
			data[43935] <= 8'h10 ;
			data[43936] <= 8'h10 ;
			data[43937] <= 8'h10 ;
			data[43938] <= 8'h10 ;
			data[43939] <= 8'h10 ;
			data[43940] <= 8'h10 ;
			data[43941] <= 8'h10 ;
			data[43942] <= 8'h10 ;
			data[43943] <= 8'h10 ;
			data[43944] <= 8'h10 ;
			data[43945] <= 8'h10 ;
			data[43946] <= 8'h10 ;
			data[43947] <= 8'h10 ;
			data[43948] <= 8'h10 ;
			data[43949] <= 8'h10 ;
			data[43950] <= 8'h10 ;
			data[43951] <= 8'h10 ;
			data[43952] <= 8'h10 ;
			data[43953] <= 8'h10 ;
			data[43954] <= 8'h10 ;
			data[43955] <= 8'h10 ;
			data[43956] <= 8'h10 ;
			data[43957] <= 8'h10 ;
			data[43958] <= 8'h10 ;
			data[43959] <= 8'h10 ;
			data[43960] <= 8'h10 ;
			data[43961] <= 8'h10 ;
			data[43962] <= 8'h10 ;
			data[43963] <= 8'h10 ;
			data[43964] <= 8'h10 ;
			data[43965] <= 8'h10 ;
			data[43966] <= 8'h10 ;
			data[43967] <= 8'h10 ;
			data[43968] <= 8'h10 ;
			data[43969] <= 8'h10 ;
			data[43970] <= 8'h10 ;
			data[43971] <= 8'h10 ;
			data[43972] <= 8'h10 ;
			data[43973] <= 8'h10 ;
			data[43974] <= 8'h10 ;
			data[43975] <= 8'h10 ;
			data[43976] <= 8'h10 ;
			data[43977] <= 8'h10 ;
			data[43978] <= 8'h10 ;
			data[43979] <= 8'h10 ;
			data[43980] <= 8'h10 ;
			data[43981] <= 8'h10 ;
			data[43982] <= 8'h10 ;
			data[43983] <= 8'h10 ;
			data[43984] <= 8'h10 ;
			data[43985] <= 8'h10 ;
			data[43986] <= 8'h10 ;
			data[43987] <= 8'h10 ;
			data[43988] <= 8'h10 ;
			data[43989] <= 8'h10 ;
			data[43990] <= 8'h10 ;
			data[43991] <= 8'h10 ;
			data[43992] <= 8'h10 ;
			data[43993] <= 8'h10 ;
			data[43994] <= 8'h10 ;
			data[43995] <= 8'h10 ;
			data[43996] <= 8'h10 ;
			data[43997] <= 8'h10 ;
			data[43998] <= 8'h10 ;
			data[43999] <= 8'h10 ;
			data[44000] <= 8'h10 ;
			data[44001] <= 8'h10 ;
			data[44002] <= 8'h10 ;
			data[44003] <= 8'h10 ;
			data[44004] <= 8'h10 ;
			data[44005] <= 8'h10 ;
			data[44006] <= 8'h10 ;
			data[44007] <= 8'h10 ;
			data[44008] <= 8'h10 ;
			data[44009] <= 8'h10 ;
			data[44010] <= 8'h10 ;
			data[44011] <= 8'h10 ;
			data[44012] <= 8'h10 ;
			data[44013] <= 8'h10 ;
			data[44014] <= 8'h10 ;
			data[44015] <= 8'h10 ;
			data[44016] <= 8'h10 ;
			data[44017] <= 8'h10 ;
			data[44018] <= 8'h10 ;
			data[44019] <= 8'h10 ;
			data[44020] <= 8'h10 ;
			data[44021] <= 8'h10 ;
			data[44022] <= 8'h10 ;
			data[44023] <= 8'h10 ;
			data[44024] <= 8'h10 ;
			data[44025] <= 8'h10 ;
			data[44026] <= 8'h10 ;
			data[44027] <= 8'h10 ;
			data[44028] <= 8'h10 ;
			data[44029] <= 8'h10 ;
			data[44030] <= 8'h10 ;
			data[44031] <= 8'h10 ;
			data[44032] <= 8'h10 ;
			data[44033] <= 8'h10 ;
			data[44034] <= 8'h10 ;
			data[44035] <= 8'h10 ;
			data[44036] <= 8'h10 ;
			data[44037] <= 8'h10 ;
			data[44038] <= 8'h10 ;
			data[44039] <= 8'h10 ;
			data[44040] <= 8'h10 ;
			data[44041] <= 8'h10 ;
			data[44042] <= 8'h10 ;
			data[44043] <= 8'h10 ;
			data[44044] <= 8'h10 ;
			data[44045] <= 8'h10 ;
			data[44046] <= 8'h10 ;
			data[44047] <= 8'h10 ;
			data[44048] <= 8'h10 ;
			data[44049] <= 8'h10 ;
			data[44050] <= 8'h10 ;
			data[44051] <= 8'h10 ;
			data[44052] <= 8'h10 ;
			data[44053] <= 8'h10 ;
			data[44054] <= 8'h10 ;
			data[44055] <= 8'h10 ;
			data[44056] <= 8'h10 ;
			data[44057] <= 8'h10 ;
			data[44058] <= 8'h10 ;
			data[44059] <= 8'h10 ;
			data[44060] <= 8'h10 ;
			data[44061] <= 8'h10 ;
			data[44062] <= 8'h10 ;
			data[44063] <= 8'h10 ;
			data[44064] <= 8'h10 ;
			data[44065] <= 8'h10 ;
			data[44066] <= 8'h10 ;
			data[44067] <= 8'h10 ;
			data[44068] <= 8'h10 ;
			data[44069] <= 8'h10 ;
			data[44070] <= 8'h10 ;
			data[44071] <= 8'h10 ;
			data[44072] <= 8'h10 ;
			data[44073] <= 8'h10 ;
			data[44074] <= 8'h10 ;
			data[44075] <= 8'h10 ;
			data[44076] <= 8'h10 ;
			data[44077] <= 8'h10 ;
			data[44078] <= 8'h10 ;
			data[44079] <= 8'h10 ;
			data[44080] <= 8'h10 ;
			data[44081] <= 8'h10 ;
			data[44082] <= 8'h10 ;
			data[44083] <= 8'h10 ;
			data[44084] <= 8'h10 ;
			data[44085] <= 8'h10 ;
			data[44086] <= 8'h10 ;
			data[44087] <= 8'h10 ;
			data[44088] <= 8'h10 ;
			data[44089] <= 8'h10 ;
			data[44090] <= 8'h10 ;
			data[44091] <= 8'h10 ;
			data[44092] <= 8'h10 ;
			data[44093] <= 8'h10 ;
			data[44094] <= 8'h10 ;
			data[44095] <= 8'h10 ;
			data[44096] <= 8'h10 ;
			data[44097] <= 8'h10 ;
			data[44098] <= 8'h10 ;
			data[44099] <= 8'h10 ;
			data[44100] <= 8'h10 ;
			data[44101] <= 8'h10 ;
			data[44102] <= 8'h10 ;
			data[44103] <= 8'h10 ;
			data[44104] <= 8'h10 ;
			data[44105] <= 8'h10 ;
			data[44106] <= 8'h10 ;
			data[44107] <= 8'h10 ;
			data[44108] <= 8'h10 ;
			data[44109] <= 8'h10 ;
			data[44110] <= 8'h10 ;
			data[44111] <= 8'h10 ;
			data[44112] <= 8'h10 ;
			data[44113] <= 8'h10 ;
			data[44114] <= 8'h10 ;
			data[44115] <= 8'h10 ;
			data[44116] <= 8'h10 ;
			data[44117] <= 8'h10 ;
			data[44118] <= 8'h10 ;
			data[44119] <= 8'h10 ;
			data[44120] <= 8'h10 ;
			data[44121] <= 8'h10 ;
			data[44122] <= 8'h10 ;
			data[44123] <= 8'h10 ;
			data[44124] <= 8'h10 ;
			data[44125] <= 8'h10 ;
			data[44126] <= 8'h10 ;
			data[44127] <= 8'h10 ;
			data[44128] <= 8'h10 ;
			data[44129] <= 8'h10 ;
			data[44130] <= 8'h10 ;
			data[44131] <= 8'h10 ;
			data[44132] <= 8'h10 ;
			data[44133] <= 8'h10 ;
			data[44134] <= 8'h10 ;
			data[44135] <= 8'h10 ;
			data[44136] <= 8'h10 ;
			data[44137] <= 8'h10 ;
			data[44138] <= 8'h10 ;
			data[44139] <= 8'h10 ;
			data[44140] <= 8'h10 ;
			data[44141] <= 8'h10 ;
			data[44142] <= 8'h10 ;
			data[44143] <= 8'h10 ;
			data[44144] <= 8'h10 ;
			data[44145] <= 8'h10 ;
			data[44146] <= 8'h10 ;
			data[44147] <= 8'h10 ;
			data[44148] <= 8'h10 ;
			data[44149] <= 8'h10 ;
			data[44150] <= 8'h10 ;
			data[44151] <= 8'h10 ;
			data[44152] <= 8'h10 ;
			data[44153] <= 8'h10 ;
			data[44154] <= 8'h10 ;
			data[44155] <= 8'h10 ;
			data[44156] <= 8'h10 ;
			data[44157] <= 8'h10 ;
			data[44158] <= 8'h10 ;
			data[44159] <= 8'h10 ;
			data[44160] <= 8'h10 ;
			data[44161] <= 8'h10 ;
			data[44162] <= 8'h10 ;
			data[44163] <= 8'h10 ;
			data[44164] <= 8'h10 ;
			data[44165] <= 8'h10 ;
			data[44166] <= 8'h10 ;
			data[44167] <= 8'h10 ;
			data[44168] <= 8'h10 ;
			data[44169] <= 8'h10 ;
			data[44170] <= 8'h10 ;
			data[44171] <= 8'h10 ;
			data[44172] <= 8'h10 ;
			data[44173] <= 8'h10 ;
			data[44174] <= 8'h10 ;
			data[44175] <= 8'h10 ;
			data[44176] <= 8'h10 ;
			data[44177] <= 8'h10 ;
			data[44178] <= 8'h10 ;
			data[44179] <= 8'h10 ;
			data[44180] <= 8'h10 ;
			data[44181] <= 8'h10 ;
			data[44182] <= 8'h10 ;
			data[44183] <= 8'h10 ;
			data[44184] <= 8'h10 ;
			data[44185] <= 8'h10 ;
			data[44186] <= 8'h10 ;
			data[44187] <= 8'h10 ;
			data[44188] <= 8'h10 ;
			data[44189] <= 8'h10 ;
			data[44190] <= 8'h10 ;
			data[44191] <= 8'h10 ;
			data[44192] <= 8'h10 ;
			data[44193] <= 8'h10 ;
			data[44194] <= 8'h10 ;
			data[44195] <= 8'h10 ;
			data[44196] <= 8'h10 ;
			data[44197] <= 8'h10 ;
			data[44198] <= 8'h10 ;
			data[44199] <= 8'h10 ;
			data[44200] <= 8'h10 ;
			data[44201] <= 8'h10 ;
			data[44202] <= 8'h10 ;
			data[44203] <= 8'h10 ;
			data[44204] <= 8'h10 ;
			data[44205] <= 8'h10 ;
			data[44206] <= 8'h10 ;
			data[44207] <= 8'h10 ;
			data[44208] <= 8'h10 ;
			data[44209] <= 8'h10 ;
			data[44210] <= 8'h10 ;
			data[44211] <= 8'h10 ;
			data[44212] <= 8'h10 ;
			data[44213] <= 8'h10 ;
			data[44214] <= 8'h10 ;
			data[44215] <= 8'h10 ;
			data[44216] <= 8'h10 ;
			data[44217] <= 8'h10 ;
			data[44218] <= 8'h10 ;
			data[44219] <= 8'h10 ;
			data[44220] <= 8'h10 ;
			data[44221] <= 8'h10 ;
			data[44222] <= 8'h10 ;
			data[44223] <= 8'h10 ;
			data[44224] <= 8'h10 ;
			data[44225] <= 8'h10 ;
			data[44226] <= 8'h10 ;
			data[44227] <= 8'h10 ;
			data[44228] <= 8'h10 ;
			data[44229] <= 8'h10 ;
			data[44230] <= 8'h10 ;
			data[44231] <= 8'h10 ;
			data[44232] <= 8'h10 ;
			data[44233] <= 8'h10 ;
			data[44234] <= 8'h10 ;
			data[44235] <= 8'h10 ;
			data[44236] <= 8'h10 ;
			data[44237] <= 8'h10 ;
			data[44238] <= 8'h10 ;
			data[44239] <= 8'h10 ;
			data[44240] <= 8'h10 ;
			data[44241] <= 8'h10 ;
			data[44242] <= 8'h10 ;
			data[44243] <= 8'h10 ;
			data[44244] <= 8'h10 ;
			data[44245] <= 8'h10 ;
			data[44246] <= 8'h10 ;
			data[44247] <= 8'h10 ;
			data[44248] <= 8'h10 ;
			data[44249] <= 8'h10 ;
			data[44250] <= 8'h10 ;
			data[44251] <= 8'h10 ;
			data[44252] <= 8'h10 ;
			data[44253] <= 8'h10 ;
			data[44254] <= 8'h10 ;
			data[44255] <= 8'h10 ;
			data[44256] <= 8'h10 ;
			data[44257] <= 8'h10 ;
			data[44258] <= 8'h10 ;
			data[44259] <= 8'h10 ;
			data[44260] <= 8'h10 ;
			data[44261] <= 8'h10 ;
			data[44262] <= 8'h10 ;
			data[44263] <= 8'h10 ;
			data[44264] <= 8'h10 ;
			data[44265] <= 8'h10 ;
			data[44266] <= 8'h10 ;
			data[44267] <= 8'h10 ;
			data[44268] <= 8'h10 ;
			data[44269] <= 8'h10 ;
			data[44270] <= 8'h10 ;
			data[44271] <= 8'h10 ;
			data[44272] <= 8'h10 ;
			data[44273] <= 8'h10 ;
			data[44274] <= 8'h10 ;
			data[44275] <= 8'h10 ;
			data[44276] <= 8'h10 ;
			data[44277] <= 8'h10 ;
			data[44278] <= 8'h10 ;
			data[44279] <= 8'h10 ;
			data[44280] <= 8'h10 ;
			data[44281] <= 8'h10 ;
			data[44282] <= 8'h10 ;
			data[44283] <= 8'h10 ;
			data[44284] <= 8'h10 ;
			data[44285] <= 8'h10 ;
			data[44286] <= 8'h10 ;
			data[44287] <= 8'h10 ;
			data[44288] <= 8'h10 ;
			data[44289] <= 8'h10 ;
			data[44290] <= 8'h10 ;
			data[44291] <= 8'h10 ;
			data[44292] <= 8'h10 ;
			data[44293] <= 8'h10 ;
			data[44294] <= 8'h10 ;
			data[44295] <= 8'h10 ;
			data[44296] <= 8'h10 ;
			data[44297] <= 8'h10 ;
			data[44298] <= 8'h10 ;
			data[44299] <= 8'h10 ;
			data[44300] <= 8'h10 ;
			data[44301] <= 8'h10 ;
			data[44302] <= 8'h10 ;
			data[44303] <= 8'h10 ;
			data[44304] <= 8'h10 ;
			data[44305] <= 8'h10 ;
			data[44306] <= 8'h10 ;
			data[44307] <= 8'h10 ;
			data[44308] <= 8'h10 ;
			data[44309] <= 8'h10 ;
			data[44310] <= 8'h10 ;
			data[44311] <= 8'h10 ;
			data[44312] <= 8'h10 ;
			data[44313] <= 8'h10 ;
			data[44314] <= 8'h10 ;
			data[44315] <= 8'h10 ;
			data[44316] <= 8'h10 ;
			data[44317] <= 8'h10 ;
			data[44318] <= 8'h10 ;
			data[44319] <= 8'h10 ;
			data[44320] <= 8'h10 ;
			data[44321] <= 8'h10 ;
			data[44322] <= 8'h10 ;
			data[44323] <= 8'h10 ;
			data[44324] <= 8'h10 ;
			data[44325] <= 8'h10 ;
			data[44326] <= 8'h10 ;
			data[44327] <= 8'h10 ;
			data[44328] <= 8'h10 ;
			data[44329] <= 8'h10 ;
			data[44330] <= 8'h10 ;
			data[44331] <= 8'h10 ;
			data[44332] <= 8'h10 ;
			data[44333] <= 8'h10 ;
			data[44334] <= 8'h10 ;
			data[44335] <= 8'h10 ;
			data[44336] <= 8'h10 ;
			data[44337] <= 8'h10 ;
			data[44338] <= 8'h10 ;
			data[44339] <= 8'h10 ;
			data[44340] <= 8'h10 ;
			data[44341] <= 8'h10 ;
			data[44342] <= 8'h10 ;
			data[44343] <= 8'h10 ;
			data[44344] <= 8'h10 ;
			data[44345] <= 8'h10 ;
			data[44346] <= 8'h10 ;
			data[44347] <= 8'h10 ;
			data[44348] <= 8'h10 ;
			data[44349] <= 8'h10 ;
			data[44350] <= 8'h10 ;
			data[44351] <= 8'h10 ;
			data[44352] <= 8'h10 ;
			data[44353] <= 8'h10 ;
			data[44354] <= 8'h10 ;
			data[44355] <= 8'h10 ;
			data[44356] <= 8'h10 ;
			data[44357] <= 8'h10 ;
			data[44358] <= 8'h10 ;
			data[44359] <= 8'h10 ;
			data[44360] <= 8'h10 ;
			data[44361] <= 8'h10 ;
			data[44362] <= 8'h10 ;
			data[44363] <= 8'h10 ;
			data[44364] <= 8'h10 ;
			data[44365] <= 8'h10 ;
			data[44366] <= 8'h10 ;
			data[44367] <= 8'h10 ;
			data[44368] <= 8'h10 ;
			data[44369] <= 8'h10 ;
			data[44370] <= 8'h10 ;
			data[44371] <= 8'h10 ;
			data[44372] <= 8'h10 ;
			data[44373] <= 8'h10 ;
			data[44374] <= 8'h10 ;
			data[44375] <= 8'h10 ;
			data[44376] <= 8'h10 ;
			data[44377] <= 8'h10 ;
			data[44378] <= 8'h10 ;
			data[44379] <= 8'h10 ;
			data[44380] <= 8'h10 ;
			data[44381] <= 8'h10 ;
			data[44382] <= 8'h10 ;
			data[44383] <= 8'h10 ;
			data[44384] <= 8'h10 ;
			data[44385] <= 8'h10 ;
			data[44386] <= 8'h10 ;
			data[44387] <= 8'h10 ;
			data[44388] <= 8'h10 ;
			data[44389] <= 8'h10 ;
			data[44390] <= 8'h10 ;
			data[44391] <= 8'h10 ;
			data[44392] <= 8'h10 ;
			data[44393] <= 8'h10 ;
			data[44394] <= 8'h10 ;
			data[44395] <= 8'h10 ;
			data[44396] <= 8'h10 ;
			data[44397] <= 8'h10 ;
			data[44398] <= 8'h10 ;
			data[44399] <= 8'h10 ;
			data[44400] <= 8'h10 ;
			data[44401] <= 8'h10 ;
			data[44402] <= 8'h10 ;
			data[44403] <= 8'h10 ;
			data[44404] <= 8'h10 ;
			data[44405] <= 8'h10 ;
			data[44406] <= 8'h10 ;
			data[44407] <= 8'h10 ;
			data[44408] <= 8'h10 ;
			data[44409] <= 8'h10 ;
			data[44410] <= 8'h10 ;
			data[44411] <= 8'h10 ;
			data[44412] <= 8'h10 ;
			data[44413] <= 8'h10 ;
			data[44414] <= 8'h10 ;
			data[44415] <= 8'h10 ;
			data[44416] <= 8'h10 ;
			data[44417] <= 8'h10 ;
			data[44418] <= 8'h10 ;
			data[44419] <= 8'h10 ;
			data[44420] <= 8'h10 ;
			data[44421] <= 8'h10 ;
			data[44422] <= 8'h10 ;
			data[44423] <= 8'h10 ;
			data[44424] <= 8'h10 ;
			data[44425] <= 8'h10 ;
			data[44426] <= 8'h10 ;
			data[44427] <= 8'h10 ;
			data[44428] <= 8'h10 ;
			data[44429] <= 8'h10 ;
			data[44430] <= 8'h10 ;
			data[44431] <= 8'h10 ;
			data[44432] <= 8'h10 ;
			data[44433] <= 8'h10 ;
			data[44434] <= 8'h10 ;
			data[44435] <= 8'h10 ;
			data[44436] <= 8'h10 ;
			data[44437] <= 8'h10 ;
			data[44438] <= 8'h10 ;
			data[44439] <= 8'h10 ;
			data[44440] <= 8'h10 ;
			data[44441] <= 8'h10 ;
			data[44442] <= 8'h10 ;
			data[44443] <= 8'h10 ;
			data[44444] <= 8'h10 ;
			data[44445] <= 8'h10 ;
			data[44446] <= 8'h10 ;
			data[44447] <= 8'h10 ;
			data[44448] <= 8'h10 ;
			data[44449] <= 8'h10 ;
			data[44450] <= 8'h10 ;
			data[44451] <= 8'h10 ;
			data[44452] <= 8'h10 ;
			data[44453] <= 8'h10 ;
			data[44454] <= 8'h10 ;
			data[44455] <= 8'h10 ;
			data[44456] <= 8'h10 ;
			data[44457] <= 8'h10 ;
			data[44458] <= 8'h10 ;
			data[44459] <= 8'h10 ;
			data[44460] <= 8'h10 ;
			data[44461] <= 8'h10 ;
			data[44462] <= 8'h10 ;
			data[44463] <= 8'h10 ;
			data[44464] <= 8'h10 ;
			data[44465] <= 8'h10 ;
			data[44466] <= 8'h10 ;
			data[44467] <= 8'h10 ;
			data[44468] <= 8'h10 ;
			data[44469] <= 8'h10 ;
			data[44470] <= 8'h10 ;
			data[44471] <= 8'h10 ;
			data[44472] <= 8'h10 ;
			data[44473] <= 8'h10 ;
			data[44474] <= 8'h10 ;
			data[44475] <= 8'h10 ;
			data[44476] <= 8'h10 ;
			data[44477] <= 8'h10 ;
			data[44478] <= 8'h10 ;
			data[44479] <= 8'h10 ;
			data[44480] <= 8'h10 ;
			data[44481] <= 8'h10 ;
			data[44482] <= 8'h10 ;
			data[44483] <= 8'h10 ;
			data[44484] <= 8'h10 ;
			data[44485] <= 8'h10 ;
			data[44486] <= 8'h10 ;
			data[44487] <= 8'h10 ;
			data[44488] <= 8'h10 ;
			data[44489] <= 8'h10 ;
			data[44490] <= 8'h10 ;
			data[44491] <= 8'h10 ;
			data[44492] <= 8'h10 ;
			data[44493] <= 8'h10 ;
			data[44494] <= 8'h10 ;
			data[44495] <= 8'h10 ;
			data[44496] <= 8'h10 ;
			data[44497] <= 8'h10 ;
			data[44498] <= 8'h10 ;
			data[44499] <= 8'h10 ;
			data[44500] <= 8'h10 ;
			data[44501] <= 8'h10 ;
			data[44502] <= 8'h10 ;
			data[44503] <= 8'h10 ;
			data[44504] <= 8'h10 ;
			data[44505] <= 8'h10 ;
			data[44506] <= 8'h10 ;
			data[44507] <= 8'h10 ;
			data[44508] <= 8'h10 ;
			data[44509] <= 8'h10 ;
			data[44510] <= 8'h10 ;
			data[44511] <= 8'h10 ;
			data[44512] <= 8'h10 ;
			data[44513] <= 8'h10 ;
			data[44514] <= 8'h10 ;
			data[44515] <= 8'h10 ;
			data[44516] <= 8'h10 ;
			data[44517] <= 8'h10 ;
			data[44518] <= 8'h10 ;
			data[44519] <= 8'h10 ;
			data[44520] <= 8'h10 ;
			data[44521] <= 8'h10 ;
			data[44522] <= 8'h10 ;
			data[44523] <= 8'h10 ;
			data[44524] <= 8'h10 ;
			data[44525] <= 8'h10 ;
			data[44526] <= 8'h10 ;
			data[44527] <= 8'h10 ;
			data[44528] <= 8'h10 ;
			data[44529] <= 8'h10 ;
			data[44530] <= 8'h10 ;
			data[44531] <= 8'h10 ;
			data[44532] <= 8'h10 ;
			data[44533] <= 8'h10 ;
			data[44534] <= 8'h10 ;
			data[44535] <= 8'h10 ;
			data[44536] <= 8'h10 ;
			data[44537] <= 8'h10 ;
			data[44538] <= 8'h10 ;
			data[44539] <= 8'h10 ;
			data[44540] <= 8'h10 ;
			data[44541] <= 8'h10 ;
			data[44542] <= 8'h10 ;
			data[44543] <= 8'h10 ;
			data[44544] <= 8'h10 ;
			data[44545] <= 8'h10 ;
			data[44546] <= 8'h10 ;
			data[44547] <= 8'h10 ;
			data[44548] <= 8'h10 ;
			data[44549] <= 8'h10 ;
			data[44550] <= 8'h10 ;
			data[44551] <= 8'h10 ;
			data[44552] <= 8'h10 ;
			data[44553] <= 8'h10 ;
			data[44554] <= 8'h10 ;
			data[44555] <= 8'h10 ;
			data[44556] <= 8'h10 ;
			data[44557] <= 8'h10 ;
			data[44558] <= 8'h10 ;
			data[44559] <= 8'h10 ;
			data[44560] <= 8'h10 ;
			data[44561] <= 8'h10 ;
			data[44562] <= 8'h10 ;
			data[44563] <= 8'h10 ;
			data[44564] <= 8'h10 ;
			data[44565] <= 8'h10 ;
			data[44566] <= 8'h10 ;
			data[44567] <= 8'h10 ;
			data[44568] <= 8'h10 ;
			data[44569] <= 8'h10 ;
			data[44570] <= 8'h10 ;
			data[44571] <= 8'h10 ;
			data[44572] <= 8'h10 ;
			data[44573] <= 8'h10 ;
			data[44574] <= 8'h10 ;
			data[44575] <= 8'h10 ;
			data[44576] <= 8'h10 ;
			data[44577] <= 8'h10 ;
			data[44578] <= 8'h10 ;
			data[44579] <= 8'h10 ;
			data[44580] <= 8'h10 ;
			data[44581] <= 8'h10 ;
			data[44582] <= 8'h10 ;
			data[44583] <= 8'h10 ;
			data[44584] <= 8'h10 ;
			data[44585] <= 8'h10 ;
			data[44586] <= 8'h10 ;
			data[44587] <= 8'h10 ;
			data[44588] <= 8'h10 ;
			data[44589] <= 8'h10 ;
			data[44590] <= 8'h10 ;
			data[44591] <= 8'h10 ;
			data[44592] <= 8'h10 ;
			data[44593] <= 8'h10 ;
			data[44594] <= 8'h10 ;
			data[44595] <= 8'h10 ;
			data[44596] <= 8'h10 ;
			data[44597] <= 8'h10 ;
			data[44598] <= 8'h10 ;
			data[44599] <= 8'h10 ;
			data[44600] <= 8'h10 ;
			data[44601] <= 8'h10 ;
			data[44602] <= 8'h10 ;
			data[44603] <= 8'h10 ;
			data[44604] <= 8'h10 ;
			data[44605] <= 8'h10 ;
			data[44606] <= 8'h10 ;
			data[44607] <= 8'h10 ;
			data[44608] <= 8'h10 ;
			data[44609] <= 8'h10 ;
			data[44610] <= 8'h10 ;
			data[44611] <= 8'h10 ;
			data[44612] <= 8'h10 ;
			data[44613] <= 8'h10 ;
			data[44614] <= 8'h10 ;
			data[44615] <= 8'h10 ;
			data[44616] <= 8'h10 ;
			data[44617] <= 8'h10 ;
			data[44618] <= 8'h10 ;
			data[44619] <= 8'h10 ;
			data[44620] <= 8'h10 ;
			data[44621] <= 8'h10 ;
			data[44622] <= 8'h10 ;
			data[44623] <= 8'h10 ;
			data[44624] <= 8'h10 ;
			data[44625] <= 8'h10 ;
			data[44626] <= 8'h10 ;
			data[44627] <= 8'h10 ;
			data[44628] <= 8'h10 ;
			data[44629] <= 8'h10 ;
			data[44630] <= 8'h10 ;
			data[44631] <= 8'h10 ;
			data[44632] <= 8'h10 ;
			data[44633] <= 8'h10 ;
			data[44634] <= 8'h10 ;
			data[44635] <= 8'h10 ;
			data[44636] <= 8'h10 ;
			data[44637] <= 8'h10 ;
			data[44638] <= 8'h10 ;
			data[44639] <= 8'h10 ;
			data[44640] <= 8'h10 ;
			data[44641] <= 8'h10 ;
			data[44642] <= 8'h10 ;
			data[44643] <= 8'h10 ;
			data[44644] <= 8'h10 ;
			data[44645] <= 8'h10 ;
			data[44646] <= 8'h10 ;
			data[44647] <= 8'h10 ;
			data[44648] <= 8'h10 ;
			data[44649] <= 8'h10 ;
			data[44650] <= 8'h10 ;
			data[44651] <= 8'h10 ;
			data[44652] <= 8'h10 ;
			data[44653] <= 8'h10 ;
			data[44654] <= 8'h10 ;
			data[44655] <= 8'h10 ;
			data[44656] <= 8'h10 ;
			data[44657] <= 8'h10 ;
			data[44658] <= 8'h10 ;
			data[44659] <= 8'h10 ;
			data[44660] <= 8'h10 ;
			data[44661] <= 8'h10 ;
			data[44662] <= 8'h10 ;
			data[44663] <= 8'h10 ;
			data[44664] <= 8'h10 ;
			data[44665] <= 8'h10 ;
			data[44666] <= 8'h10 ;
			data[44667] <= 8'h10 ;
			data[44668] <= 8'h10 ;
			data[44669] <= 8'h10 ;
			data[44670] <= 8'h10 ;
			data[44671] <= 8'h10 ;
			data[44672] <= 8'h10 ;
			data[44673] <= 8'h10 ;
			data[44674] <= 8'h10 ;
			data[44675] <= 8'h10 ;
			data[44676] <= 8'h10 ;
			data[44677] <= 8'h10 ;
			data[44678] <= 8'h10 ;
			data[44679] <= 8'h10 ;
			data[44680] <= 8'h10 ;
			data[44681] <= 8'h10 ;
			data[44682] <= 8'h10 ;
			data[44683] <= 8'h10 ;
			data[44684] <= 8'h10 ;
			data[44685] <= 8'h10 ;
			data[44686] <= 8'h10 ;
			data[44687] <= 8'h10 ;
			data[44688] <= 8'h10 ;
			data[44689] <= 8'h10 ;
			data[44690] <= 8'h10 ;
			data[44691] <= 8'h10 ;
			data[44692] <= 8'h10 ;
			data[44693] <= 8'h10 ;
			data[44694] <= 8'h10 ;
			data[44695] <= 8'h10 ;
			data[44696] <= 8'h10 ;
			data[44697] <= 8'h10 ;
			data[44698] <= 8'h10 ;
			data[44699] <= 8'h10 ;
			data[44700] <= 8'h10 ;
			data[44701] <= 8'h10 ;
			data[44702] <= 8'h10 ;
			data[44703] <= 8'h10 ;
			data[44704] <= 8'h10 ;
			data[44705] <= 8'h10 ;
			data[44706] <= 8'h10 ;
			data[44707] <= 8'h10 ;
			data[44708] <= 8'h10 ;
			data[44709] <= 8'h10 ;
			data[44710] <= 8'h10 ;
			data[44711] <= 8'h10 ;
			data[44712] <= 8'h10 ;
			data[44713] <= 8'h10 ;
			data[44714] <= 8'h10 ;
			data[44715] <= 8'h10 ;
			data[44716] <= 8'h10 ;
			data[44717] <= 8'h10 ;
			data[44718] <= 8'h10 ;
			data[44719] <= 8'h10 ;
			data[44720] <= 8'h10 ;
			data[44721] <= 8'h10 ;
			data[44722] <= 8'h10 ;
			data[44723] <= 8'h10 ;
			data[44724] <= 8'h10 ;
			data[44725] <= 8'h10 ;
			data[44726] <= 8'h10 ;
			data[44727] <= 8'h10 ;
			data[44728] <= 8'h10 ;
			data[44729] <= 8'h10 ;
			data[44730] <= 8'h10 ;
			data[44731] <= 8'h10 ;
			data[44732] <= 8'h10 ;
			data[44733] <= 8'h10 ;
			data[44734] <= 8'h10 ;
			data[44735] <= 8'h10 ;
			data[44736] <= 8'h10 ;
			data[44737] <= 8'h10 ;
			data[44738] <= 8'h10 ;
			data[44739] <= 8'h10 ;
			data[44740] <= 8'h10 ;
			data[44741] <= 8'h10 ;
			data[44742] <= 8'h10 ;
			data[44743] <= 8'h10 ;
			data[44744] <= 8'h10 ;
			data[44745] <= 8'h10 ;
			data[44746] <= 8'h10 ;
			data[44747] <= 8'h10 ;
			data[44748] <= 8'h10 ;
			data[44749] <= 8'h10 ;
			data[44750] <= 8'h10 ;
			data[44751] <= 8'h10 ;
			data[44752] <= 8'h10 ;
			data[44753] <= 8'h10 ;
			data[44754] <= 8'h10 ;
			data[44755] <= 8'h10 ;
			data[44756] <= 8'h10 ;
			data[44757] <= 8'h10 ;
			data[44758] <= 8'h10 ;
			data[44759] <= 8'h10 ;
			data[44760] <= 8'h10 ;
			data[44761] <= 8'h10 ;
			data[44762] <= 8'h10 ;
			data[44763] <= 8'h10 ;
			data[44764] <= 8'h10 ;
			data[44765] <= 8'h10 ;
			data[44766] <= 8'h10 ;
			data[44767] <= 8'h10 ;
			data[44768] <= 8'h10 ;
			data[44769] <= 8'h10 ;
			data[44770] <= 8'h10 ;
			data[44771] <= 8'h10 ;
			data[44772] <= 8'h10 ;
			data[44773] <= 8'h10 ;
			data[44774] <= 8'h10 ;
			data[44775] <= 8'h10 ;
			data[44776] <= 8'h10 ;
			data[44777] <= 8'h10 ;
			data[44778] <= 8'h10 ;
			data[44779] <= 8'h10 ;
			data[44780] <= 8'h10 ;
			data[44781] <= 8'h10 ;
			data[44782] <= 8'h10 ;
			data[44783] <= 8'h10 ;
			data[44784] <= 8'h10 ;
			data[44785] <= 8'h10 ;
			data[44786] <= 8'h10 ;
			data[44787] <= 8'h10 ;
			data[44788] <= 8'h10 ;
			data[44789] <= 8'h10 ;
			data[44790] <= 8'h10 ;
			data[44791] <= 8'h10 ;
			data[44792] <= 8'h10 ;
			data[44793] <= 8'h10 ;
			data[44794] <= 8'h10 ;
			data[44795] <= 8'h10 ;
			data[44796] <= 8'h10 ;
			data[44797] <= 8'h10 ;
			data[44798] <= 8'h10 ;
			data[44799] <= 8'h10 ;
			data[44800] <= 8'h10 ;
			data[44801] <= 8'h10 ;
			data[44802] <= 8'h10 ;
			data[44803] <= 8'h10 ;
			data[44804] <= 8'h10 ;
			data[44805] <= 8'h10 ;
			data[44806] <= 8'h10 ;
			data[44807] <= 8'h10 ;
			data[44808] <= 8'h10 ;
			data[44809] <= 8'h10 ;
			data[44810] <= 8'h10 ;
			data[44811] <= 8'h10 ;
			data[44812] <= 8'h10 ;
			data[44813] <= 8'h10 ;
			data[44814] <= 8'h10 ;
			data[44815] <= 8'h10 ;
			data[44816] <= 8'h10 ;
			data[44817] <= 8'h10 ;
			data[44818] <= 8'h10 ;
			data[44819] <= 8'h10 ;
			data[44820] <= 8'h10 ;
			data[44821] <= 8'h10 ;
			data[44822] <= 8'h10 ;
			data[44823] <= 8'h10 ;
			data[44824] <= 8'h10 ;
			data[44825] <= 8'h10 ;
			data[44826] <= 8'h10 ;
			data[44827] <= 8'h10 ;
			data[44828] <= 8'h10 ;
			data[44829] <= 8'h10 ;
			data[44830] <= 8'h10 ;
			data[44831] <= 8'h10 ;
			data[44832] <= 8'h10 ;
			data[44833] <= 8'h10 ;
			data[44834] <= 8'h10 ;
			data[44835] <= 8'h10 ;
			data[44836] <= 8'h10 ;
			data[44837] <= 8'h10 ;
			data[44838] <= 8'h10 ;
			data[44839] <= 8'h10 ;
			data[44840] <= 8'h10 ;
			data[44841] <= 8'h10 ;
			data[44842] <= 8'h10 ;
			data[44843] <= 8'h10 ;
			data[44844] <= 8'h10 ;
			data[44845] <= 8'h10 ;
			data[44846] <= 8'h10 ;
			data[44847] <= 8'h10 ;
			data[44848] <= 8'h10 ;
			data[44849] <= 8'h10 ;
			data[44850] <= 8'h10 ;
			data[44851] <= 8'h10 ;
			data[44852] <= 8'h10 ;
			data[44853] <= 8'h10 ;
			data[44854] <= 8'h10 ;
			data[44855] <= 8'h10 ;
			data[44856] <= 8'h10 ;
			data[44857] <= 8'h10 ;
			data[44858] <= 8'h10 ;
			data[44859] <= 8'h10 ;
			data[44860] <= 8'h10 ;
			data[44861] <= 8'h10 ;
			data[44862] <= 8'h10 ;
			data[44863] <= 8'h10 ;
			data[44864] <= 8'h10 ;
			data[44865] <= 8'h10 ;
			data[44866] <= 8'h10 ;
			data[44867] <= 8'h10 ;
			data[44868] <= 8'h10 ;
			data[44869] <= 8'h10 ;
			data[44870] <= 8'h10 ;
			data[44871] <= 8'h10 ;
			data[44872] <= 8'h10 ;
			data[44873] <= 8'h10 ;
			data[44874] <= 8'h10 ;
			data[44875] <= 8'h10 ;
			data[44876] <= 8'h10 ;
			data[44877] <= 8'h10 ;
			data[44878] <= 8'h10 ;
			data[44879] <= 8'h10 ;
			data[44880] <= 8'h10 ;
			data[44881] <= 8'h10 ;
			data[44882] <= 8'h10 ;
			data[44883] <= 8'h10 ;
			data[44884] <= 8'h10 ;
			data[44885] <= 8'h10 ;
			data[44886] <= 8'h10 ;
			data[44887] <= 8'h10 ;
			data[44888] <= 8'h10 ;
			data[44889] <= 8'h10 ;
			data[44890] <= 8'h10 ;
			data[44891] <= 8'h10 ;
			data[44892] <= 8'h10 ;
			data[44893] <= 8'h10 ;
			data[44894] <= 8'h10 ;
			data[44895] <= 8'h10 ;
			data[44896] <= 8'h10 ;
			data[44897] <= 8'h10 ;
			data[44898] <= 8'h10 ;
			data[44899] <= 8'h10 ;
			data[44900] <= 8'h10 ;
			data[44901] <= 8'h10 ;
			data[44902] <= 8'h10 ;
			data[44903] <= 8'h10 ;
			data[44904] <= 8'h10 ;
			data[44905] <= 8'h10 ;
			data[44906] <= 8'h10 ;
			data[44907] <= 8'h10 ;
			data[44908] <= 8'h10 ;
			data[44909] <= 8'h10 ;
			data[44910] <= 8'h10 ;
			data[44911] <= 8'h10 ;
			data[44912] <= 8'h10 ;
			data[44913] <= 8'h10 ;
			data[44914] <= 8'h10 ;
			data[44915] <= 8'h10 ;
			data[44916] <= 8'h10 ;
			data[44917] <= 8'h10 ;
			data[44918] <= 8'h10 ;
			data[44919] <= 8'h10 ;
			data[44920] <= 8'h10 ;
			data[44921] <= 8'h10 ;
			data[44922] <= 8'h10 ;
			data[44923] <= 8'h10 ;
			data[44924] <= 8'h10 ;
			data[44925] <= 8'h10 ;
			data[44926] <= 8'h10 ;
			data[44927] <= 8'h10 ;
			data[44928] <= 8'h10 ;
			data[44929] <= 8'h10 ;
			data[44930] <= 8'h10 ;
			data[44931] <= 8'h10 ;
			data[44932] <= 8'h10 ;
			data[44933] <= 8'h10 ;
			data[44934] <= 8'h10 ;
			data[44935] <= 8'h10 ;
			data[44936] <= 8'h10 ;
			data[44937] <= 8'h10 ;
			data[44938] <= 8'h10 ;
			data[44939] <= 8'h10 ;
			data[44940] <= 8'h10 ;
			data[44941] <= 8'h10 ;
			data[44942] <= 8'h10 ;
			data[44943] <= 8'h10 ;
			data[44944] <= 8'h10 ;
			data[44945] <= 8'h10 ;
			data[44946] <= 8'h10 ;
			data[44947] <= 8'h10 ;
			data[44948] <= 8'h10 ;
			data[44949] <= 8'h10 ;
			data[44950] <= 8'h10 ;
			data[44951] <= 8'h10 ;
			data[44952] <= 8'h10 ;
			data[44953] <= 8'h10 ;
			data[44954] <= 8'h10 ;
			data[44955] <= 8'h10 ;
			data[44956] <= 8'h10 ;
			data[44957] <= 8'h10 ;
			data[44958] <= 8'h10 ;
			data[44959] <= 8'h10 ;
			data[44960] <= 8'h10 ;
			data[44961] <= 8'h10 ;
			data[44962] <= 8'h10 ;
			data[44963] <= 8'h10 ;
			data[44964] <= 8'h10 ;
			data[44965] <= 8'h10 ;
			data[44966] <= 8'h10 ;
			data[44967] <= 8'h10 ;
			data[44968] <= 8'h10 ;
			data[44969] <= 8'h10 ;
			data[44970] <= 8'h10 ;
			data[44971] <= 8'h10 ;
			data[44972] <= 8'h10 ;
			data[44973] <= 8'h10 ;
			data[44974] <= 8'h10 ;
			data[44975] <= 8'h10 ;
			data[44976] <= 8'h10 ;
			data[44977] <= 8'h10 ;
			data[44978] <= 8'h10 ;
			data[44979] <= 8'h10 ;
			data[44980] <= 8'h10 ;
			data[44981] <= 8'h10 ;
			data[44982] <= 8'h10 ;
			data[44983] <= 8'h10 ;
			data[44984] <= 8'h10 ;
			data[44985] <= 8'h10 ;
			data[44986] <= 8'h10 ;
			data[44987] <= 8'h10 ;
			data[44988] <= 8'h10 ;
			data[44989] <= 8'h10 ;
			data[44990] <= 8'h10 ;
			data[44991] <= 8'h10 ;
			data[44992] <= 8'h10 ;
			data[44993] <= 8'h10 ;
			data[44994] <= 8'h10 ;
			data[44995] <= 8'h10 ;
			data[44996] <= 8'h10 ;
			data[44997] <= 8'h10 ;
			data[44998] <= 8'h10 ;
			data[44999] <= 8'h10 ;
			data[45000] <= 8'h10 ;
			data[45001] <= 8'h10 ;
			data[45002] <= 8'h10 ;
			data[45003] <= 8'h10 ;
			data[45004] <= 8'h10 ;
			data[45005] <= 8'h10 ;
			data[45006] <= 8'h10 ;
			data[45007] <= 8'h10 ;
			data[45008] <= 8'h10 ;
			data[45009] <= 8'h10 ;
			data[45010] <= 8'h10 ;
			data[45011] <= 8'h10 ;
			data[45012] <= 8'h10 ;
			data[45013] <= 8'h10 ;
			data[45014] <= 8'h10 ;
			data[45015] <= 8'h10 ;
			data[45016] <= 8'h10 ;
			data[45017] <= 8'h10 ;
			data[45018] <= 8'h10 ;
			data[45019] <= 8'h10 ;
			data[45020] <= 8'h10 ;
			data[45021] <= 8'h10 ;
			data[45022] <= 8'h10 ;
			data[45023] <= 8'h10 ;
			data[45024] <= 8'h10 ;
			data[45025] <= 8'h10 ;
			data[45026] <= 8'h10 ;
			data[45027] <= 8'h10 ;
			data[45028] <= 8'h10 ;
			data[45029] <= 8'h10 ;
			data[45030] <= 8'h10 ;
			data[45031] <= 8'h10 ;
			data[45032] <= 8'h10 ;
			data[45033] <= 8'h10 ;
			data[45034] <= 8'h10 ;
			data[45035] <= 8'h10 ;
			data[45036] <= 8'h10 ;
			data[45037] <= 8'h10 ;
			data[45038] <= 8'h10 ;
			data[45039] <= 8'h10 ;
			data[45040] <= 8'h10 ;
			data[45041] <= 8'h10 ;
			data[45042] <= 8'h10 ;
			data[45043] <= 8'h10 ;
			data[45044] <= 8'h10 ;
			data[45045] <= 8'h10 ;
			data[45046] <= 8'h10 ;
			data[45047] <= 8'h10 ;
			data[45048] <= 8'h10 ;
			data[45049] <= 8'h10 ;
			data[45050] <= 8'h10 ;
			data[45051] <= 8'h10 ;
			data[45052] <= 8'h10 ;
			data[45053] <= 8'h10 ;
			data[45054] <= 8'h10 ;
			data[45055] <= 8'h10 ;
			data[45056] <= 8'h10 ;
			data[45057] <= 8'h10 ;
			data[45058] <= 8'h10 ;
			data[45059] <= 8'h10 ;
			data[45060] <= 8'h10 ;
			data[45061] <= 8'h10 ;
			data[45062] <= 8'h10 ;
			data[45063] <= 8'h10 ;
			data[45064] <= 8'h10 ;
			data[45065] <= 8'h10 ;
			data[45066] <= 8'h10 ;
			data[45067] <= 8'h10 ;
			data[45068] <= 8'h10 ;
			data[45069] <= 8'h10 ;
			data[45070] <= 8'h10 ;
			data[45071] <= 8'h10 ;
			data[45072] <= 8'h10 ;
			data[45073] <= 8'h10 ;
			data[45074] <= 8'h10 ;
			data[45075] <= 8'h10 ;
			data[45076] <= 8'h10 ;
			data[45077] <= 8'h10 ;
			data[45078] <= 8'h10 ;
			data[45079] <= 8'h10 ;
			data[45080] <= 8'h10 ;
			data[45081] <= 8'h10 ;
			data[45082] <= 8'h10 ;
			data[45083] <= 8'h10 ;
			data[45084] <= 8'h10 ;
			data[45085] <= 8'h10 ;
			data[45086] <= 8'h10 ;
			data[45087] <= 8'h10 ;
			data[45088] <= 8'h10 ;
			data[45089] <= 8'h10 ;
			data[45090] <= 8'h10 ;
			data[45091] <= 8'h10 ;
			data[45092] <= 8'h10 ;
			data[45093] <= 8'h10 ;
			data[45094] <= 8'h10 ;
			data[45095] <= 8'h10 ;
			data[45096] <= 8'h10 ;
			data[45097] <= 8'h10 ;
			data[45098] <= 8'h10 ;
			data[45099] <= 8'h10 ;
			data[45100] <= 8'h10 ;
			data[45101] <= 8'h10 ;
			data[45102] <= 8'h10 ;
			data[45103] <= 8'h10 ;
			data[45104] <= 8'h10 ;
			data[45105] <= 8'h10 ;
			data[45106] <= 8'h10 ;
			data[45107] <= 8'h10 ;
			data[45108] <= 8'h10 ;
			data[45109] <= 8'h10 ;
			data[45110] <= 8'h10 ;
			data[45111] <= 8'h10 ;
			data[45112] <= 8'h10 ;
			data[45113] <= 8'h10 ;
			data[45114] <= 8'h10 ;
			data[45115] <= 8'h10 ;
			data[45116] <= 8'h10 ;
			data[45117] <= 8'h10 ;
			data[45118] <= 8'h10 ;
			data[45119] <= 8'h10 ;
			data[45120] <= 8'h10 ;
			data[45121] <= 8'h10 ;
			data[45122] <= 8'h10 ;
			data[45123] <= 8'h10 ;
			data[45124] <= 8'h10 ;
			data[45125] <= 8'h10 ;
			data[45126] <= 8'h10 ;
			data[45127] <= 8'h10 ;
			data[45128] <= 8'h10 ;
			data[45129] <= 8'h10 ;
			data[45130] <= 8'h10 ;
			data[45131] <= 8'h10 ;
			data[45132] <= 8'h10 ;
			data[45133] <= 8'h10 ;
			data[45134] <= 8'h10 ;
			data[45135] <= 8'h10 ;
			data[45136] <= 8'h10 ;
			data[45137] <= 8'h10 ;
			data[45138] <= 8'h10 ;
			data[45139] <= 8'h10 ;
			data[45140] <= 8'h10 ;
			data[45141] <= 8'h10 ;
			data[45142] <= 8'h10 ;
			data[45143] <= 8'h10 ;
			data[45144] <= 8'h10 ;
			data[45145] <= 8'h10 ;
			data[45146] <= 8'h10 ;
			data[45147] <= 8'h10 ;
			data[45148] <= 8'h10 ;
			data[45149] <= 8'h10 ;
			data[45150] <= 8'h10 ;
			data[45151] <= 8'h10 ;
			data[45152] <= 8'h10 ;
			data[45153] <= 8'h10 ;
			data[45154] <= 8'h10 ;
			data[45155] <= 8'h10 ;
			data[45156] <= 8'h10 ;
			data[45157] <= 8'h10 ;
			data[45158] <= 8'h10 ;
			data[45159] <= 8'h10 ;
			data[45160] <= 8'h10 ;
			data[45161] <= 8'h10 ;
			data[45162] <= 8'h10 ;
			data[45163] <= 8'h10 ;
			data[45164] <= 8'h10 ;
			data[45165] <= 8'h10 ;
			data[45166] <= 8'h10 ;
			data[45167] <= 8'h10 ;
			data[45168] <= 8'h10 ;
			data[45169] <= 8'h10 ;
			data[45170] <= 8'h10 ;
			data[45171] <= 8'h10 ;
			data[45172] <= 8'h10 ;
			data[45173] <= 8'h10 ;
			data[45174] <= 8'h10 ;
			data[45175] <= 8'h10 ;
			data[45176] <= 8'h10 ;
			data[45177] <= 8'h10 ;
			data[45178] <= 8'h10 ;
			data[45179] <= 8'h10 ;
			data[45180] <= 8'h10 ;
			data[45181] <= 8'h10 ;
			data[45182] <= 8'h10 ;
			data[45183] <= 8'h10 ;
			data[45184] <= 8'h10 ;
			data[45185] <= 8'h10 ;
			data[45186] <= 8'h10 ;
			data[45187] <= 8'h10 ;
			data[45188] <= 8'h10 ;
			data[45189] <= 8'h10 ;
			data[45190] <= 8'h10 ;
			data[45191] <= 8'h10 ;
			data[45192] <= 8'h10 ;
			data[45193] <= 8'h10 ;
			data[45194] <= 8'h10 ;
			data[45195] <= 8'h10 ;
			data[45196] <= 8'h10 ;
			data[45197] <= 8'h10 ;
			data[45198] <= 8'h10 ;
			data[45199] <= 8'h10 ;
			data[45200] <= 8'h10 ;
			data[45201] <= 8'h10 ;
			data[45202] <= 8'h10 ;
			data[45203] <= 8'h10 ;
			data[45204] <= 8'h10 ;
			data[45205] <= 8'h10 ;
			data[45206] <= 8'h10 ;
			data[45207] <= 8'h10 ;
			data[45208] <= 8'h10 ;
			data[45209] <= 8'h10 ;
			data[45210] <= 8'h10 ;
			data[45211] <= 8'h10 ;
			data[45212] <= 8'h10 ;
			data[45213] <= 8'h10 ;
			data[45214] <= 8'h10 ;
			data[45215] <= 8'h10 ;
			data[45216] <= 8'h10 ;
			data[45217] <= 8'h10 ;
			data[45218] <= 8'h10 ;
			data[45219] <= 8'h10 ;
			data[45220] <= 8'h10 ;
			data[45221] <= 8'h10 ;
			data[45222] <= 8'h10 ;
			data[45223] <= 8'h10 ;
			data[45224] <= 8'h10 ;
			data[45225] <= 8'h10 ;
			data[45226] <= 8'h10 ;
			data[45227] <= 8'h10 ;
			data[45228] <= 8'h10 ;
			data[45229] <= 8'h10 ;
			data[45230] <= 8'h10 ;
			data[45231] <= 8'h10 ;
			data[45232] <= 8'h10 ;
			data[45233] <= 8'h10 ;
			data[45234] <= 8'h10 ;
			data[45235] <= 8'h10 ;
			data[45236] <= 8'h10 ;
			data[45237] <= 8'h10 ;
			data[45238] <= 8'h10 ;
			data[45239] <= 8'h10 ;
			data[45240] <= 8'h10 ;
			data[45241] <= 8'h10 ;
			data[45242] <= 8'h10 ;
			data[45243] <= 8'h10 ;
			data[45244] <= 8'h10 ;
			data[45245] <= 8'h10 ;
			data[45246] <= 8'h10 ;
			data[45247] <= 8'h10 ;
			data[45248] <= 8'h10 ;
			data[45249] <= 8'h10 ;
			data[45250] <= 8'h10 ;
			data[45251] <= 8'h10 ;
			data[45252] <= 8'h10 ;
			data[45253] <= 8'h10 ;
			data[45254] <= 8'h10 ;
			data[45255] <= 8'h10 ;
			data[45256] <= 8'h10 ;
			data[45257] <= 8'h10 ;
			data[45258] <= 8'h10 ;
			data[45259] <= 8'h10 ;
			data[45260] <= 8'h10 ;
			data[45261] <= 8'h10 ;
			data[45262] <= 8'h10 ;
			data[45263] <= 8'h10 ;
			data[45264] <= 8'h10 ;
			data[45265] <= 8'h10 ;
			data[45266] <= 8'h10 ;
			data[45267] <= 8'h10 ;
			data[45268] <= 8'h10 ;
			data[45269] <= 8'h10 ;
			data[45270] <= 8'h10 ;
			data[45271] <= 8'h10 ;
			data[45272] <= 8'h10 ;
			data[45273] <= 8'h10 ;
			data[45274] <= 8'h10 ;
			data[45275] <= 8'h10 ;
			data[45276] <= 8'h10 ;
			data[45277] <= 8'h10 ;
			data[45278] <= 8'h10 ;
			data[45279] <= 8'h10 ;
			data[45280] <= 8'h10 ;
			data[45281] <= 8'h10 ;
			data[45282] <= 8'h10 ;
			data[45283] <= 8'h10 ;
			data[45284] <= 8'h10 ;
			data[45285] <= 8'h10 ;
			data[45286] <= 8'h10 ;
			data[45287] <= 8'h10 ;
			data[45288] <= 8'h10 ;
			data[45289] <= 8'h10 ;
			data[45290] <= 8'h10 ;
			data[45291] <= 8'h10 ;
			data[45292] <= 8'h10 ;
			data[45293] <= 8'h10 ;
			data[45294] <= 8'h10 ;
			data[45295] <= 8'h10 ;
			data[45296] <= 8'h10 ;
			data[45297] <= 8'h10 ;
			data[45298] <= 8'h10 ;
			data[45299] <= 8'h10 ;
			data[45300] <= 8'h10 ;
			data[45301] <= 8'h10 ;
			data[45302] <= 8'h10 ;
			data[45303] <= 8'h10 ;
			data[45304] <= 8'h10 ;
			data[45305] <= 8'h10 ;
			data[45306] <= 8'h10 ;
			data[45307] <= 8'h10 ;
			data[45308] <= 8'h10 ;
			data[45309] <= 8'h10 ;
			data[45310] <= 8'h10 ;
			data[45311] <= 8'h10 ;
			data[45312] <= 8'h10 ;
			data[45313] <= 8'h10 ;
			data[45314] <= 8'h10 ;
			data[45315] <= 8'h10 ;
			data[45316] <= 8'h10 ;
			data[45317] <= 8'h10 ;
			data[45318] <= 8'h10 ;
			data[45319] <= 8'h10 ;
			data[45320] <= 8'h10 ;
			data[45321] <= 8'h10 ;
			data[45322] <= 8'h10 ;
			data[45323] <= 8'h10 ;
			data[45324] <= 8'h10 ;
			data[45325] <= 8'h10 ;
			data[45326] <= 8'h10 ;
			data[45327] <= 8'h10 ;
			data[45328] <= 8'h10 ;
			data[45329] <= 8'h10 ;
			data[45330] <= 8'h10 ;
			data[45331] <= 8'h10 ;
			data[45332] <= 8'h10 ;
			data[45333] <= 8'h10 ;
			data[45334] <= 8'h10 ;
			data[45335] <= 8'h10 ;
			data[45336] <= 8'h10 ;
			data[45337] <= 8'h10 ;
			data[45338] <= 8'h10 ;
			data[45339] <= 8'h10 ;
			data[45340] <= 8'h10 ;
			data[45341] <= 8'h10 ;
			data[45342] <= 8'h10 ;
			data[45343] <= 8'h10 ;
			data[45344] <= 8'h10 ;
			data[45345] <= 8'h10 ;
			data[45346] <= 8'h10 ;
			data[45347] <= 8'h10 ;
			data[45348] <= 8'h10 ;
			data[45349] <= 8'h10 ;
			data[45350] <= 8'h10 ;
			data[45351] <= 8'h10 ;
			data[45352] <= 8'h10 ;
			data[45353] <= 8'h10 ;
			data[45354] <= 8'h10 ;
			data[45355] <= 8'h10 ;
			data[45356] <= 8'h10 ;
			data[45357] <= 8'h10 ;
			data[45358] <= 8'h10 ;
			data[45359] <= 8'h10 ;
			data[45360] <= 8'h10 ;
			data[45361] <= 8'h10 ;
			data[45362] <= 8'h10 ;
			data[45363] <= 8'h10 ;
			data[45364] <= 8'h10 ;
			data[45365] <= 8'h10 ;
			data[45366] <= 8'h10 ;
			data[45367] <= 8'h10 ;
			data[45368] <= 8'h10 ;
			data[45369] <= 8'h10 ;
			data[45370] <= 8'h10 ;
			data[45371] <= 8'h10 ;
			data[45372] <= 8'h10 ;
			data[45373] <= 8'h10 ;
			data[45374] <= 8'h10 ;
			data[45375] <= 8'h10 ;
			data[45376] <= 8'h10 ;
			data[45377] <= 8'h10 ;
			data[45378] <= 8'h10 ;
			data[45379] <= 8'h10 ;
			data[45380] <= 8'h10 ;
			data[45381] <= 8'h10 ;
			data[45382] <= 8'h10 ;
			data[45383] <= 8'h10 ;
			data[45384] <= 8'h10 ;
			data[45385] <= 8'h10 ;
			data[45386] <= 8'h10 ;
			data[45387] <= 8'h10 ;
			data[45388] <= 8'h10 ;
			data[45389] <= 8'h10 ;
			data[45390] <= 8'h10 ;
			data[45391] <= 8'h10 ;
			data[45392] <= 8'h10 ;
			data[45393] <= 8'h10 ;
			data[45394] <= 8'h10 ;
			data[45395] <= 8'h10 ;
			data[45396] <= 8'h10 ;
			data[45397] <= 8'h10 ;
			data[45398] <= 8'h10 ;
			data[45399] <= 8'h10 ;
			data[45400] <= 8'h10 ;
			data[45401] <= 8'h10 ;
			data[45402] <= 8'h10 ;
			data[45403] <= 8'h10 ;
			data[45404] <= 8'h10 ;
			data[45405] <= 8'h10 ;
			data[45406] <= 8'h10 ;
			data[45407] <= 8'h10 ;
			data[45408] <= 8'h10 ;
			data[45409] <= 8'h10 ;
			data[45410] <= 8'h10 ;
			data[45411] <= 8'h10 ;
			data[45412] <= 8'h10 ;
			data[45413] <= 8'h10 ;
			data[45414] <= 8'h10 ;
			data[45415] <= 8'h10 ;
			data[45416] <= 8'h10 ;
			data[45417] <= 8'h10 ;
			data[45418] <= 8'h10 ;
			data[45419] <= 8'h10 ;
			data[45420] <= 8'h10 ;
			data[45421] <= 8'h10 ;
			data[45422] <= 8'h10 ;
			data[45423] <= 8'h10 ;
			data[45424] <= 8'h10 ;
			data[45425] <= 8'h10 ;
			data[45426] <= 8'h10 ;
			data[45427] <= 8'h10 ;
			data[45428] <= 8'h10 ;
			data[45429] <= 8'h10 ;
			data[45430] <= 8'h10 ;
			data[45431] <= 8'h10 ;
			data[45432] <= 8'h10 ;
			data[45433] <= 8'h10 ;
			data[45434] <= 8'h10 ;
			data[45435] <= 8'h10 ;
			data[45436] <= 8'h10 ;
			data[45437] <= 8'h10 ;
			data[45438] <= 8'h10 ;
			data[45439] <= 8'h10 ;
			data[45440] <= 8'h10 ;
			data[45441] <= 8'h10 ;
			data[45442] <= 8'h10 ;
			data[45443] <= 8'h10 ;
			data[45444] <= 8'h10 ;
			data[45445] <= 8'h10 ;
			data[45446] <= 8'h10 ;
			data[45447] <= 8'h10 ;
			data[45448] <= 8'h10 ;
			data[45449] <= 8'h10 ;
			data[45450] <= 8'h10 ;
			data[45451] <= 8'h10 ;
			data[45452] <= 8'h10 ;
			data[45453] <= 8'h10 ;
			data[45454] <= 8'h10 ;
			data[45455] <= 8'h10 ;
			data[45456] <= 8'h10 ;
			data[45457] <= 8'h10 ;
			data[45458] <= 8'h10 ;
			data[45459] <= 8'h10 ;
			data[45460] <= 8'h10 ;
			data[45461] <= 8'h10 ;
			data[45462] <= 8'h10 ;
			data[45463] <= 8'h10 ;
			data[45464] <= 8'h10 ;
			data[45465] <= 8'h10 ;
			data[45466] <= 8'h10 ;
			data[45467] <= 8'h10 ;
			data[45468] <= 8'h10 ;
			data[45469] <= 8'h10 ;
			data[45470] <= 8'h10 ;
			data[45471] <= 8'h10 ;
			data[45472] <= 8'h10 ;
			data[45473] <= 8'h10 ;
			data[45474] <= 8'h10 ;
			data[45475] <= 8'h10 ;
			data[45476] <= 8'h10 ;
			data[45477] <= 8'h10 ;
			data[45478] <= 8'h10 ;
			data[45479] <= 8'h10 ;
			data[45480] <= 8'h10 ;
			data[45481] <= 8'h10 ;
			data[45482] <= 8'h10 ;
			data[45483] <= 8'h10 ;
			data[45484] <= 8'h10 ;
			data[45485] <= 8'h10 ;
			data[45486] <= 8'h10 ;
			data[45487] <= 8'h10 ;
			data[45488] <= 8'h10 ;
			data[45489] <= 8'h10 ;
			data[45490] <= 8'h10 ;
			data[45491] <= 8'h10 ;
			data[45492] <= 8'h10 ;
			data[45493] <= 8'h10 ;
			data[45494] <= 8'h10 ;
			data[45495] <= 8'h10 ;
			data[45496] <= 8'h10 ;
			data[45497] <= 8'h10 ;
			data[45498] <= 8'h10 ;
			data[45499] <= 8'h10 ;
			data[45500] <= 8'h10 ;
			data[45501] <= 8'h10 ;
			data[45502] <= 8'h10 ;
			data[45503] <= 8'h10 ;
			data[45504] <= 8'h10 ;
			data[45505] <= 8'h10 ;
			data[45506] <= 8'h10 ;
			data[45507] <= 8'h10 ;
			data[45508] <= 8'h10 ;
			data[45509] <= 8'h10 ;
			data[45510] <= 8'h10 ;
			data[45511] <= 8'h10 ;
			data[45512] <= 8'h10 ;
			data[45513] <= 8'h10 ;
			data[45514] <= 8'h10 ;
			data[45515] <= 8'h10 ;
			data[45516] <= 8'h10 ;
			data[45517] <= 8'h10 ;
			data[45518] <= 8'h10 ;
			data[45519] <= 8'h10 ;
			data[45520] <= 8'h10 ;
			data[45521] <= 8'h10 ;
			data[45522] <= 8'h10 ;
			data[45523] <= 8'h10 ;
			data[45524] <= 8'h10 ;
			data[45525] <= 8'h10 ;
			data[45526] <= 8'h10 ;
			data[45527] <= 8'h10 ;
			data[45528] <= 8'h10 ;
			data[45529] <= 8'h10 ;
			data[45530] <= 8'h10 ;
			data[45531] <= 8'h10 ;
			data[45532] <= 8'h10 ;
			data[45533] <= 8'h10 ;
			data[45534] <= 8'h10 ;
			data[45535] <= 8'h10 ;
			data[45536] <= 8'h10 ;
			data[45537] <= 8'h10 ;
			data[45538] <= 8'h10 ;
			data[45539] <= 8'h10 ;
			data[45540] <= 8'h10 ;
			data[45541] <= 8'h10 ;
			data[45542] <= 8'h10 ;
			data[45543] <= 8'h10 ;
			data[45544] <= 8'h10 ;
			data[45545] <= 8'h10 ;
			data[45546] <= 8'h10 ;
			data[45547] <= 8'h10 ;
			data[45548] <= 8'h10 ;
			data[45549] <= 8'h10 ;
			data[45550] <= 8'h10 ;
			data[45551] <= 8'h10 ;
			data[45552] <= 8'h10 ;
			data[45553] <= 8'h10 ;
			data[45554] <= 8'h10 ;
			data[45555] <= 8'h10 ;
			data[45556] <= 8'h10 ;
			data[45557] <= 8'h10 ;
			data[45558] <= 8'h10 ;
			data[45559] <= 8'h10 ;
			data[45560] <= 8'h10 ;
			data[45561] <= 8'h10 ;
			data[45562] <= 8'h10 ;
			data[45563] <= 8'h10 ;
			data[45564] <= 8'h10 ;
			data[45565] <= 8'h10 ;
			data[45566] <= 8'h10 ;
			data[45567] <= 8'h10 ;
			data[45568] <= 8'h10 ;
			data[45569] <= 8'h10 ;
			data[45570] <= 8'h10 ;
			data[45571] <= 8'h10 ;
			data[45572] <= 8'h10 ;
			data[45573] <= 8'h10 ;
			data[45574] <= 8'h10 ;
			data[45575] <= 8'h10 ;
			data[45576] <= 8'h10 ;
			data[45577] <= 8'h10 ;
			data[45578] <= 8'h10 ;
			data[45579] <= 8'h10 ;
			data[45580] <= 8'h10 ;
			data[45581] <= 8'h10 ;
			data[45582] <= 8'h10 ;
			data[45583] <= 8'h10 ;
			data[45584] <= 8'h10 ;
			data[45585] <= 8'h10 ;
			data[45586] <= 8'h10 ;
			data[45587] <= 8'h10 ;
			data[45588] <= 8'h10 ;
			data[45589] <= 8'h10 ;
			data[45590] <= 8'h10 ;
			data[45591] <= 8'h10 ;
			data[45592] <= 8'h10 ;
			data[45593] <= 8'h10 ;
			data[45594] <= 8'h10 ;
			data[45595] <= 8'h10 ;
			data[45596] <= 8'h10 ;
			data[45597] <= 8'h10 ;
			data[45598] <= 8'h10 ;
			data[45599] <= 8'h10 ;
			data[45600] <= 8'h10 ;
			data[45601] <= 8'h10 ;
			data[45602] <= 8'h10 ;
			data[45603] <= 8'h10 ;
			data[45604] <= 8'h10 ;
			data[45605] <= 8'h10 ;
			data[45606] <= 8'h10 ;
			data[45607] <= 8'h10 ;
			data[45608] <= 8'h10 ;
			data[45609] <= 8'h10 ;
			data[45610] <= 8'h10 ;
			data[45611] <= 8'h10 ;
			data[45612] <= 8'h10 ;
			data[45613] <= 8'h10 ;
			data[45614] <= 8'h10 ;
			data[45615] <= 8'h10 ;
			data[45616] <= 8'h10 ;
			data[45617] <= 8'h10 ;
			data[45618] <= 8'h10 ;
			data[45619] <= 8'h10 ;
			data[45620] <= 8'h10 ;
			data[45621] <= 8'h10 ;
			data[45622] <= 8'h10 ;
			data[45623] <= 8'h10 ;
			data[45624] <= 8'h10 ;
			data[45625] <= 8'h10 ;
			data[45626] <= 8'h10 ;
			data[45627] <= 8'h10 ;
			data[45628] <= 8'h10 ;
			data[45629] <= 8'h10 ;
			data[45630] <= 8'h10 ;
			data[45631] <= 8'h10 ;
			data[45632] <= 8'h10 ;
			data[45633] <= 8'h10 ;
			data[45634] <= 8'h10 ;
			data[45635] <= 8'h10 ;
			data[45636] <= 8'h10 ;
			data[45637] <= 8'h10 ;
			data[45638] <= 8'h10 ;
			data[45639] <= 8'h10 ;
			data[45640] <= 8'h10 ;
			data[45641] <= 8'h10 ;
			data[45642] <= 8'h10 ;
			data[45643] <= 8'h10 ;
			data[45644] <= 8'h10 ;
			data[45645] <= 8'h10 ;
			data[45646] <= 8'h10 ;
			data[45647] <= 8'h10 ;
			data[45648] <= 8'h10 ;
			data[45649] <= 8'h10 ;
			data[45650] <= 8'h10 ;
			data[45651] <= 8'h10 ;
			data[45652] <= 8'h10 ;
			data[45653] <= 8'h10 ;
			data[45654] <= 8'h10 ;
			data[45655] <= 8'h10 ;
			data[45656] <= 8'h10 ;
			data[45657] <= 8'h10 ;
			data[45658] <= 8'h10 ;
			data[45659] <= 8'h10 ;
			data[45660] <= 8'h10 ;
			data[45661] <= 8'h10 ;
			data[45662] <= 8'h10 ;
			data[45663] <= 8'h10 ;
			data[45664] <= 8'h10 ;
			data[45665] <= 8'h10 ;
			data[45666] <= 8'h10 ;
			data[45667] <= 8'h10 ;
			data[45668] <= 8'h10 ;
			data[45669] <= 8'h10 ;
			data[45670] <= 8'h10 ;
			data[45671] <= 8'h10 ;
			data[45672] <= 8'h10 ;
			data[45673] <= 8'h10 ;
			data[45674] <= 8'h10 ;
			data[45675] <= 8'h10 ;
			data[45676] <= 8'h10 ;
			data[45677] <= 8'h10 ;
			data[45678] <= 8'h10 ;
			data[45679] <= 8'h10 ;
			data[45680] <= 8'h10 ;
			data[45681] <= 8'h10 ;
			data[45682] <= 8'h10 ;
			data[45683] <= 8'h10 ;
			data[45684] <= 8'h10 ;
			data[45685] <= 8'h10 ;
			data[45686] <= 8'h10 ;
			data[45687] <= 8'h10 ;
			data[45688] <= 8'h10 ;
			data[45689] <= 8'h10 ;
			data[45690] <= 8'h10 ;
			data[45691] <= 8'h10 ;
			data[45692] <= 8'h10 ;
			data[45693] <= 8'h10 ;
			data[45694] <= 8'h10 ;
			data[45695] <= 8'h10 ;
			data[45696] <= 8'h10 ;
			data[45697] <= 8'h10 ;
			data[45698] <= 8'h10 ;
			data[45699] <= 8'h10 ;
			data[45700] <= 8'h10 ;
			data[45701] <= 8'h10 ;
			data[45702] <= 8'h10 ;
			data[45703] <= 8'h10 ;
			data[45704] <= 8'h10 ;
			data[45705] <= 8'h10 ;
			data[45706] <= 8'h10 ;
			data[45707] <= 8'h10 ;
			data[45708] <= 8'h10 ;
			data[45709] <= 8'h10 ;
			data[45710] <= 8'h10 ;
			data[45711] <= 8'h10 ;
			data[45712] <= 8'h10 ;
			data[45713] <= 8'h10 ;
			data[45714] <= 8'h10 ;
			data[45715] <= 8'h10 ;
			data[45716] <= 8'h10 ;
			data[45717] <= 8'h10 ;
			data[45718] <= 8'h10 ;
			data[45719] <= 8'h10 ;
			data[45720] <= 8'h10 ;
			data[45721] <= 8'h10 ;
			data[45722] <= 8'h10 ;
			data[45723] <= 8'h10 ;
			data[45724] <= 8'h10 ;
			data[45725] <= 8'h10 ;
			data[45726] <= 8'h10 ;
			data[45727] <= 8'h10 ;
			data[45728] <= 8'h10 ;
			data[45729] <= 8'h10 ;
			data[45730] <= 8'h10 ;
			data[45731] <= 8'h10 ;
			data[45732] <= 8'h10 ;
			data[45733] <= 8'h10 ;
			data[45734] <= 8'h10 ;
			data[45735] <= 8'h10 ;
			data[45736] <= 8'h10 ;
			data[45737] <= 8'h10 ;
			data[45738] <= 8'h10 ;
			data[45739] <= 8'h10 ;
			data[45740] <= 8'h10 ;
			data[45741] <= 8'h10 ;
			data[45742] <= 8'h10 ;
			data[45743] <= 8'h10 ;
			data[45744] <= 8'h10 ;
			data[45745] <= 8'h10 ;
			data[45746] <= 8'h10 ;
			data[45747] <= 8'h10 ;
			data[45748] <= 8'h10 ;
			data[45749] <= 8'h10 ;
			data[45750] <= 8'h10 ;
			data[45751] <= 8'h10 ;
			data[45752] <= 8'h10 ;
			data[45753] <= 8'h10 ;
			data[45754] <= 8'h10 ;
			data[45755] <= 8'h10 ;
			data[45756] <= 8'h10 ;
			data[45757] <= 8'h10 ;
			data[45758] <= 8'h10 ;
			data[45759] <= 8'h10 ;
			data[45760] <= 8'h10 ;
			data[45761] <= 8'h10 ;
			data[45762] <= 8'h10 ;
			data[45763] <= 8'h10 ;
			data[45764] <= 8'h10 ;
			data[45765] <= 8'h10 ;
			data[45766] <= 8'h10 ;
			data[45767] <= 8'h10 ;
			data[45768] <= 8'h10 ;
			data[45769] <= 8'h10 ;
			data[45770] <= 8'h10 ;
			data[45771] <= 8'h10 ;
			data[45772] <= 8'h10 ;
			data[45773] <= 8'h10 ;
			data[45774] <= 8'h10 ;
			data[45775] <= 8'h10 ;
			data[45776] <= 8'h10 ;
			data[45777] <= 8'h10 ;
			data[45778] <= 8'h10 ;
			data[45779] <= 8'h10 ;
			data[45780] <= 8'h10 ;
			data[45781] <= 8'h10 ;
			data[45782] <= 8'h10 ;
			data[45783] <= 8'h10 ;
			data[45784] <= 8'h10 ;
			data[45785] <= 8'h10 ;
			data[45786] <= 8'h10 ;
			data[45787] <= 8'h10 ;
			data[45788] <= 8'h10 ;
			data[45789] <= 8'h10 ;
			data[45790] <= 8'h10 ;
			data[45791] <= 8'h10 ;
			data[45792] <= 8'h10 ;
			data[45793] <= 8'h10 ;
			data[45794] <= 8'h10 ;
			data[45795] <= 8'h10 ;
			data[45796] <= 8'h10 ;
			data[45797] <= 8'h10 ;
			data[45798] <= 8'h10 ;
			data[45799] <= 8'h10 ;
			data[45800] <= 8'h10 ;
			data[45801] <= 8'h10 ;
			data[45802] <= 8'h10 ;
			data[45803] <= 8'h10 ;
			data[45804] <= 8'h10 ;
			data[45805] <= 8'h10 ;
			data[45806] <= 8'h10 ;
			data[45807] <= 8'h10 ;
			data[45808] <= 8'h10 ;
			data[45809] <= 8'h10 ;
			data[45810] <= 8'h10 ;
			data[45811] <= 8'h10 ;
			data[45812] <= 8'h10 ;
			data[45813] <= 8'h10 ;
			data[45814] <= 8'h10 ;
			data[45815] <= 8'h10 ;
			data[45816] <= 8'h10 ;
			data[45817] <= 8'h10 ;
			data[45818] <= 8'h10 ;
			data[45819] <= 8'h10 ;
			data[45820] <= 8'h10 ;
			data[45821] <= 8'h10 ;
			data[45822] <= 8'h10 ;
			data[45823] <= 8'h10 ;
			data[45824] <= 8'h10 ;
			data[45825] <= 8'h10 ;
			data[45826] <= 8'h10 ;
			data[45827] <= 8'h10 ;
			data[45828] <= 8'h10 ;
			data[45829] <= 8'h10 ;
			data[45830] <= 8'h10 ;
			data[45831] <= 8'h10 ;
			data[45832] <= 8'h10 ;
			data[45833] <= 8'h10 ;
			data[45834] <= 8'h10 ;
			data[45835] <= 8'h10 ;
			data[45836] <= 8'h10 ;
			data[45837] <= 8'h10 ;
			data[45838] <= 8'h10 ;
			data[45839] <= 8'h10 ;
			data[45840] <= 8'h10 ;
			data[45841] <= 8'h10 ;
			data[45842] <= 8'h10 ;
			data[45843] <= 8'h10 ;
			data[45844] <= 8'h10 ;
			data[45845] <= 8'h10 ;
			data[45846] <= 8'h10 ;
			data[45847] <= 8'h10 ;
			data[45848] <= 8'h10 ;
			data[45849] <= 8'h10 ;
			data[45850] <= 8'h10 ;
			data[45851] <= 8'h10 ;
			data[45852] <= 8'h10 ;
			data[45853] <= 8'h10 ;
			data[45854] <= 8'h10 ;
			data[45855] <= 8'h10 ;
			data[45856] <= 8'h10 ;
			data[45857] <= 8'h10 ;
			data[45858] <= 8'h10 ;
			data[45859] <= 8'h10 ;
			data[45860] <= 8'h10 ;
			data[45861] <= 8'h10 ;
			data[45862] <= 8'h10 ;
			data[45863] <= 8'h10 ;
			data[45864] <= 8'h10 ;
			data[45865] <= 8'h10 ;
			data[45866] <= 8'h10 ;
			data[45867] <= 8'h10 ;
			data[45868] <= 8'h10 ;
			data[45869] <= 8'h10 ;
			data[45870] <= 8'h10 ;
			data[45871] <= 8'h10 ;
			data[45872] <= 8'h10 ;
			data[45873] <= 8'h10 ;
			data[45874] <= 8'h10 ;
			data[45875] <= 8'h10 ;
			data[45876] <= 8'h10 ;
			data[45877] <= 8'h10 ;
			data[45878] <= 8'h10 ;
			data[45879] <= 8'h10 ;
			data[45880] <= 8'h10 ;
			data[45881] <= 8'h10 ;
			data[45882] <= 8'h10 ;
			data[45883] <= 8'h10 ;
			data[45884] <= 8'h10 ;
			data[45885] <= 8'h10 ;
			data[45886] <= 8'h10 ;
			data[45887] <= 8'h10 ;
			data[45888] <= 8'h10 ;
			data[45889] <= 8'h10 ;
			data[45890] <= 8'h10 ;
			data[45891] <= 8'h10 ;
			data[45892] <= 8'h10 ;
			data[45893] <= 8'h10 ;
			data[45894] <= 8'h10 ;
			data[45895] <= 8'h10 ;
			data[45896] <= 8'h10 ;
			data[45897] <= 8'h10 ;
			data[45898] <= 8'h10 ;
			data[45899] <= 8'h10 ;
			data[45900] <= 8'h10 ;
			data[45901] <= 8'h10 ;
			data[45902] <= 8'h10 ;
			data[45903] <= 8'h10 ;
			data[45904] <= 8'h10 ;
			data[45905] <= 8'h10 ;
			data[45906] <= 8'h10 ;
			data[45907] <= 8'h10 ;
			data[45908] <= 8'h10 ;
			data[45909] <= 8'h10 ;
			data[45910] <= 8'h10 ;
			data[45911] <= 8'h10 ;
			data[45912] <= 8'h10 ;
			data[45913] <= 8'h10 ;
			data[45914] <= 8'h10 ;
			data[45915] <= 8'h10 ;
			data[45916] <= 8'h10 ;
			data[45917] <= 8'h10 ;
			data[45918] <= 8'h10 ;
			data[45919] <= 8'h10 ;
			data[45920] <= 8'h10 ;
			data[45921] <= 8'h10 ;
			data[45922] <= 8'h10 ;
			data[45923] <= 8'h10 ;
			data[45924] <= 8'h10 ;
			data[45925] <= 8'h10 ;
			data[45926] <= 8'h10 ;
			data[45927] <= 8'h10 ;
			data[45928] <= 8'h10 ;
			data[45929] <= 8'h10 ;
			data[45930] <= 8'h10 ;
			data[45931] <= 8'h10 ;
			data[45932] <= 8'h10 ;
			data[45933] <= 8'h10 ;
			data[45934] <= 8'h10 ;
			data[45935] <= 8'h10 ;
			data[45936] <= 8'h10 ;
			data[45937] <= 8'h10 ;
			data[45938] <= 8'h10 ;
			data[45939] <= 8'h10 ;
			data[45940] <= 8'h10 ;
			data[45941] <= 8'h10 ;
			data[45942] <= 8'h10 ;
			data[45943] <= 8'h10 ;
			data[45944] <= 8'h10 ;
			data[45945] <= 8'h10 ;
			data[45946] <= 8'h10 ;
			data[45947] <= 8'h10 ;
			data[45948] <= 8'h10 ;
			data[45949] <= 8'h10 ;
			data[45950] <= 8'h10 ;
			data[45951] <= 8'h10 ;
			data[45952] <= 8'h10 ;
			data[45953] <= 8'h10 ;
			data[45954] <= 8'h10 ;
			data[45955] <= 8'h10 ;
			data[45956] <= 8'h10 ;
			data[45957] <= 8'h10 ;
			data[45958] <= 8'h10 ;
			data[45959] <= 8'h10 ;
			data[45960] <= 8'h10 ;
			data[45961] <= 8'h10 ;
			data[45962] <= 8'h10 ;
			data[45963] <= 8'h10 ;
			data[45964] <= 8'h10 ;
			data[45965] <= 8'h10 ;
			data[45966] <= 8'h10 ;
			data[45967] <= 8'h10 ;
			data[45968] <= 8'h10 ;
			data[45969] <= 8'h10 ;
			data[45970] <= 8'h10 ;
			data[45971] <= 8'h10 ;
			data[45972] <= 8'h10 ;
			data[45973] <= 8'h10 ;
			data[45974] <= 8'h10 ;
			data[45975] <= 8'h10 ;
			data[45976] <= 8'h10 ;
			data[45977] <= 8'h10 ;
			data[45978] <= 8'h10 ;
			data[45979] <= 8'h10 ;
			data[45980] <= 8'h10 ;
			data[45981] <= 8'h10 ;
			data[45982] <= 8'h10 ;
			data[45983] <= 8'h10 ;
			data[45984] <= 8'h10 ;
			data[45985] <= 8'h10 ;
			data[45986] <= 8'h10 ;
			data[45987] <= 8'h10 ;
			data[45988] <= 8'h10 ;
			data[45989] <= 8'h10 ;
			data[45990] <= 8'h10 ;
			data[45991] <= 8'h10 ;
			data[45992] <= 8'h10 ;
			data[45993] <= 8'h10 ;
			data[45994] <= 8'h10 ;
			data[45995] <= 8'h10 ;
			data[45996] <= 8'h10 ;
			data[45997] <= 8'h10 ;
			data[45998] <= 8'h10 ;
			data[45999] <= 8'h10 ;
			data[46000] <= 8'h10 ;
			data[46001] <= 8'h10 ;
			data[46002] <= 8'h10 ;
			data[46003] <= 8'h10 ;
			data[46004] <= 8'h10 ;
			data[46005] <= 8'h10 ;
			data[46006] <= 8'h10 ;
			data[46007] <= 8'h10 ;
			data[46008] <= 8'h10 ;
			data[46009] <= 8'h10 ;
			data[46010] <= 8'h10 ;
			data[46011] <= 8'h10 ;
			data[46012] <= 8'h10 ;
			data[46013] <= 8'h10 ;
			data[46014] <= 8'h10 ;
			data[46015] <= 8'h10 ;
			data[46016] <= 8'h10 ;
			data[46017] <= 8'h10 ;
			data[46018] <= 8'h10 ;
			data[46019] <= 8'h10 ;
			data[46020] <= 8'h10 ;
			data[46021] <= 8'h10 ;
			data[46022] <= 8'h10 ;
			data[46023] <= 8'h10 ;
			data[46024] <= 8'h10 ;
			data[46025] <= 8'h10 ;
			data[46026] <= 8'h10 ;
			data[46027] <= 8'h10 ;
			data[46028] <= 8'h10 ;
			data[46029] <= 8'h10 ;
			data[46030] <= 8'h10 ;
			data[46031] <= 8'h10 ;
			data[46032] <= 8'h10 ;
			data[46033] <= 8'h10 ;
			data[46034] <= 8'h10 ;
			data[46035] <= 8'h10 ;
			data[46036] <= 8'h10 ;
			data[46037] <= 8'h10 ;
			data[46038] <= 8'h10 ;
			data[46039] <= 8'h10 ;
			data[46040] <= 8'h10 ;
			data[46041] <= 8'h10 ;
			data[46042] <= 8'h10 ;
			data[46043] <= 8'h10 ;
			data[46044] <= 8'h10 ;
			data[46045] <= 8'h10 ;
			data[46046] <= 8'h10 ;
			data[46047] <= 8'h10 ;
			data[46048] <= 8'h10 ;
			data[46049] <= 8'h10 ;
			data[46050] <= 8'h10 ;
			data[46051] <= 8'h10 ;
			data[46052] <= 8'h10 ;
			data[46053] <= 8'h10 ;
			data[46054] <= 8'h10 ;
			data[46055] <= 8'h10 ;
			data[46056] <= 8'h10 ;
			data[46057] <= 8'h10 ;
			data[46058] <= 8'h10 ;
			data[46059] <= 8'h10 ;
			data[46060] <= 8'h10 ;
			data[46061] <= 8'h10 ;
			data[46062] <= 8'h10 ;
			data[46063] <= 8'h10 ;
			data[46064] <= 8'h10 ;
			data[46065] <= 8'h10 ;
			data[46066] <= 8'h10 ;
			data[46067] <= 8'h10 ;
			data[46068] <= 8'h10 ;
			data[46069] <= 8'h10 ;
			data[46070] <= 8'h10 ;
			data[46071] <= 8'h10 ;
			data[46072] <= 8'h10 ;
			data[46073] <= 8'h10 ;
			data[46074] <= 8'h10 ;
			data[46075] <= 8'h10 ;
			data[46076] <= 8'h10 ;
			data[46077] <= 8'h10 ;
			data[46078] <= 8'h10 ;
			data[46079] <= 8'h10 ;
			data[46080] <= 8'h10 ;
			data[46081] <= 8'h10 ;
			data[46082] <= 8'h10 ;
			data[46083] <= 8'h10 ;
			data[46084] <= 8'h10 ;
			data[46085] <= 8'h10 ;
			data[46086] <= 8'h10 ;
			data[46087] <= 8'h10 ;
			data[46088] <= 8'h10 ;
			data[46089] <= 8'h10 ;
			data[46090] <= 8'h10 ;
			data[46091] <= 8'h10 ;
			data[46092] <= 8'h10 ;
			data[46093] <= 8'h10 ;
			data[46094] <= 8'h10 ;
			data[46095] <= 8'h10 ;
			data[46096] <= 8'h10 ;
			data[46097] <= 8'h10 ;
			data[46098] <= 8'h10 ;
			data[46099] <= 8'h10 ;
			data[46100] <= 8'h10 ;
			data[46101] <= 8'h10 ;
			data[46102] <= 8'h10 ;
			data[46103] <= 8'h10 ;
			data[46104] <= 8'h10 ;
			data[46105] <= 8'h10 ;
			data[46106] <= 8'h10 ;
			data[46107] <= 8'h10 ;
			data[46108] <= 8'h10 ;
			data[46109] <= 8'h10 ;
			data[46110] <= 8'h10 ;
			data[46111] <= 8'h10 ;
			data[46112] <= 8'h10 ;
			data[46113] <= 8'h10 ;
			data[46114] <= 8'h10 ;
			data[46115] <= 8'h10 ;
			data[46116] <= 8'h10 ;
			data[46117] <= 8'h10 ;
			data[46118] <= 8'h10 ;
			data[46119] <= 8'h10 ;
			data[46120] <= 8'h10 ;
			data[46121] <= 8'h10 ;
			data[46122] <= 8'h10 ;
			data[46123] <= 8'h10 ;
			data[46124] <= 8'h10 ;
			data[46125] <= 8'h10 ;
			data[46126] <= 8'h10 ;
			data[46127] <= 8'h10 ;
			data[46128] <= 8'h10 ;
			data[46129] <= 8'h10 ;
			data[46130] <= 8'h10 ;
			data[46131] <= 8'h10 ;
			data[46132] <= 8'h10 ;
			data[46133] <= 8'h10 ;
			data[46134] <= 8'h10 ;
			data[46135] <= 8'h10 ;
			data[46136] <= 8'h10 ;
			data[46137] <= 8'h10 ;
			data[46138] <= 8'h10 ;
			data[46139] <= 8'h10 ;
			data[46140] <= 8'h10 ;
			data[46141] <= 8'h10 ;
			data[46142] <= 8'h10 ;
			data[46143] <= 8'h10 ;
			data[46144] <= 8'h10 ;
			data[46145] <= 8'h10 ;
			data[46146] <= 8'h10 ;
			data[46147] <= 8'h10 ;
			data[46148] <= 8'h10 ;
			data[46149] <= 8'h10 ;
			data[46150] <= 8'h10 ;
			data[46151] <= 8'h10 ;
			data[46152] <= 8'h10 ;
			data[46153] <= 8'h10 ;
			data[46154] <= 8'h10 ;
			data[46155] <= 8'h10 ;
			data[46156] <= 8'h10 ;
			data[46157] <= 8'h10 ;
			data[46158] <= 8'h10 ;
			data[46159] <= 8'h10 ;
			data[46160] <= 8'h10 ;
			data[46161] <= 8'h10 ;
			data[46162] <= 8'h10 ;
			data[46163] <= 8'h10 ;
			data[46164] <= 8'h10 ;
			data[46165] <= 8'h10 ;
			data[46166] <= 8'h10 ;
			data[46167] <= 8'h10 ;
			data[46168] <= 8'h10 ;
			data[46169] <= 8'h10 ;
			data[46170] <= 8'h10 ;
			data[46171] <= 8'h10 ;
			data[46172] <= 8'h10 ;
			data[46173] <= 8'h10 ;
			data[46174] <= 8'h10 ;
			data[46175] <= 8'h10 ;
			data[46176] <= 8'h10 ;
			data[46177] <= 8'h10 ;
			data[46178] <= 8'h10 ;
			data[46179] <= 8'h10 ;
			data[46180] <= 8'h10 ;
			data[46181] <= 8'h10 ;
			data[46182] <= 8'h10 ;
			data[46183] <= 8'h10 ;
			data[46184] <= 8'h10 ;
			data[46185] <= 8'h10 ;
			data[46186] <= 8'h10 ;
			data[46187] <= 8'h10 ;
			data[46188] <= 8'h10 ;
			data[46189] <= 8'h10 ;
			data[46190] <= 8'h10 ;
			data[46191] <= 8'h10 ;
			data[46192] <= 8'h10 ;
			data[46193] <= 8'h10 ;
			data[46194] <= 8'h10 ;
			data[46195] <= 8'h10 ;
			data[46196] <= 8'h10 ;
			data[46197] <= 8'h10 ;
			data[46198] <= 8'h10 ;
			data[46199] <= 8'h10 ;
			data[46200] <= 8'h10 ;
			data[46201] <= 8'h10 ;
			data[46202] <= 8'h10 ;
			data[46203] <= 8'h10 ;
			data[46204] <= 8'h10 ;
			data[46205] <= 8'h10 ;
			data[46206] <= 8'h10 ;
			data[46207] <= 8'h10 ;
			data[46208] <= 8'h10 ;
			data[46209] <= 8'h10 ;
			data[46210] <= 8'h10 ;
			data[46211] <= 8'h10 ;
			data[46212] <= 8'h10 ;
			data[46213] <= 8'h10 ;
			data[46214] <= 8'h10 ;
			data[46215] <= 8'h10 ;
			data[46216] <= 8'h10 ;
			data[46217] <= 8'h10 ;
			data[46218] <= 8'h10 ;
			data[46219] <= 8'h10 ;
			data[46220] <= 8'h10 ;
			data[46221] <= 8'h10 ;
			data[46222] <= 8'h10 ;
			data[46223] <= 8'h10 ;
			data[46224] <= 8'h10 ;
			data[46225] <= 8'h10 ;
			data[46226] <= 8'h10 ;
			data[46227] <= 8'h10 ;
			data[46228] <= 8'h10 ;
			data[46229] <= 8'h10 ;
			data[46230] <= 8'h10 ;
			data[46231] <= 8'h10 ;
			data[46232] <= 8'h10 ;
			data[46233] <= 8'h10 ;
			data[46234] <= 8'h10 ;
			data[46235] <= 8'h10 ;
			data[46236] <= 8'h10 ;
			data[46237] <= 8'h10 ;
			data[46238] <= 8'h10 ;
			data[46239] <= 8'h10 ;
			data[46240] <= 8'h10 ;
			data[46241] <= 8'h10 ;
			data[46242] <= 8'h10 ;
			data[46243] <= 8'h10 ;
			data[46244] <= 8'h10 ;
			data[46245] <= 8'h10 ;
			data[46246] <= 8'h10 ;
			data[46247] <= 8'h10 ;
			data[46248] <= 8'h10 ;
			data[46249] <= 8'h10 ;
			data[46250] <= 8'h10 ;
			data[46251] <= 8'h10 ;
			data[46252] <= 8'h10 ;
			data[46253] <= 8'h10 ;
			data[46254] <= 8'h10 ;
			data[46255] <= 8'h10 ;
			data[46256] <= 8'h10 ;
			data[46257] <= 8'h10 ;
			data[46258] <= 8'h10 ;
			data[46259] <= 8'h10 ;
			data[46260] <= 8'h10 ;
			data[46261] <= 8'h10 ;
			data[46262] <= 8'h10 ;
			data[46263] <= 8'h10 ;
			data[46264] <= 8'h10 ;
			data[46265] <= 8'h10 ;
			data[46266] <= 8'h10 ;
			data[46267] <= 8'h10 ;
			data[46268] <= 8'h10 ;
			data[46269] <= 8'h10 ;
			data[46270] <= 8'h10 ;
			data[46271] <= 8'h10 ;
			data[46272] <= 8'h10 ;
			data[46273] <= 8'h10 ;
			data[46274] <= 8'h10 ;
			data[46275] <= 8'h10 ;
			data[46276] <= 8'h10 ;
			data[46277] <= 8'h10 ;
			data[46278] <= 8'h10 ;
			data[46279] <= 8'h10 ;
			data[46280] <= 8'h10 ;
			data[46281] <= 8'h10 ;
			data[46282] <= 8'h10 ;
			data[46283] <= 8'h10 ;
			data[46284] <= 8'h10 ;
			data[46285] <= 8'h10 ;
			data[46286] <= 8'h10 ;
			data[46287] <= 8'h10 ;
			data[46288] <= 8'h10 ;
			data[46289] <= 8'h10 ;
			data[46290] <= 8'h10 ;
			data[46291] <= 8'h10 ;
			data[46292] <= 8'h10 ;
			data[46293] <= 8'h10 ;
			data[46294] <= 8'h10 ;
			data[46295] <= 8'h10 ;
			data[46296] <= 8'h10 ;
			data[46297] <= 8'h10 ;
			data[46298] <= 8'h10 ;
			data[46299] <= 8'h10 ;
			data[46300] <= 8'h10 ;
			data[46301] <= 8'h10 ;
			data[46302] <= 8'h10 ;
			data[46303] <= 8'h10 ;
			data[46304] <= 8'h10 ;
			data[46305] <= 8'h10 ;
			data[46306] <= 8'h10 ;
			data[46307] <= 8'h10 ;
			data[46308] <= 8'h10 ;
			data[46309] <= 8'h10 ;
			data[46310] <= 8'h10 ;
			data[46311] <= 8'h10 ;
			data[46312] <= 8'h10 ;
			data[46313] <= 8'h10 ;
			data[46314] <= 8'h10 ;
			data[46315] <= 8'h10 ;
			data[46316] <= 8'h10 ;
			data[46317] <= 8'h10 ;
			data[46318] <= 8'h10 ;
			data[46319] <= 8'h10 ;
			data[46320] <= 8'h10 ;
			data[46321] <= 8'h10 ;
			data[46322] <= 8'h10 ;
			data[46323] <= 8'h10 ;
			data[46324] <= 8'h10 ;
			data[46325] <= 8'h10 ;
			data[46326] <= 8'h10 ;
			data[46327] <= 8'h10 ;
			data[46328] <= 8'h10 ;
			data[46329] <= 8'h10 ;
			data[46330] <= 8'h10 ;
			data[46331] <= 8'h10 ;
			data[46332] <= 8'h10 ;
			data[46333] <= 8'h10 ;
			data[46334] <= 8'h10 ;
			data[46335] <= 8'h10 ;
			data[46336] <= 8'h10 ;
			data[46337] <= 8'h10 ;
			data[46338] <= 8'h10 ;
			data[46339] <= 8'h10 ;
			data[46340] <= 8'h10 ;
			data[46341] <= 8'h10 ;
			data[46342] <= 8'h10 ;
			data[46343] <= 8'h10 ;
			data[46344] <= 8'h10 ;
			data[46345] <= 8'h10 ;
			data[46346] <= 8'h10 ;
			data[46347] <= 8'h10 ;
			data[46348] <= 8'h10 ;
			data[46349] <= 8'h10 ;
			data[46350] <= 8'h10 ;
			data[46351] <= 8'h10 ;
			data[46352] <= 8'h10 ;
			data[46353] <= 8'h10 ;
			data[46354] <= 8'h10 ;
			data[46355] <= 8'h10 ;
			data[46356] <= 8'h10 ;
			data[46357] <= 8'h10 ;
			data[46358] <= 8'h10 ;
			data[46359] <= 8'h10 ;
			data[46360] <= 8'h10 ;
			data[46361] <= 8'h10 ;
			data[46362] <= 8'h10 ;
			data[46363] <= 8'h10 ;
			data[46364] <= 8'h10 ;
			data[46365] <= 8'h10 ;
			data[46366] <= 8'h10 ;
			data[46367] <= 8'h10 ;
			data[46368] <= 8'h10 ;
			data[46369] <= 8'h10 ;
			data[46370] <= 8'h10 ;
			data[46371] <= 8'h10 ;
			data[46372] <= 8'h10 ;
			data[46373] <= 8'h10 ;
			data[46374] <= 8'h10 ;
			data[46375] <= 8'h10 ;
			data[46376] <= 8'h10 ;
			data[46377] <= 8'h10 ;
			data[46378] <= 8'h10 ;
			data[46379] <= 8'h10 ;
			data[46380] <= 8'h10 ;
			data[46381] <= 8'h10 ;
			data[46382] <= 8'h10 ;
			data[46383] <= 8'h10 ;
			data[46384] <= 8'h10 ;
			data[46385] <= 8'h10 ;
			data[46386] <= 8'h10 ;
			data[46387] <= 8'h10 ;
			data[46388] <= 8'h10 ;
			data[46389] <= 8'h10 ;
			data[46390] <= 8'h10 ;
			data[46391] <= 8'h10 ;
			data[46392] <= 8'h10 ;
			data[46393] <= 8'h10 ;
			data[46394] <= 8'h10 ;
			data[46395] <= 8'h10 ;
			data[46396] <= 8'h10 ;
			data[46397] <= 8'h10 ;
			data[46398] <= 8'h10 ;
			data[46399] <= 8'h10 ;
			data[46400] <= 8'h10 ;
			data[46401] <= 8'h10 ;
			data[46402] <= 8'h10 ;
			data[46403] <= 8'h10 ;
			data[46404] <= 8'h10 ;
			data[46405] <= 8'h10 ;
			data[46406] <= 8'h10 ;
			data[46407] <= 8'h10 ;
			data[46408] <= 8'h10 ;
			data[46409] <= 8'h10 ;
			data[46410] <= 8'h10 ;
			data[46411] <= 8'h10 ;
			data[46412] <= 8'h10 ;
			data[46413] <= 8'h10 ;
			data[46414] <= 8'h10 ;
			data[46415] <= 8'h10 ;
			data[46416] <= 8'h10 ;
			data[46417] <= 8'h10 ;
			data[46418] <= 8'h10 ;
			data[46419] <= 8'h10 ;
			data[46420] <= 8'h10 ;
			data[46421] <= 8'h10 ;
			data[46422] <= 8'h10 ;
			data[46423] <= 8'h10 ;
			data[46424] <= 8'h10 ;
			data[46425] <= 8'h10 ;
			data[46426] <= 8'h10 ;
			data[46427] <= 8'h10 ;
			data[46428] <= 8'h10 ;
			data[46429] <= 8'h10 ;
			data[46430] <= 8'h10 ;
			data[46431] <= 8'h10 ;
			data[46432] <= 8'h10 ;
			data[46433] <= 8'h10 ;
			data[46434] <= 8'h10 ;
			data[46435] <= 8'h10 ;
			data[46436] <= 8'h10 ;
			data[46437] <= 8'h10 ;
			data[46438] <= 8'h10 ;
			data[46439] <= 8'h10 ;
			data[46440] <= 8'h10 ;
			data[46441] <= 8'h10 ;
			data[46442] <= 8'h10 ;
			data[46443] <= 8'h10 ;
			data[46444] <= 8'h10 ;
			data[46445] <= 8'h10 ;
			data[46446] <= 8'h10 ;
			data[46447] <= 8'h10 ;
			data[46448] <= 8'h10 ;
			data[46449] <= 8'h10 ;
			data[46450] <= 8'h10 ;
			data[46451] <= 8'h10 ;
			data[46452] <= 8'h10 ;
			data[46453] <= 8'h10 ;
			data[46454] <= 8'h10 ;
			data[46455] <= 8'h10 ;
			data[46456] <= 8'h10 ;
			data[46457] <= 8'h10 ;
			data[46458] <= 8'h10 ;
			data[46459] <= 8'h10 ;
			data[46460] <= 8'h10 ;
			data[46461] <= 8'h10 ;
			data[46462] <= 8'h10 ;
			data[46463] <= 8'h10 ;
			data[46464] <= 8'h10 ;
			data[46465] <= 8'h10 ;
			data[46466] <= 8'h10 ;
			data[46467] <= 8'h10 ;
			data[46468] <= 8'h10 ;
			data[46469] <= 8'h10 ;
			data[46470] <= 8'h10 ;
			data[46471] <= 8'h10 ;
			data[46472] <= 8'h10 ;
			data[46473] <= 8'h10 ;
			data[46474] <= 8'h10 ;
			data[46475] <= 8'h10 ;
			data[46476] <= 8'h10 ;
			data[46477] <= 8'h10 ;
			data[46478] <= 8'h10 ;
			data[46479] <= 8'h10 ;
			data[46480] <= 8'h10 ;
			data[46481] <= 8'h10 ;
			data[46482] <= 8'h10 ;
			data[46483] <= 8'h10 ;
			data[46484] <= 8'h10 ;
			data[46485] <= 8'h10 ;
			data[46486] <= 8'h10 ;
			data[46487] <= 8'h10 ;
			data[46488] <= 8'h10 ;
			data[46489] <= 8'h10 ;
			data[46490] <= 8'h10 ;
			data[46491] <= 8'h10 ;
			data[46492] <= 8'h10 ;
			data[46493] <= 8'h10 ;
			data[46494] <= 8'h10 ;
			data[46495] <= 8'h10 ;
			data[46496] <= 8'h10 ;
			data[46497] <= 8'h10 ;
			data[46498] <= 8'h10 ;
			data[46499] <= 8'h10 ;
			data[46500] <= 8'h10 ;
			data[46501] <= 8'h10 ;
			data[46502] <= 8'h10 ;
			data[46503] <= 8'h10 ;
			data[46504] <= 8'h10 ;
			data[46505] <= 8'h10 ;
			data[46506] <= 8'h10 ;
			data[46507] <= 8'h10 ;
			data[46508] <= 8'h10 ;
			data[46509] <= 8'h10 ;
			data[46510] <= 8'h10 ;
			data[46511] <= 8'h10 ;
			data[46512] <= 8'h10 ;
			data[46513] <= 8'h10 ;
			data[46514] <= 8'h10 ;
			data[46515] <= 8'h10 ;
			data[46516] <= 8'h10 ;
			data[46517] <= 8'h10 ;
			data[46518] <= 8'h10 ;
			data[46519] <= 8'h10 ;
			data[46520] <= 8'h10 ;
			data[46521] <= 8'h10 ;
			data[46522] <= 8'h10 ;
			data[46523] <= 8'h10 ;
			data[46524] <= 8'h10 ;
			data[46525] <= 8'h10 ;
			data[46526] <= 8'h10 ;
			data[46527] <= 8'h10 ;
			data[46528] <= 8'h10 ;
			data[46529] <= 8'h10 ;
			data[46530] <= 8'h10 ;
			data[46531] <= 8'h10 ;
			data[46532] <= 8'h10 ;
			data[46533] <= 8'h10 ;
			data[46534] <= 8'h10 ;
			data[46535] <= 8'h10 ;
			data[46536] <= 8'h10 ;
			data[46537] <= 8'h10 ;
			data[46538] <= 8'h10 ;
			data[46539] <= 8'h10 ;
			data[46540] <= 8'h10 ;
			data[46541] <= 8'h10 ;
			data[46542] <= 8'h10 ;
			data[46543] <= 8'h10 ;
			data[46544] <= 8'h10 ;
			data[46545] <= 8'h10 ;
			data[46546] <= 8'h10 ;
			data[46547] <= 8'h10 ;
			data[46548] <= 8'h10 ;
			data[46549] <= 8'h10 ;
			data[46550] <= 8'h10 ;
			data[46551] <= 8'h10 ;
			data[46552] <= 8'h10 ;
			data[46553] <= 8'h10 ;
			data[46554] <= 8'h10 ;
			data[46555] <= 8'h10 ;
			data[46556] <= 8'h10 ;
			data[46557] <= 8'h10 ;
			data[46558] <= 8'h10 ;
			data[46559] <= 8'h10 ;
			data[46560] <= 8'h10 ;
			data[46561] <= 8'h10 ;
			data[46562] <= 8'h10 ;
			data[46563] <= 8'h10 ;
			data[46564] <= 8'h10 ;
			data[46565] <= 8'h10 ;
			data[46566] <= 8'h10 ;
			data[46567] <= 8'h10 ;
			data[46568] <= 8'h10 ;
			data[46569] <= 8'h10 ;
			data[46570] <= 8'h10 ;
			data[46571] <= 8'h10 ;
			data[46572] <= 8'h10 ;
			data[46573] <= 8'h10 ;
			data[46574] <= 8'h10 ;
			data[46575] <= 8'h10 ;
			data[46576] <= 8'h10 ;
			data[46577] <= 8'h10 ;
			data[46578] <= 8'h10 ;
			data[46579] <= 8'h10 ;
			data[46580] <= 8'h10 ;
			data[46581] <= 8'h10 ;
			data[46582] <= 8'h10 ;
			data[46583] <= 8'h10 ;
			data[46584] <= 8'h10 ;
			data[46585] <= 8'h10 ;
			data[46586] <= 8'h10 ;
			data[46587] <= 8'h10 ;
			data[46588] <= 8'h10 ;
			data[46589] <= 8'h10 ;
			data[46590] <= 8'h10 ;
			data[46591] <= 8'h10 ;
			data[46592] <= 8'h10 ;
			data[46593] <= 8'h10 ;
			data[46594] <= 8'h10 ;
			data[46595] <= 8'h10 ;
			data[46596] <= 8'h10 ;
			data[46597] <= 8'h10 ;
			data[46598] <= 8'h10 ;
			data[46599] <= 8'h10 ;
			data[46600] <= 8'h10 ;
			data[46601] <= 8'h10 ;
			data[46602] <= 8'h10 ;
			data[46603] <= 8'h10 ;
			data[46604] <= 8'h10 ;
			data[46605] <= 8'h10 ;
			data[46606] <= 8'h10 ;
			data[46607] <= 8'h10 ;
			data[46608] <= 8'h10 ;
			data[46609] <= 8'h10 ;
			data[46610] <= 8'h10 ;
			data[46611] <= 8'h10 ;
			data[46612] <= 8'h10 ;
			data[46613] <= 8'h10 ;
			data[46614] <= 8'h10 ;
			data[46615] <= 8'h10 ;
			data[46616] <= 8'h10 ;
			data[46617] <= 8'h10 ;
			data[46618] <= 8'h10 ;
			data[46619] <= 8'h10 ;
			data[46620] <= 8'h10 ;
			data[46621] <= 8'h10 ;
			data[46622] <= 8'h10 ;
			data[46623] <= 8'h10 ;
			data[46624] <= 8'h10 ;
			data[46625] <= 8'h10 ;
			data[46626] <= 8'h10 ;
			data[46627] <= 8'h10 ;
			data[46628] <= 8'h10 ;
			data[46629] <= 8'h10 ;
			data[46630] <= 8'h10 ;
			data[46631] <= 8'h10 ;
			data[46632] <= 8'h10 ;
			data[46633] <= 8'h10 ;
			data[46634] <= 8'h10 ;
			data[46635] <= 8'h10 ;
			data[46636] <= 8'h10 ;
			data[46637] <= 8'h10 ;
			data[46638] <= 8'h10 ;
			data[46639] <= 8'h10 ;
			data[46640] <= 8'h10 ;
			data[46641] <= 8'h10 ;
			data[46642] <= 8'h10 ;
			data[46643] <= 8'h10 ;
			data[46644] <= 8'h10 ;
			data[46645] <= 8'h10 ;
			data[46646] <= 8'h10 ;
			data[46647] <= 8'h10 ;
			data[46648] <= 8'h10 ;
			data[46649] <= 8'h10 ;
			data[46650] <= 8'h10 ;
			data[46651] <= 8'h10 ;
			data[46652] <= 8'h10 ;
			data[46653] <= 8'h10 ;
			data[46654] <= 8'h10 ;
			data[46655] <= 8'h10 ;
			data[46656] <= 8'h10 ;
			data[46657] <= 8'h10 ;
			data[46658] <= 8'h10 ;
			data[46659] <= 8'h10 ;
			data[46660] <= 8'h10 ;
			data[46661] <= 8'h10 ;
			data[46662] <= 8'h10 ;
			data[46663] <= 8'h10 ;
			data[46664] <= 8'h10 ;
			data[46665] <= 8'h10 ;
			data[46666] <= 8'h10 ;
			data[46667] <= 8'h10 ;
			data[46668] <= 8'h10 ;
			data[46669] <= 8'h10 ;
			data[46670] <= 8'h10 ;
			data[46671] <= 8'h10 ;
			data[46672] <= 8'h10 ;
			data[46673] <= 8'h10 ;
			data[46674] <= 8'h10 ;
			data[46675] <= 8'h10 ;
			data[46676] <= 8'h10 ;
			data[46677] <= 8'h10 ;
			data[46678] <= 8'h10 ;
			data[46679] <= 8'h10 ;
			data[46680] <= 8'h10 ;
			data[46681] <= 8'h10 ;
			data[46682] <= 8'h10 ;
			data[46683] <= 8'h10 ;
			data[46684] <= 8'h10 ;
			data[46685] <= 8'h10 ;
			data[46686] <= 8'h10 ;
			data[46687] <= 8'h10 ;
			data[46688] <= 8'h10 ;
			data[46689] <= 8'h10 ;
			data[46690] <= 8'h10 ;
			data[46691] <= 8'h10 ;
			data[46692] <= 8'h10 ;
			data[46693] <= 8'h10 ;
			data[46694] <= 8'h10 ;
			data[46695] <= 8'h10 ;
			data[46696] <= 8'h10 ;
			data[46697] <= 8'h10 ;
			data[46698] <= 8'h10 ;
			data[46699] <= 8'h10 ;
			data[46700] <= 8'h10 ;
			data[46701] <= 8'h10 ;
			data[46702] <= 8'h10 ;
			data[46703] <= 8'h10 ;
			data[46704] <= 8'h10 ;
			data[46705] <= 8'h10 ;
			data[46706] <= 8'h10 ;
			data[46707] <= 8'h10 ;
			data[46708] <= 8'h10 ;
			data[46709] <= 8'h10 ;
			data[46710] <= 8'h10 ;
			data[46711] <= 8'h10 ;
			data[46712] <= 8'h10 ;
			data[46713] <= 8'h10 ;
			data[46714] <= 8'h10 ;
			data[46715] <= 8'h10 ;
			data[46716] <= 8'h10 ;
			data[46717] <= 8'h10 ;
			data[46718] <= 8'h10 ;
			data[46719] <= 8'h10 ;
			data[46720] <= 8'h10 ;
			data[46721] <= 8'h10 ;
			data[46722] <= 8'h10 ;
			data[46723] <= 8'h10 ;
			data[46724] <= 8'h10 ;
			data[46725] <= 8'h10 ;
			data[46726] <= 8'h10 ;
			data[46727] <= 8'h10 ;
			data[46728] <= 8'h10 ;
			data[46729] <= 8'h10 ;
			data[46730] <= 8'h10 ;
			data[46731] <= 8'h10 ;
			data[46732] <= 8'h10 ;
			data[46733] <= 8'h10 ;
			data[46734] <= 8'h10 ;
			data[46735] <= 8'h10 ;
			data[46736] <= 8'h10 ;
			data[46737] <= 8'h10 ;
			data[46738] <= 8'h10 ;
			data[46739] <= 8'h10 ;
			data[46740] <= 8'h10 ;
			data[46741] <= 8'h10 ;
			data[46742] <= 8'h10 ;
			data[46743] <= 8'h10 ;
			data[46744] <= 8'h10 ;
			data[46745] <= 8'h10 ;
			data[46746] <= 8'h10 ;
			data[46747] <= 8'h10 ;
			data[46748] <= 8'h10 ;
			data[46749] <= 8'h10 ;
			data[46750] <= 8'h10 ;
			data[46751] <= 8'h10 ;
			data[46752] <= 8'h10 ;
			data[46753] <= 8'h10 ;
			data[46754] <= 8'h10 ;
			data[46755] <= 8'h10 ;
			data[46756] <= 8'h10 ;
			data[46757] <= 8'h10 ;
			data[46758] <= 8'h10 ;
			data[46759] <= 8'h10 ;
			data[46760] <= 8'h10 ;
			data[46761] <= 8'h10 ;
			data[46762] <= 8'h10 ;
			data[46763] <= 8'h10 ;
			data[46764] <= 8'h10 ;
			data[46765] <= 8'h10 ;
			data[46766] <= 8'h10 ;
			data[46767] <= 8'h10 ;
			data[46768] <= 8'h10 ;
			data[46769] <= 8'h10 ;
			data[46770] <= 8'h10 ;
			data[46771] <= 8'h10 ;
			data[46772] <= 8'h10 ;
			data[46773] <= 8'h10 ;
			data[46774] <= 8'h10 ;
			data[46775] <= 8'h10 ;
			data[46776] <= 8'h10 ;
			data[46777] <= 8'h10 ;
			data[46778] <= 8'h10 ;
			data[46779] <= 8'h10 ;
			data[46780] <= 8'h10 ;
			data[46781] <= 8'h10 ;
			data[46782] <= 8'h10 ;
			data[46783] <= 8'h10 ;
			data[46784] <= 8'h10 ;
			data[46785] <= 8'h10 ;
			data[46786] <= 8'h10 ;
			data[46787] <= 8'h10 ;
			data[46788] <= 8'h10 ;
			data[46789] <= 8'h10 ;
			data[46790] <= 8'h10 ;
			data[46791] <= 8'h10 ;
			data[46792] <= 8'h10 ;
			data[46793] <= 8'h10 ;
			data[46794] <= 8'h10 ;
			data[46795] <= 8'h10 ;
			data[46796] <= 8'h10 ;
			data[46797] <= 8'h10 ;
			data[46798] <= 8'h10 ;
			data[46799] <= 8'h10 ;
			data[46800] <= 8'h10 ;
			data[46801] <= 8'h10 ;
			data[46802] <= 8'h10 ;
			data[46803] <= 8'h10 ;
			data[46804] <= 8'h10 ;
			data[46805] <= 8'h10 ;
			data[46806] <= 8'h10 ;
			data[46807] <= 8'h10 ;
			data[46808] <= 8'h10 ;
			data[46809] <= 8'h10 ;
			data[46810] <= 8'h10 ;
			data[46811] <= 8'h10 ;
			data[46812] <= 8'h10 ;
			data[46813] <= 8'h10 ;
			data[46814] <= 8'h10 ;
			data[46815] <= 8'h10 ;
			data[46816] <= 8'h10 ;
			data[46817] <= 8'h10 ;
			data[46818] <= 8'h10 ;
			data[46819] <= 8'h10 ;
			data[46820] <= 8'h10 ;
			data[46821] <= 8'h10 ;
			data[46822] <= 8'h10 ;
			data[46823] <= 8'h10 ;
			data[46824] <= 8'h10 ;
			data[46825] <= 8'h10 ;
			data[46826] <= 8'h10 ;
			data[46827] <= 8'h10 ;
			data[46828] <= 8'h10 ;
			data[46829] <= 8'h10 ;
			data[46830] <= 8'h10 ;
			data[46831] <= 8'h10 ;
			data[46832] <= 8'h10 ;
			data[46833] <= 8'h10 ;
			data[46834] <= 8'h10 ;
			data[46835] <= 8'h10 ;
			data[46836] <= 8'h10 ;
			data[46837] <= 8'h10 ;
			data[46838] <= 8'h10 ;
			data[46839] <= 8'h10 ;
			data[46840] <= 8'h10 ;
			data[46841] <= 8'h10 ;
			data[46842] <= 8'h10 ;
			data[46843] <= 8'h10 ;
			data[46844] <= 8'h10 ;
			data[46845] <= 8'h10 ;
			data[46846] <= 8'h10 ;
			data[46847] <= 8'h10 ;
			data[46848] <= 8'h10 ;
			data[46849] <= 8'h10 ;
			data[46850] <= 8'h10 ;
			data[46851] <= 8'h10 ;
			data[46852] <= 8'h10 ;
			data[46853] <= 8'h10 ;
			data[46854] <= 8'h10 ;
			data[46855] <= 8'h10 ;
			data[46856] <= 8'h10 ;
			data[46857] <= 8'h10 ;
			data[46858] <= 8'h10 ;
			data[46859] <= 8'h10 ;
			data[46860] <= 8'h10 ;
			data[46861] <= 8'h10 ;
			data[46862] <= 8'h10 ;
			data[46863] <= 8'h10 ;
			data[46864] <= 8'h10 ;
			data[46865] <= 8'h10 ;
			data[46866] <= 8'h10 ;
			data[46867] <= 8'h10 ;
			data[46868] <= 8'h10 ;
			data[46869] <= 8'h10 ;
			data[46870] <= 8'h10 ;
			data[46871] <= 8'h10 ;
			data[46872] <= 8'h10 ;
			data[46873] <= 8'h10 ;
			data[46874] <= 8'h10 ;
			data[46875] <= 8'h10 ;
			data[46876] <= 8'h10 ;
			data[46877] <= 8'h10 ;
			data[46878] <= 8'h10 ;
			data[46879] <= 8'h10 ;
			data[46880] <= 8'h10 ;
			data[46881] <= 8'h10 ;
			data[46882] <= 8'h10 ;
			data[46883] <= 8'h10 ;
			data[46884] <= 8'h10 ;
			data[46885] <= 8'h10 ;
			data[46886] <= 8'h10 ;
			data[46887] <= 8'h10 ;
			data[46888] <= 8'h10 ;
			data[46889] <= 8'h10 ;
			data[46890] <= 8'h10 ;
			data[46891] <= 8'h10 ;
			data[46892] <= 8'h10 ;
			data[46893] <= 8'h10 ;
			data[46894] <= 8'h10 ;
			data[46895] <= 8'h10 ;
			data[46896] <= 8'h10 ;
			data[46897] <= 8'h10 ;
			data[46898] <= 8'h10 ;
			data[46899] <= 8'h10 ;
			data[46900] <= 8'h10 ;
			data[46901] <= 8'h10 ;
			data[46902] <= 8'h10 ;
			data[46903] <= 8'h10 ;
			data[46904] <= 8'h10 ;
			data[46905] <= 8'h10 ;
			data[46906] <= 8'h10 ;
			data[46907] <= 8'h10 ;
			data[46908] <= 8'h10 ;
			data[46909] <= 8'h10 ;
			data[46910] <= 8'h10 ;
			data[46911] <= 8'h10 ;
			data[46912] <= 8'h10 ;
			data[46913] <= 8'h10 ;
			data[46914] <= 8'h10 ;
			data[46915] <= 8'h10 ;
			data[46916] <= 8'h10 ;
			data[46917] <= 8'h10 ;
			data[46918] <= 8'h10 ;
			data[46919] <= 8'h10 ;
			data[46920] <= 8'h10 ;
			data[46921] <= 8'h10 ;
			data[46922] <= 8'h10 ;
			data[46923] <= 8'h10 ;
			data[46924] <= 8'h10 ;
			data[46925] <= 8'h10 ;
			data[46926] <= 8'h10 ;
			data[46927] <= 8'h10 ;
			data[46928] <= 8'h10 ;
			data[46929] <= 8'h10 ;
			data[46930] <= 8'h10 ;
			data[46931] <= 8'h10 ;
			data[46932] <= 8'h10 ;
			data[46933] <= 8'h10 ;
			data[46934] <= 8'h10 ;
			data[46935] <= 8'h10 ;
			data[46936] <= 8'h10 ;
			data[46937] <= 8'h10 ;
			data[46938] <= 8'h10 ;
			data[46939] <= 8'h10 ;
			data[46940] <= 8'h10 ;
			data[46941] <= 8'h10 ;
			data[46942] <= 8'h10 ;
			data[46943] <= 8'h10 ;
			data[46944] <= 8'h10 ;
			data[46945] <= 8'h10 ;
			data[46946] <= 8'h10 ;
			data[46947] <= 8'h10 ;
			data[46948] <= 8'h10 ;
			data[46949] <= 8'h10 ;
			data[46950] <= 8'h10 ;
			data[46951] <= 8'h10 ;
			data[46952] <= 8'h10 ;
			data[46953] <= 8'h10 ;
			data[46954] <= 8'h10 ;
			data[46955] <= 8'h10 ;
			data[46956] <= 8'h10 ;
			data[46957] <= 8'h10 ;
			data[46958] <= 8'h10 ;
			data[46959] <= 8'h10 ;
			data[46960] <= 8'h10 ;
			data[46961] <= 8'h10 ;
			data[46962] <= 8'h10 ;
			data[46963] <= 8'h10 ;
			data[46964] <= 8'h10 ;
			data[46965] <= 8'h10 ;
			data[46966] <= 8'h10 ;
			data[46967] <= 8'h10 ;
			data[46968] <= 8'h10 ;
			data[46969] <= 8'h10 ;
			data[46970] <= 8'h10 ;
			data[46971] <= 8'h10 ;
			data[46972] <= 8'h10 ;
			data[46973] <= 8'h10 ;
			data[46974] <= 8'h10 ;
			data[46975] <= 8'h10 ;
			data[46976] <= 8'h10 ;
			data[46977] <= 8'h10 ;
			data[46978] <= 8'h10 ;
			data[46979] <= 8'h10 ;
			data[46980] <= 8'h10 ;
			data[46981] <= 8'h10 ;
			data[46982] <= 8'h10 ;
			data[46983] <= 8'h10 ;
			data[46984] <= 8'h10 ;
			data[46985] <= 8'h10 ;
			data[46986] <= 8'h10 ;
			data[46987] <= 8'h10 ;
			data[46988] <= 8'h10 ;
			data[46989] <= 8'h10 ;
			data[46990] <= 8'h10 ;
			data[46991] <= 8'h10 ;
			data[46992] <= 8'h10 ;
			data[46993] <= 8'h10 ;
			data[46994] <= 8'h10 ;
			data[46995] <= 8'h10 ;
			data[46996] <= 8'h10 ;
			data[46997] <= 8'h10 ;
			data[46998] <= 8'h10 ;
			data[46999] <= 8'h10 ;
			data[47000] <= 8'h10 ;
			data[47001] <= 8'h10 ;
			data[47002] <= 8'h10 ;
			data[47003] <= 8'h10 ;
			data[47004] <= 8'h10 ;
			data[47005] <= 8'h10 ;
			data[47006] <= 8'h10 ;
			data[47007] <= 8'h10 ;
			data[47008] <= 8'h10 ;
			data[47009] <= 8'h10 ;
			data[47010] <= 8'h10 ;
			data[47011] <= 8'h10 ;
			data[47012] <= 8'h10 ;
			data[47013] <= 8'h10 ;
			data[47014] <= 8'h10 ;
			data[47015] <= 8'h10 ;
			data[47016] <= 8'h10 ;
			data[47017] <= 8'h10 ;
			data[47018] <= 8'h10 ;
			data[47019] <= 8'h10 ;
			data[47020] <= 8'h10 ;
			data[47021] <= 8'h10 ;
			data[47022] <= 8'h10 ;
			data[47023] <= 8'h10 ;
			data[47024] <= 8'h10 ;
			data[47025] <= 8'h10 ;
			data[47026] <= 8'h10 ;
			data[47027] <= 8'h10 ;
			data[47028] <= 8'h10 ;
			data[47029] <= 8'h10 ;
			data[47030] <= 8'h10 ;
			data[47031] <= 8'h10 ;
			data[47032] <= 8'h10 ;
			data[47033] <= 8'h10 ;
			data[47034] <= 8'h10 ;
			data[47035] <= 8'h10 ;
			data[47036] <= 8'h10 ;
			data[47037] <= 8'h10 ;
			data[47038] <= 8'h10 ;
			data[47039] <= 8'h10 ;
			data[47040] <= 8'h10 ;
			data[47041] <= 8'h10 ;
			data[47042] <= 8'h10 ;
			data[47043] <= 8'h10 ;
			data[47044] <= 8'h10 ;
			data[47045] <= 8'h10 ;
			data[47046] <= 8'h10 ;
			data[47047] <= 8'h10 ;
			data[47048] <= 8'h10 ;
			data[47049] <= 8'h10 ;
			data[47050] <= 8'h10 ;
			data[47051] <= 8'h10 ;
			data[47052] <= 8'h10 ;
			data[47053] <= 8'h10 ;
			data[47054] <= 8'h10 ;
			data[47055] <= 8'h10 ;
			data[47056] <= 8'h10 ;
			data[47057] <= 8'h10 ;
			data[47058] <= 8'h10 ;
			data[47059] <= 8'h10 ;
			data[47060] <= 8'h10 ;
			data[47061] <= 8'h10 ;
			data[47062] <= 8'h10 ;
			data[47063] <= 8'h10 ;
			data[47064] <= 8'h10 ;
			data[47065] <= 8'h10 ;
			data[47066] <= 8'h10 ;
			data[47067] <= 8'h10 ;
			data[47068] <= 8'h10 ;
			data[47069] <= 8'h10 ;
			data[47070] <= 8'h10 ;
			data[47071] <= 8'h10 ;
			data[47072] <= 8'h10 ;
			data[47073] <= 8'h10 ;
			data[47074] <= 8'h10 ;
			data[47075] <= 8'h10 ;
			data[47076] <= 8'h10 ;
			data[47077] <= 8'h10 ;
			data[47078] <= 8'h10 ;
			data[47079] <= 8'h10 ;
			data[47080] <= 8'h10 ;
			data[47081] <= 8'h10 ;
			data[47082] <= 8'h10 ;
			data[47083] <= 8'h10 ;
			data[47084] <= 8'h10 ;
			data[47085] <= 8'h10 ;
			data[47086] <= 8'h10 ;
			data[47087] <= 8'h10 ;
			data[47088] <= 8'h10 ;
			data[47089] <= 8'h10 ;
			data[47090] <= 8'h10 ;
			data[47091] <= 8'h10 ;
			data[47092] <= 8'h10 ;
			data[47093] <= 8'h10 ;
			data[47094] <= 8'h10 ;
			data[47095] <= 8'h10 ;
			data[47096] <= 8'h10 ;
			data[47097] <= 8'h10 ;
			data[47098] <= 8'h10 ;
			data[47099] <= 8'h10 ;
			data[47100] <= 8'h10 ;
			data[47101] <= 8'h10 ;
			data[47102] <= 8'h10 ;
			data[47103] <= 8'h10 ;
			data[47104] <= 8'h10 ;
			data[47105] <= 8'h10 ;
			data[47106] <= 8'h10 ;
			data[47107] <= 8'h10 ;
			data[47108] <= 8'h10 ;
			data[47109] <= 8'h10 ;
			data[47110] <= 8'h10 ;
			data[47111] <= 8'h10 ;
			data[47112] <= 8'h10 ;
			data[47113] <= 8'h10 ;
			data[47114] <= 8'h10 ;
			data[47115] <= 8'h10 ;
			data[47116] <= 8'h10 ;
			data[47117] <= 8'h10 ;
			data[47118] <= 8'h10 ;
			data[47119] <= 8'h10 ;
			data[47120] <= 8'h10 ;
			data[47121] <= 8'h10 ;
			data[47122] <= 8'h10 ;
			data[47123] <= 8'h10 ;
			data[47124] <= 8'h10 ;
			data[47125] <= 8'h10 ;
			data[47126] <= 8'h10 ;
			data[47127] <= 8'h10 ;
			data[47128] <= 8'h10 ;
			data[47129] <= 8'h10 ;
			data[47130] <= 8'h10 ;
			data[47131] <= 8'h10 ;
			data[47132] <= 8'h10 ;
			data[47133] <= 8'h10 ;
			data[47134] <= 8'h10 ;
			data[47135] <= 8'h10 ;
			data[47136] <= 8'h10 ;
			data[47137] <= 8'h10 ;
			data[47138] <= 8'h10 ;
			data[47139] <= 8'h10 ;
			data[47140] <= 8'h10 ;
			data[47141] <= 8'h10 ;
			data[47142] <= 8'h10 ;
			data[47143] <= 8'h10 ;
			data[47144] <= 8'h10 ;
			data[47145] <= 8'h10 ;
			data[47146] <= 8'h10 ;
			data[47147] <= 8'h10 ;
			data[47148] <= 8'h10 ;
			data[47149] <= 8'h10 ;
			data[47150] <= 8'h10 ;
			data[47151] <= 8'h10 ;
			data[47152] <= 8'h10 ;
			data[47153] <= 8'h10 ;
			data[47154] <= 8'h10 ;
			data[47155] <= 8'h10 ;
			data[47156] <= 8'h10 ;
			data[47157] <= 8'h10 ;
			data[47158] <= 8'h10 ;
			data[47159] <= 8'h10 ;
			data[47160] <= 8'h10 ;
			data[47161] <= 8'h10 ;
			data[47162] <= 8'h10 ;
			data[47163] <= 8'h10 ;
			data[47164] <= 8'h10 ;
			data[47165] <= 8'h10 ;
			data[47166] <= 8'h10 ;
			data[47167] <= 8'h10 ;
			data[47168] <= 8'h10 ;
			data[47169] <= 8'h10 ;
			data[47170] <= 8'h10 ;
			data[47171] <= 8'h10 ;
			data[47172] <= 8'h10 ;
			data[47173] <= 8'h10 ;
			data[47174] <= 8'h10 ;
			data[47175] <= 8'h10 ;
			data[47176] <= 8'h10 ;
			data[47177] <= 8'h10 ;
			data[47178] <= 8'h10 ;
			data[47179] <= 8'h10 ;
			data[47180] <= 8'h10 ;
			data[47181] <= 8'h10 ;
			data[47182] <= 8'h10 ;
			data[47183] <= 8'h10 ;
			data[47184] <= 8'h10 ;
			data[47185] <= 8'h10 ;
			data[47186] <= 8'h10 ;
			data[47187] <= 8'h10 ;
			data[47188] <= 8'h10 ;
			data[47189] <= 8'h10 ;
			data[47190] <= 8'h10 ;
			data[47191] <= 8'h10 ;
			data[47192] <= 8'h10 ;
			data[47193] <= 8'h10 ;
			data[47194] <= 8'h10 ;
			data[47195] <= 8'h10 ;
			data[47196] <= 8'h10 ;
			data[47197] <= 8'h10 ;
			data[47198] <= 8'h10 ;
			data[47199] <= 8'h10 ;
			data[47200] <= 8'h10 ;
			data[47201] <= 8'h10 ;
			data[47202] <= 8'h10 ;
			data[47203] <= 8'h10 ;
			data[47204] <= 8'h10 ;
			data[47205] <= 8'h10 ;
			data[47206] <= 8'h10 ;
			data[47207] <= 8'h10 ;
			data[47208] <= 8'h10 ;
			data[47209] <= 8'h10 ;
			data[47210] <= 8'h10 ;
			data[47211] <= 8'h10 ;
			data[47212] <= 8'h10 ;
			data[47213] <= 8'h10 ;
			data[47214] <= 8'h10 ;
			data[47215] <= 8'h10 ;
			data[47216] <= 8'h10 ;
			data[47217] <= 8'h10 ;
			data[47218] <= 8'h10 ;
			data[47219] <= 8'h10 ;
			data[47220] <= 8'h10 ;
			data[47221] <= 8'h10 ;
			data[47222] <= 8'h10 ;
			data[47223] <= 8'h10 ;
			data[47224] <= 8'h10 ;
			data[47225] <= 8'h10 ;
			data[47226] <= 8'h10 ;
			data[47227] <= 8'h10 ;
			data[47228] <= 8'h10 ;
			data[47229] <= 8'h10 ;
			data[47230] <= 8'h10 ;
			data[47231] <= 8'h10 ;
			data[47232] <= 8'h10 ;
			data[47233] <= 8'h10 ;
			data[47234] <= 8'h10 ;
			data[47235] <= 8'h10 ;
			data[47236] <= 8'h10 ;
			data[47237] <= 8'h10 ;
			data[47238] <= 8'h10 ;
			data[47239] <= 8'h10 ;
			data[47240] <= 8'h10 ;
			data[47241] <= 8'h10 ;
			data[47242] <= 8'h10 ;
			data[47243] <= 8'h10 ;
			data[47244] <= 8'h10 ;
			data[47245] <= 8'h10 ;
			data[47246] <= 8'h10 ;
			data[47247] <= 8'h10 ;
			data[47248] <= 8'h10 ;
			data[47249] <= 8'h10 ;
			data[47250] <= 8'h10 ;
			data[47251] <= 8'h10 ;
			data[47252] <= 8'h10 ;
			data[47253] <= 8'h10 ;
			data[47254] <= 8'h10 ;
			data[47255] <= 8'h10 ;
			data[47256] <= 8'h10 ;
			data[47257] <= 8'h10 ;
			data[47258] <= 8'h10 ;
			data[47259] <= 8'h10 ;
			data[47260] <= 8'h10 ;
			data[47261] <= 8'h10 ;
			data[47262] <= 8'h10 ;
			data[47263] <= 8'h10 ;
			data[47264] <= 8'h10 ;
			data[47265] <= 8'h10 ;
			data[47266] <= 8'h10 ;
			data[47267] <= 8'h10 ;
			data[47268] <= 8'h10 ;
			data[47269] <= 8'h10 ;
			data[47270] <= 8'h10 ;
			data[47271] <= 8'h10 ;
			data[47272] <= 8'h10 ;
			data[47273] <= 8'h10 ;
			data[47274] <= 8'h10 ;
			data[47275] <= 8'h10 ;
			data[47276] <= 8'h10 ;
			data[47277] <= 8'h10 ;
			data[47278] <= 8'h10 ;
			data[47279] <= 8'h10 ;
			data[47280] <= 8'h10 ;
			data[47281] <= 8'h10 ;
			data[47282] <= 8'h10 ;
			data[47283] <= 8'h10 ;
			data[47284] <= 8'h10 ;
			data[47285] <= 8'h10 ;
			data[47286] <= 8'h10 ;
			data[47287] <= 8'h10 ;
			data[47288] <= 8'h10 ;
			data[47289] <= 8'h10 ;
			data[47290] <= 8'h10 ;
			data[47291] <= 8'h10 ;
			data[47292] <= 8'h10 ;
			data[47293] <= 8'h10 ;
			data[47294] <= 8'h10 ;
			data[47295] <= 8'h10 ;
			data[47296] <= 8'h10 ;
			data[47297] <= 8'h10 ;
			data[47298] <= 8'h10 ;
			data[47299] <= 8'h10 ;
			data[47300] <= 8'h10 ;
			data[47301] <= 8'h10 ;
			data[47302] <= 8'h10 ;
			data[47303] <= 8'h10 ;
			data[47304] <= 8'h10 ;
			data[47305] <= 8'h10 ;
			data[47306] <= 8'h10 ;
			data[47307] <= 8'h10 ;
			data[47308] <= 8'h10 ;
			data[47309] <= 8'h10 ;
			data[47310] <= 8'h10 ;
			data[47311] <= 8'h10 ;
			data[47312] <= 8'h10 ;
			data[47313] <= 8'h10 ;
			data[47314] <= 8'h10 ;
			data[47315] <= 8'h10 ;
			data[47316] <= 8'h10 ;
			data[47317] <= 8'h10 ;
			data[47318] <= 8'h10 ;
			data[47319] <= 8'h10 ;
			data[47320] <= 8'h10 ;
			data[47321] <= 8'h10 ;
			data[47322] <= 8'h10 ;
			data[47323] <= 8'h10 ;
			data[47324] <= 8'h10 ;
			data[47325] <= 8'h10 ;
			data[47326] <= 8'h10 ;
			data[47327] <= 8'h10 ;
			data[47328] <= 8'h10 ;
			data[47329] <= 8'h10 ;
			data[47330] <= 8'h10 ;
			data[47331] <= 8'h10 ;
			data[47332] <= 8'h10 ;
			data[47333] <= 8'h10 ;
			data[47334] <= 8'h10 ;
			data[47335] <= 8'h10 ;
			data[47336] <= 8'h10 ;
			data[47337] <= 8'h10 ;
			data[47338] <= 8'h10 ;
			data[47339] <= 8'h10 ;
			data[47340] <= 8'h10 ;
			data[47341] <= 8'h10 ;
			data[47342] <= 8'h10 ;
			data[47343] <= 8'h10 ;
			data[47344] <= 8'h10 ;
			data[47345] <= 8'h10 ;
			data[47346] <= 8'h10 ;
			data[47347] <= 8'h10 ;
			data[47348] <= 8'h10 ;
			data[47349] <= 8'h10 ;
			data[47350] <= 8'h10 ;
			data[47351] <= 8'h10 ;
			data[47352] <= 8'h10 ;
			data[47353] <= 8'h10 ;
			data[47354] <= 8'h10 ;
			data[47355] <= 8'h10 ;
			data[47356] <= 8'h10 ;
			data[47357] <= 8'h10 ;
			data[47358] <= 8'h10 ;
			data[47359] <= 8'h10 ;
			data[47360] <= 8'h10 ;
			data[47361] <= 8'h10 ;
			data[47362] <= 8'h10 ;
			data[47363] <= 8'h10 ;
			data[47364] <= 8'h10 ;
			data[47365] <= 8'h10 ;
			data[47366] <= 8'h10 ;
			data[47367] <= 8'h10 ;
			data[47368] <= 8'h10 ;
			data[47369] <= 8'h10 ;
			data[47370] <= 8'h10 ;
			data[47371] <= 8'h10 ;
			data[47372] <= 8'h10 ;
			data[47373] <= 8'h10 ;
			data[47374] <= 8'h10 ;
			data[47375] <= 8'h10 ;
			data[47376] <= 8'h10 ;
			data[47377] <= 8'h10 ;
			data[47378] <= 8'h10 ;
			data[47379] <= 8'h10 ;
			data[47380] <= 8'h10 ;
			data[47381] <= 8'h10 ;
			data[47382] <= 8'h10 ;
			data[47383] <= 8'h10 ;
			data[47384] <= 8'h10 ;
			data[47385] <= 8'h10 ;
			data[47386] <= 8'h10 ;
			data[47387] <= 8'h10 ;
			data[47388] <= 8'h10 ;
			data[47389] <= 8'h10 ;
			data[47390] <= 8'h10 ;
			data[47391] <= 8'h10 ;
			data[47392] <= 8'h10 ;
			data[47393] <= 8'h10 ;
			data[47394] <= 8'h10 ;
			data[47395] <= 8'h10 ;
			data[47396] <= 8'h10 ;
			data[47397] <= 8'h10 ;
			data[47398] <= 8'h10 ;
			data[47399] <= 8'h10 ;
			data[47400] <= 8'h10 ;
			data[47401] <= 8'h10 ;
			data[47402] <= 8'h10 ;
			data[47403] <= 8'h10 ;
			data[47404] <= 8'h10 ;
			data[47405] <= 8'h10 ;
			data[47406] <= 8'h10 ;
			data[47407] <= 8'h10 ;
			data[47408] <= 8'h10 ;
			data[47409] <= 8'h10 ;
			data[47410] <= 8'h10 ;
			data[47411] <= 8'h10 ;
			data[47412] <= 8'h10 ;
			data[47413] <= 8'h10 ;
			data[47414] <= 8'h10 ;
			data[47415] <= 8'h10 ;
			data[47416] <= 8'h10 ;
			data[47417] <= 8'h10 ;
			data[47418] <= 8'h10 ;
			data[47419] <= 8'h10 ;
			data[47420] <= 8'h10 ;
			data[47421] <= 8'h10 ;
			data[47422] <= 8'h10 ;
			data[47423] <= 8'h10 ;
			data[47424] <= 8'h10 ;
			data[47425] <= 8'h10 ;
			data[47426] <= 8'h10 ;
			data[47427] <= 8'h10 ;
			data[47428] <= 8'h10 ;
			data[47429] <= 8'h10 ;
			data[47430] <= 8'h10 ;
			data[47431] <= 8'h10 ;
			data[47432] <= 8'h10 ;
			data[47433] <= 8'h10 ;
			data[47434] <= 8'h10 ;
			data[47435] <= 8'h10 ;
			data[47436] <= 8'h10 ;
			data[47437] <= 8'h10 ;
			data[47438] <= 8'h10 ;
			data[47439] <= 8'h10 ;
			data[47440] <= 8'h10 ;
			data[47441] <= 8'h10 ;
			data[47442] <= 8'h10 ;
			data[47443] <= 8'h10 ;
			data[47444] <= 8'h10 ;
			data[47445] <= 8'h10 ;
			data[47446] <= 8'h10 ;
			data[47447] <= 8'h10 ;
			data[47448] <= 8'h10 ;
			data[47449] <= 8'h10 ;
			data[47450] <= 8'h10 ;
			data[47451] <= 8'h10 ;
			data[47452] <= 8'h10 ;
			data[47453] <= 8'h10 ;
			data[47454] <= 8'h10 ;
			data[47455] <= 8'h10 ;
			data[47456] <= 8'h10 ;
			data[47457] <= 8'h10 ;
			data[47458] <= 8'h10 ;
			data[47459] <= 8'h10 ;
			data[47460] <= 8'h10 ;
			data[47461] <= 8'h10 ;
			data[47462] <= 8'h10 ;
			data[47463] <= 8'h10 ;
			data[47464] <= 8'h10 ;
			data[47465] <= 8'h10 ;
			data[47466] <= 8'h10 ;
			data[47467] <= 8'h10 ;
			data[47468] <= 8'h10 ;
			data[47469] <= 8'h10 ;
			data[47470] <= 8'h10 ;
			data[47471] <= 8'h10 ;
			data[47472] <= 8'h10 ;
			data[47473] <= 8'h10 ;
			data[47474] <= 8'h10 ;
			data[47475] <= 8'h10 ;
			data[47476] <= 8'h10 ;
			data[47477] <= 8'h10 ;
			data[47478] <= 8'h10 ;
			data[47479] <= 8'h10 ;
			data[47480] <= 8'h10 ;
			data[47481] <= 8'h10 ;
			data[47482] <= 8'h10 ;
			data[47483] <= 8'h10 ;
			data[47484] <= 8'h10 ;
			data[47485] <= 8'h10 ;
			data[47486] <= 8'h10 ;
			data[47487] <= 8'h10 ;
			data[47488] <= 8'h10 ;
			data[47489] <= 8'h10 ;
			data[47490] <= 8'h10 ;
			data[47491] <= 8'h10 ;
			data[47492] <= 8'h10 ;
			data[47493] <= 8'h10 ;
			data[47494] <= 8'h10 ;
			data[47495] <= 8'h10 ;
			data[47496] <= 8'h10 ;
			data[47497] <= 8'h10 ;
			data[47498] <= 8'h10 ;
			data[47499] <= 8'h10 ;
			data[47500] <= 8'h10 ;
			data[47501] <= 8'h10 ;
			data[47502] <= 8'h10 ;
			data[47503] <= 8'h10 ;
			data[47504] <= 8'h10 ;
			data[47505] <= 8'h10 ;
			data[47506] <= 8'h10 ;
			data[47507] <= 8'h10 ;
			data[47508] <= 8'h10 ;
			data[47509] <= 8'h10 ;
			data[47510] <= 8'h10 ;
			data[47511] <= 8'h10 ;
			data[47512] <= 8'h10 ;
			data[47513] <= 8'h10 ;
			data[47514] <= 8'h10 ;
			data[47515] <= 8'h10 ;
			data[47516] <= 8'h10 ;
			data[47517] <= 8'h10 ;
			data[47518] <= 8'h10 ;
			data[47519] <= 8'h10 ;
			data[47520] <= 8'h10 ;
			data[47521] <= 8'h10 ;
			data[47522] <= 8'h10 ;
			data[47523] <= 8'h10 ;
			data[47524] <= 8'h10 ;
			data[47525] <= 8'h10 ;
			data[47526] <= 8'h10 ;
			data[47527] <= 8'h10 ;
			data[47528] <= 8'h10 ;
			data[47529] <= 8'h10 ;
			data[47530] <= 8'h10 ;
			data[47531] <= 8'h10 ;
			data[47532] <= 8'h10 ;
			data[47533] <= 8'h10 ;
			data[47534] <= 8'h10 ;
			data[47535] <= 8'h10 ;
			data[47536] <= 8'h10 ;
			data[47537] <= 8'h10 ;
			data[47538] <= 8'h10 ;
			data[47539] <= 8'h10 ;
			data[47540] <= 8'h10 ;
			data[47541] <= 8'h10 ;
			data[47542] <= 8'h10 ;
			data[47543] <= 8'h10 ;
			data[47544] <= 8'h10 ;
			data[47545] <= 8'h10 ;
			data[47546] <= 8'h10 ;
			data[47547] <= 8'h10 ;
			data[47548] <= 8'h10 ;
			data[47549] <= 8'h10 ;
			data[47550] <= 8'h10 ;
			data[47551] <= 8'h10 ;
			data[47552] <= 8'h10 ;
			data[47553] <= 8'h10 ;
			data[47554] <= 8'h10 ;
			data[47555] <= 8'h10 ;
			data[47556] <= 8'h10 ;
			data[47557] <= 8'h10 ;
			data[47558] <= 8'h10 ;
			data[47559] <= 8'h10 ;
			data[47560] <= 8'h10 ;
			data[47561] <= 8'h10 ;
			data[47562] <= 8'h10 ;
			data[47563] <= 8'h10 ;
			data[47564] <= 8'h10 ;
			data[47565] <= 8'h10 ;
			data[47566] <= 8'h10 ;
			data[47567] <= 8'h10 ;
			data[47568] <= 8'h10 ;
			data[47569] <= 8'h10 ;
			data[47570] <= 8'h10 ;
			data[47571] <= 8'h10 ;
			data[47572] <= 8'h10 ;
			data[47573] <= 8'h10 ;
			data[47574] <= 8'h10 ;
			data[47575] <= 8'h10 ;
			data[47576] <= 8'h10 ;
			data[47577] <= 8'h10 ;
			data[47578] <= 8'h10 ;
			data[47579] <= 8'h10 ;
			data[47580] <= 8'h10 ;
			data[47581] <= 8'h10 ;
			data[47582] <= 8'h10 ;
			data[47583] <= 8'h10 ;
			data[47584] <= 8'h10 ;
			data[47585] <= 8'h10 ;
			data[47586] <= 8'h10 ;
			data[47587] <= 8'h10 ;
			data[47588] <= 8'h10 ;
			data[47589] <= 8'h10 ;
			data[47590] <= 8'h10 ;
			data[47591] <= 8'h10 ;
			data[47592] <= 8'h10 ;
			data[47593] <= 8'h10 ;
			data[47594] <= 8'h10 ;
			data[47595] <= 8'h10 ;
			data[47596] <= 8'h10 ;
			data[47597] <= 8'h10 ;
			data[47598] <= 8'h10 ;
			data[47599] <= 8'h10 ;
			data[47600] <= 8'h10 ;
			data[47601] <= 8'h10 ;
			data[47602] <= 8'h10 ;
			data[47603] <= 8'h10 ;
			data[47604] <= 8'h10 ;
			data[47605] <= 8'h10 ;
			data[47606] <= 8'h10 ;
			data[47607] <= 8'h10 ;
			data[47608] <= 8'h10 ;
			data[47609] <= 8'h10 ;
			data[47610] <= 8'h10 ;
			data[47611] <= 8'h10 ;
			data[47612] <= 8'h10 ;
			data[47613] <= 8'h10 ;
			data[47614] <= 8'h10 ;
			data[47615] <= 8'h10 ;
			data[47616] <= 8'h10 ;
			data[47617] <= 8'h10 ;
			data[47618] <= 8'h10 ;
			data[47619] <= 8'h10 ;
			data[47620] <= 8'h10 ;
			data[47621] <= 8'h10 ;
			data[47622] <= 8'h10 ;
			data[47623] <= 8'h10 ;
			data[47624] <= 8'h10 ;
			data[47625] <= 8'h10 ;
			data[47626] <= 8'h10 ;
			data[47627] <= 8'h10 ;
			data[47628] <= 8'h10 ;
			data[47629] <= 8'h10 ;
			data[47630] <= 8'h10 ;
			data[47631] <= 8'h10 ;
			data[47632] <= 8'h10 ;
			data[47633] <= 8'h10 ;
			data[47634] <= 8'h10 ;
			data[47635] <= 8'h10 ;
			data[47636] <= 8'h10 ;
			data[47637] <= 8'h10 ;
			data[47638] <= 8'h10 ;
			data[47639] <= 8'h10 ;
			data[47640] <= 8'h10 ;
			data[47641] <= 8'h10 ;
			data[47642] <= 8'h10 ;
			data[47643] <= 8'h10 ;
			data[47644] <= 8'h10 ;
			data[47645] <= 8'h10 ;
			data[47646] <= 8'h10 ;
			data[47647] <= 8'h10 ;
			data[47648] <= 8'h10 ;
			data[47649] <= 8'h10 ;
			data[47650] <= 8'h10 ;
			data[47651] <= 8'h10 ;
			data[47652] <= 8'h10 ;
			data[47653] <= 8'h10 ;
			data[47654] <= 8'h10 ;
			data[47655] <= 8'h10 ;
			data[47656] <= 8'h10 ;
			data[47657] <= 8'h10 ;
			data[47658] <= 8'h10 ;
			data[47659] <= 8'h10 ;
			data[47660] <= 8'h10 ;
			data[47661] <= 8'h10 ;
			data[47662] <= 8'h10 ;
			data[47663] <= 8'h10 ;
			data[47664] <= 8'h10 ;
			data[47665] <= 8'h10 ;
			data[47666] <= 8'h10 ;
			data[47667] <= 8'h10 ;
			data[47668] <= 8'h10 ;
			data[47669] <= 8'h10 ;
			data[47670] <= 8'h10 ;
			data[47671] <= 8'h10 ;
			data[47672] <= 8'h10 ;
			data[47673] <= 8'h10 ;
			data[47674] <= 8'h10 ;
			data[47675] <= 8'h10 ;
			data[47676] <= 8'h10 ;
			data[47677] <= 8'h10 ;
			data[47678] <= 8'h10 ;
			data[47679] <= 8'h10 ;
			data[47680] <= 8'h10 ;
			data[47681] <= 8'h10 ;
			data[47682] <= 8'h10 ;
			data[47683] <= 8'h10 ;
			data[47684] <= 8'h10 ;
			data[47685] <= 8'h10 ;
			data[47686] <= 8'h10 ;
			data[47687] <= 8'h10 ;
			data[47688] <= 8'h10 ;
			data[47689] <= 8'h10 ;
			data[47690] <= 8'h10 ;
			data[47691] <= 8'h10 ;
			data[47692] <= 8'h10 ;
			data[47693] <= 8'h10 ;
			data[47694] <= 8'h10 ;
			data[47695] <= 8'h10 ;
			data[47696] <= 8'h10 ;
			data[47697] <= 8'h10 ;
			data[47698] <= 8'h10 ;
			data[47699] <= 8'h10 ;
			data[47700] <= 8'h10 ;
			data[47701] <= 8'h10 ;
			data[47702] <= 8'h10 ;
			data[47703] <= 8'h10 ;
			data[47704] <= 8'h10 ;
			data[47705] <= 8'h10 ;
			data[47706] <= 8'h10 ;
			data[47707] <= 8'h10 ;
			data[47708] <= 8'h10 ;
			data[47709] <= 8'h10 ;
			data[47710] <= 8'h10 ;
			data[47711] <= 8'h10 ;
			data[47712] <= 8'h10 ;
			data[47713] <= 8'h10 ;
			data[47714] <= 8'h10 ;
			data[47715] <= 8'h10 ;
			data[47716] <= 8'h10 ;
			data[47717] <= 8'h10 ;
			data[47718] <= 8'h10 ;
			data[47719] <= 8'h10 ;
			data[47720] <= 8'h10 ;
			data[47721] <= 8'h10 ;
			data[47722] <= 8'h10 ;
			data[47723] <= 8'h10 ;
			data[47724] <= 8'h10 ;
			data[47725] <= 8'h10 ;
			data[47726] <= 8'h10 ;
			data[47727] <= 8'h10 ;
			data[47728] <= 8'h10 ;
			data[47729] <= 8'h10 ;
			data[47730] <= 8'h10 ;
			data[47731] <= 8'h10 ;
			data[47732] <= 8'h10 ;
			data[47733] <= 8'h10 ;
			data[47734] <= 8'h10 ;
			data[47735] <= 8'h10 ;
			data[47736] <= 8'h10 ;
			data[47737] <= 8'h10 ;
			data[47738] <= 8'h10 ;
			data[47739] <= 8'h10 ;
			data[47740] <= 8'h10 ;
			data[47741] <= 8'h10 ;
			data[47742] <= 8'h10 ;
			data[47743] <= 8'h10 ;
			data[47744] <= 8'h10 ;
			data[47745] <= 8'h10 ;
			data[47746] <= 8'h10 ;
			data[47747] <= 8'h10 ;
			data[47748] <= 8'h10 ;
			data[47749] <= 8'h10 ;
			data[47750] <= 8'h10 ;
			data[47751] <= 8'h10 ;
			data[47752] <= 8'h10 ;
			data[47753] <= 8'h10 ;
			data[47754] <= 8'h10 ;
			data[47755] <= 8'h10 ;
			data[47756] <= 8'h10 ;
			data[47757] <= 8'h10 ;
			data[47758] <= 8'h10 ;
			data[47759] <= 8'h10 ;
			data[47760] <= 8'h10 ;
			data[47761] <= 8'h10 ;
			data[47762] <= 8'h10 ;
			data[47763] <= 8'h10 ;
			data[47764] <= 8'h10 ;
			data[47765] <= 8'h10 ;
			data[47766] <= 8'h10 ;
			data[47767] <= 8'h10 ;
			data[47768] <= 8'h10 ;
			data[47769] <= 8'h10 ;
			data[47770] <= 8'h10 ;
			data[47771] <= 8'h10 ;
			data[47772] <= 8'h10 ;
			data[47773] <= 8'h10 ;
			data[47774] <= 8'h10 ;
			data[47775] <= 8'h10 ;
			data[47776] <= 8'h10 ;
			data[47777] <= 8'h10 ;
			data[47778] <= 8'h10 ;
			data[47779] <= 8'h10 ;
			data[47780] <= 8'h10 ;
			data[47781] <= 8'h10 ;
			data[47782] <= 8'h10 ;
			data[47783] <= 8'h10 ;
			data[47784] <= 8'h10 ;
			data[47785] <= 8'h10 ;
			data[47786] <= 8'h10 ;
			data[47787] <= 8'h10 ;
			data[47788] <= 8'h10 ;
			data[47789] <= 8'h10 ;
			data[47790] <= 8'h10 ;
			data[47791] <= 8'h10 ;
			data[47792] <= 8'h10 ;
			data[47793] <= 8'h10 ;
			data[47794] <= 8'h10 ;
			data[47795] <= 8'h10 ;
			data[47796] <= 8'h10 ;
			data[47797] <= 8'h10 ;
			data[47798] <= 8'h10 ;
			data[47799] <= 8'h10 ;
			data[47800] <= 8'h10 ;
			data[47801] <= 8'h10 ;
			data[47802] <= 8'h10 ;
			data[47803] <= 8'h10 ;
			data[47804] <= 8'h10 ;
			data[47805] <= 8'h10 ;
			data[47806] <= 8'h10 ;
			data[47807] <= 8'h10 ;
			data[47808] <= 8'h10 ;
			data[47809] <= 8'h10 ;
			data[47810] <= 8'h10 ;
			data[47811] <= 8'h10 ;
			data[47812] <= 8'h10 ;
			data[47813] <= 8'h10 ;
			data[47814] <= 8'h10 ;
			data[47815] <= 8'h10 ;
			data[47816] <= 8'h10 ;
			data[47817] <= 8'h10 ;
			data[47818] <= 8'h10 ;
			data[47819] <= 8'h10 ;
			data[47820] <= 8'h10 ;
			data[47821] <= 8'h10 ;
			data[47822] <= 8'h10 ;
			data[47823] <= 8'h10 ;
			data[47824] <= 8'h10 ;
			data[47825] <= 8'h10 ;
			data[47826] <= 8'h10 ;
			data[47827] <= 8'h10 ;
			data[47828] <= 8'h10 ;
			data[47829] <= 8'h10 ;
			data[47830] <= 8'h10 ;
			data[47831] <= 8'h10 ;
			data[47832] <= 8'h10 ;
			data[47833] <= 8'h10 ;
			data[47834] <= 8'h10 ;
			data[47835] <= 8'h10 ;
			data[47836] <= 8'h10 ;
			data[47837] <= 8'h10 ;
			data[47838] <= 8'h10 ;
			data[47839] <= 8'h10 ;
			data[47840] <= 8'h10 ;
			data[47841] <= 8'h10 ;
			data[47842] <= 8'h10 ;
			data[47843] <= 8'h10 ;
			data[47844] <= 8'h10 ;
			data[47845] <= 8'h10 ;
			data[47846] <= 8'h10 ;
			data[47847] <= 8'h10 ;
			data[47848] <= 8'h10 ;
			data[47849] <= 8'h10 ;
			data[47850] <= 8'h10 ;
			data[47851] <= 8'h10 ;
			data[47852] <= 8'h10 ;
			data[47853] <= 8'h10 ;
			data[47854] <= 8'h10 ;
			data[47855] <= 8'h10 ;
			data[47856] <= 8'h10 ;
			data[47857] <= 8'h10 ;
			data[47858] <= 8'h10 ;
			data[47859] <= 8'h10 ;
			data[47860] <= 8'h10 ;
			data[47861] <= 8'h10 ;
			data[47862] <= 8'h10 ;
			data[47863] <= 8'h10 ;
			data[47864] <= 8'h10 ;
			data[47865] <= 8'h10 ;
			data[47866] <= 8'h10 ;
			data[47867] <= 8'h10 ;
			data[47868] <= 8'h10 ;
			data[47869] <= 8'h10 ;
			data[47870] <= 8'h10 ;
			data[47871] <= 8'h10 ;
			data[47872] <= 8'h10 ;
			data[47873] <= 8'h10 ;
			data[47874] <= 8'h10 ;
			data[47875] <= 8'h10 ;
			data[47876] <= 8'h10 ;
			data[47877] <= 8'h10 ;
			data[47878] <= 8'h10 ;
			data[47879] <= 8'h10 ;
			data[47880] <= 8'h10 ;
			data[47881] <= 8'h10 ;
			data[47882] <= 8'h10 ;
			data[47883] <= 8'h10 ;
			data[47884] <= 8'h10 ;
			data[47885] <= 8'h10 ;
			data[47886] <= 8'h10 ;
			data[47887] <= 8'h10 ;
			data[47888] <= 8'h10 ;
			data[47889] <= 8'h10 ;
			data[47890] <= 8'h10 ;
			data[47891] <= 8'h10 ;
			data[47892] <= 8'h10 ;
			data[47893] <= 8'h10 ;
			data[47894] <= 8'h10 ;
			data[47895] <= 8'h10 ;
			data[47896] <= 8'h10 ;
			data[47897] <= 8'h10 ;
			data[47898] <= 8'h10 ;
			data[47899] <= 8'h10 ;
			data[47900] <= 8'h10 ;
			data[47901] <= 8'h10 ;
			data[47902] <= 8'h10 ;
			data[47903] <= 8'h10 ;
			data[47904] <= 8'h10 ;
			data[47905] <= 8'h10 ;
			data[47906] <= 8'h10 ;
			data[47907] <= 8'h10 ;
			data[47908] <= 8'h10 ;
			data[47909] <= 8'h10 ;
			data[47910] <= 8'h10 ;
			data[47911] <= 8'h10 ;
			data[47912] <= 8'h10 ;
			data[47913] <= 8'h10 ;
			data[47914] <= 8'h10 ;
			data[47915] <= 8'h10 ;
			data[47916] <= 8'h10 ;
			data[47917] <= 8'h10 ;
			data[47918] <= 8'h10 ;
			data[47919] <= 8'h10 ;
			data[47920] <= 8'h10 ;
			data[47921] <= 8'h10 ;
			data[47922] <= 8'h10 ;
			data[47923] <= 8'h10 ;
			data[47924] <= 8'h10 ;
			data[47925] <= 8'h10 ;
			data[47926] <= 8'h10 ;
			data[47927] <= 8'h10 ;
			data[47928] <= 8'h10 ;
			data[47929] <= 8'h10 ;
			data[47930] <= 8'h10 ;
			data[47931] <= 8'h10 ;
			data[47932] <= 8'h10 ;
			data[47933] <= 8'h10 ;
			data[47934] <= 8'h10 ;
			data[47935] <= 8'h10 ;
			data[47936] <= 8'h10 ;
			data[47937] <= 8'h10 ;
			data[47938] <= 8'h10 ;
			data[47939] <= 8'h10 ;
			data[47940] <= 8'h10 ;
			data[47941] <= 8'h10 ;
			data[47942] <= 8'h10 ;
			data[47943] <= 8'h10 ;
			data[47944] <= 8'h10 ;
			data[47945] <= 8'h10 ;
			data[47946] <= 8'h10 ;
			data[47947] <= 8'h10 ;
			data[47948] <= 8'h10 ;
			data[47949] <= 8'h10 ;
			data[47950] <= 8'h10 ;
			data[47951] <= 8'h10 ;
			data[47952] <= 8'h10 ;
			data[47953] <= 8'h10 ;
			data[47954] <= 8'h10 ;
			data[47955] <= 8'h10 ;
			data[47956] <= 8'h10 ;
			data[47957] <= 8'h10 ;
			data[47958] <= 8'h10 ;
			data[47959] <= 8'h10 ;
			data[47960] <= 8'h10 ;
			data[47961] <= 8'h10 ;
			data[47962] <= 8'h10 ;
			data[47963] <= 8'h10 ;
			data[47964] <= 8'h10 ;
			data[47965] <= 8'h10 ;
			data[47966] <= 8'h10 ;
			data[47967] <= 8'h10 ;
			data[47968] <= 8'h10 ;
			data[47969] <= 8'h10 ;
			data[47970] <= 8'h10 ;
			data[47971] <= 8'h10 ;
			data[47972] <= 8'h10 ;
			data[47973] <= 8'h10 ;
			data[47974] <= 8'h10 ;
			data[47975] <= 8'h10 ;
			data[47976] <= 8'h10 ;
			data[47977] <= 8'h10 ;
			data[47978] <= 8'h10 ;
			data[47979] <= 8'h10 ;
			data[47980] <= 8'h10 ;
			data[47981] <= 8'h10 ;
			data[47982] <= 8'h10 ;
			data[47983] <= 8'h10 ;
			data[47984] <= 8'h10 ;
			data[47985] <= 8'h10 ;
			data[47986] <= 8'h10 ;
			data[47987] <= 8'h10 ;
			data[47988] <= 8'h10 ;
			data[47989] <= 8'h10 ;
			data[47990] <= 8'h10 ;
			data[47991] <= 8'h10 ;
			data[47992] <= 8'h10 ;
			data[47993] <= 8'h10 ;
			data[47994] <= 8'h10 ;
			data[47995] <= 8'h10 ;
			data[47996] <= 8'h10 ;
			data[47997] <= 8'h10 ;
			data[47998] <= 8'h10 ;
			data[47999] <= 8'h10 ;
			data[48000] <= 8'h10 ;
			data[48001] <= 8'h10 ;
			data[48002] <= 8'h10 ;
			data[48003] <= 8'h10 ;
			data[48004] <= 8'h10 ;
			data[48005] <= 8'h10 ;
			data[48006] <= 8'h10 ;
			data[48007] <= 8'h10 ;
			data[48008] <= 8'h10 ;
			data[48009] <= 8'h10 ;
			data[48010] <= 8'h10 ;
			data[48011] <= 8'h10 ;
			data[48012] <= 8'h10 ;
			data[48013] <= 8'h10 ;
			data[48014] <= 8'h10 ;
			data[48015] <= 8'h10 ;
			data[48016] <= 8'h10 ;
			data[48017] <= 8'h10 ;
			data[48018] <= 8'h10 ;
			data[48019] <= 8'h10 ;
			data[48020] <= 8'h10 ;
			data[48021] <= 8'h10 ;
			data[48022] <= 8'h10 ;
			data[48023] <= 8'h10 ;
			data[48024] <= 8'h10 ;
			data[48025] <= 8'h10 ;
			data[48026] <= 8'h10 ;
			data[48027] <= 8'h10 ;
			data[48028] <= 8'h10 ;
			data[48029] <= 8'h10 ;
			data[48030] <= 8'h10 ;
			data[48031] <= 8'h10 ;
			data[48032] <= 8'h10 ;
			data[48033] <= 8'h10 ;
			data[48034] <= 8'h10 ;
			data[48035] <= 8'h10 ;
			data[48036] <= 8'h10 ;
			data[48037] <= 8'h10 ;
			data[48038] <= 8'h10 ;
			data[48039] <= 8'h10 ;
			data[48040] <= 8'h10 ;
			data[48041] <= 8'h10 ;
			data[48042] <= 8'h10 ;
			data[48043] <= 8'h10 ;
			data[48044] <= 8'h10 ;
			data[48045] <= 8'h10 ;
			data[48046] <= 8'h10 ;
			data[48047] <= 8'h10 ;
			data[48048] <= 8'h10 ;
			data[48049] <= 8'h10 ;
			data[48050] <= 8'h10 ;
			data[48051] <= 8'h10 ;
			data[48052] <= 8'h10 ;
			data[48053] <= 8'h10 ;
			data[48054] <= 8'h10 ;
			data[48055] <= 8'h10 ;
			data[48056] <= 8'h10 ;
			data[48057] <= 8'h10 ;
			data[48058] <= 8'h10 ;
			data[48059] <= 8'h10 ;
			data[48060] <= 8'h10 ;
			data[48061] <= 8'h10 ;
			data[48062] <= 8'h10 ;
			data[48063] <= 8'h10 ;
			data[48064] <= 8'h10 ;
			data[48065] <= 8'h10 ;
			data[48066] <= 8'h10 ;
			data[48067] <= 8'h10 ;
			data[48068] <= 8'h10 ;
			data[48069] <= 8'h10 ;
			data[48070] <= 8'h10 ;
			data[48071] <= 8'h10 ;
			data[48072] <= 8'h10 ;
			data[48073] <= 8'h10 ;
			data[48074] <= 8'h10 ;
			data[48075] <= 8'h10 ;
			data[48076] <= 8'h10 ;
			data[48077] <= 8'h10 ;
			data[48078] <= 8'h10 ;
			data[48079] <= 8'h10 ;
			data[48080] <= 8'h10 ;
			data[48081] <= 8'h10 ;
			data[48082] <= 8'h10 ;
			data[48083] <= 8'h10 ;
			data[48084] <= 8'h10 ;
			data[48085] <= 8'h10 ;
			data[48086] <= 8'h10 ;
			data[48087] <= 8'h10 ;
			data[48088] <= 8'h10 ;
			data[48089] <= 8'h10 ;
			data[48090] <= 8'h10 ;
			data[48091] <= 8'h10 ;
			data[48092] <= 8'h10 ;
			data[48093] <= 8'h10 ;
			data[48094] <= 8'h10 ;
			data[48095] <= 8'h10 ;
			data[48096] <= 8'h10 ;
			data[48097] <= 8'h10 ;
			data[48098] <= 8'h10 ;
			data[48099] <= 8'h10 ;
			data[48100] <= 8'h10 ;
			data[48101] <= 8'h10 ;
			data[48102] <= 8'h10 ;
			data[48103] <= 8'h10 ;
			data[48104] <= 8'h10 ;
			data[48105] <= 8'h10 ;
			data[48106] <= 8'h10 ;
			data[48107] <= 8'h10 ;
			data[48108] <= 8'h10 ;
			data[48109] <= 8'h10 ;
			data[48110] <= 8'h10 ;
			data[48111] <= 8'h10 ;
			data[48112] <= 8'h10 ;
			data[48113] <= 8'h10 ;
			data[48114] <= 8'h10 ;
			data[48115] <= 8'h10 ;
			data[48116] <= 8'h10 ;
			data[48117] <= 8'h10 ;
			data[48118] <= 8'h10 ;
			data[48119] <= 8'h10 ;
			data[48120] <= 8'h10 ;
			data[48121] <= 8'h10 ;
			data[48122] <= 8'h10 ;
			data[48123] <= 8'h10 ;
			data[48124] <= 8'h10 ;
			data[48125] <= 8'h10 ;
			data[48126] <= 8'h10 ;
			data[48127] <= 8'h10 ;
			data[48128] <= 8'h10 ;
			data[48129] <= 8'h10 ;
			data[48130] <= 8'h10 ;
			data[48131] <= 8'h10 ;
			data[48132] <= 8'h10 ;
			data[48133] <= 8'h10 ;
			data[48134] <= 8'h10 ;
			data[48135] <= 8'h10 ;
			data[48136] <= 8'h10 ;
			data[48137] <= 8'h10 ;
			data[48138] <= 8'h10 ;
			data[48139] <= 8'h10 ;
			data[48140] <= 8'h10 ;
			data[48141] <= 8'h10 ;
			data[48142] <= 8'h10 ;
			data[48143] <= 8'h10 ;
			data[48144] <= 8'h10 ;
			data[48145] <= 8'h10 ;
			data[48146] <= 8'h10 ;
			data[48147] <= 8'h10 ;
			data[48148] <= 8'h10 ;
			data[48149] <= 8'h10 ;
			data[48150] <= 8'h10 ;
			data[48151] <= 8'h10 ;
			data[48152] <= 8'h10 ;
			data[48153] <= 8'h10 ;
			data[48154] <= 8'h10 ;
			data[48155] <= 8'h10 ;
			data[48156] <= 8'h10 ;
			data[48157] <= 8'h10 ;
			data[48158] <= 8'h10 ;
			data[48159] <= 8'h10 ;
			data[48160] <= 8'h10 ;
			data[48161] <= 8'h10 ;
			data[48162] <= 8'h10 ;
			data[48163] <= 8'h10 ;
			data[48164] <= 8'h10 ;
			data[48165] <= 8'h10 ;
			data[48166] <= 8'h10 ;
			data[48167] <= 8'h10 ;
			data[48168] <= 8'h10 ;
			data[48169] <= 8'h10 ;
			data[48170] <= 8'h10 ;
			data[48171] <= 8'h10 ;
			data[48172] <= 8'h10 ;
			data[48173] <= 8'h10 ;
			data[48174] <= 8'h10 ;
			data[48175] <= 8'h10 ;
			data[48176] <= 8'h10 ;
			data[48177] <= 8'h10 ;
			data[48178] <= 8'h10 ;
			data[48179] <= 8'h10 ;
			data[48180] <= 8'h10 ;
			data[48181] <= 8'h10 ;
			data[48182] <= 8'h10 ;
			data[48183] <= 8'h10 ;
			data[48184] <= 8'h10 ;
			data[48185] <= 8'h10 ;
			data[48186] <= 8'h10 ;
			data[48187] <= 8'h10 ;
			data[48188] <= 8'h10 ;
			data[48189] <= 8'h10 ;
			data[48190] <= 8'h10 ;
			data[48191] <= 8'h10 ;
			data[48192] <= 8'h10 ;
			data[48193] <= 8'h10 ;
			data[48194] <= 8'h10 ;
			data[48195] <= 8'h10 ;
			data[48196] <= 8'h10 ;
			data[48197] <= 8'h10 ;
			data[48198] <= 8'h10 ;
			data[48199] <= 8'h10 ;
			data[48200] <= 8'h10 ;
			data[48201] <= 8'h10 ;
			data[48202] <= 8'h10 ;
			data[48203] <= 8'h10 ;
			data[48204] <= 8'h10 ;
			data[48205] <= 8'h10 ;
			data[48206] <= 8'h10 ;
			data[48207] <= 8'h10 ;
			data[48208] <= 8'h10 ;
			data[48209] <= 8'h10 ;
			data[48210] <= 8'h10 ;
			data[48211] <= 8'h10 ;
			data[48212] <= 8'h10 ;
			data[48213] <= 8'h10 ;
			data[48214] <= 8'h10 ;
			data[48215] <= 8'h10 ;
			data[48216] <= 8'h10 ;
			data[48217] <= 8'h10 ;
			data[48218] <= 8'h10 ;
			data[48219] <= 8'h10 ;
			data[48220] <= 8'h10 ;
			data[48221] <= 8'h10 ;
			data[48222] <= 8'h10 ;
			data[48223] <= 8'h10 ;
			data[48224] <= 8'h10 ;
			data[48225] <= 8'h10 ;
			data[48226] <= 8'h10 ;
			data[48227] <= 8'h10 ;
			data[48228] <= 8'h10 ;
			data[48229] <= 8'h10 ;
			data[48230] <= 8'h10 ;
			data[48231] <= 8'h10 ;
			data[48232] <= 8'h10 ;
			data[48233] <= 8'h10 ;
			data[48234] <= 8'h10 ;
			data[48235] <= 8'h10 ;
			data[48236] <= 8'h10 ;
			data[48237] <= 8'h10 ;
			data[48238] <= 8'h10 ;
			data[48239] <= 8'h10 ;
			data[48240] <= 8'h10 ;
			data[48241] <= 8'h10 ;
			data[48242] <= 8'h10 ;
			data[48243] <= 8'h10 ;
			data[48244] <= 8'h10 ;
			data[48245] <= 8'h10 ;
			data[48246] <= 8'h10 ;
			data[48247] <= 8'h10 ;
			data[48248] <= 8'h10 ;
			data[48249] <= 8'h10 ;
			data[48250] <= 8'h10 ;
			data[48251] <= 8'h10 ;
			data[48252] <= 8'h10 ;
			data[48253] <= 8'h10 ;
			data[48254] <= 8'h10 ;
			data[48255] <= 8'h10 ;
			data[48256] <= 8'h10 ;
			data[48257] <= 8'h10 ;
			data[48258] <= 8'h10 ;
			data[48259] <= 8'h10 ;
			data[48260] <= 8'h10 ;
			data[48261] <= 8'h10 ;
			data[48262] <= 8'h10 ;
			data[48263] <= 8'h10 ;
			data[48264] <= 8'h10 ;
			data[48265] <= 8'h10 ;
			data[48266] <= 8'h10 ;
			data[48267] <= 8'h10 ;
			data[48268] <= 8'h10 ;
			data[48269] <= 8'h10 ;
			data[48270] <= 8'h10 ;
			data[48271] <= 8'h10 ;
			data[48272] <= 8'h10 ;
			data[48273] <= 8'h10 ;
			data[48274] <= 8'h10 ;
			data[48275] <= 8'h10 ;
			data[48276] <= 8'h10 ;
			data[48277] <= 8'h10 ;
			data[48278] <= 8'h10 ;
			data[48279] <= 8'h10 ;
			data[48280] <= 8'h10 ;
			data[48281] <= 8'h10 ;
			data[48282] <= 8'h10 ;
			data[48283] <= 8'h10 ;
			data[48284] <= 8'h10 ;
			data[48285] <= 8'h10 ;
			data[48286] <= 8'h10 ;
			data[48287] <= 8'h10 ;
			data[48288] <= 8'h10 ;
			data[48289] <= 8'h10 ;
			data[48290] <= 8'h10 ;
			data[48291] <= 8'h10 ;
			data[48292] <= 8'h10 ;
			data[48293] <= 8'h10 ;
			data[48294] <= 8'h10 ;
			data[48295] <= 8'h10 ;
			data[48296] <= 8'h10 ;
			data[48297] <= 8'h10 ;
			data[48298] <= 8'h10 ;
			data[48299] <= 8'h10 ;
			data[48300] <= 8'h10 ;
			data[48301] <= 8'h10 ;
			data[48302] <= 8'h10 ;
			data[48303] <= 8'h10 ;
			data[48304] <= 8'h10 ;
			data[48305] <= 8'h10 ;
			data[48306] <= 8'h10 ;
			data[48307] <= 8'h10 ;
			data[48308] <= 8'h10 ;
			data[48309] <= 8'h10 ;
			data[48310] <= 8'h10 ;
			data[48311] <= 8'h10 ;
			data[48312] <= 8'h10 ;
			data[48313] <= 8'h10 ;
			data[48314] <= 8'h10 ;
			data[48315] <= 8'h10 ;
			data[48316] <= 8'h10 ;
			data[48317] <= 8'h10 ;
			data[48318] <= 8'h10 ;
			data[48319] <= 8'h10 ;
			data[48320] <= 8'h10 ;
			data[48321] <= 8'h10 ;
			data[48322] <= 8'h10 ;
			data[48323] <= 8'h10 ;
			data[48324] <= 8'h10 ;
			data[48325] <= 8'h10 ;
			data[48326] <= 8'h10 ;
			data[48327] <= 8'h10 ;
			data[48328] <= 8'h10 ;
			data[48329] <= 8'h10 ;
			data[48330] <= 8'h10 ;
			data[48331] <= 8'h10 ;
			data[48332] <= 8'h10 ;
			data[48333] <= 8'h10 ;
			data[48334] <= 8'h10 ;
			data[48335] <= 8'h10 ;
			data[48336] <= 8'h10 ;
			data[48337] <= 8'h10 ;
			data[48338] <= 8'h10 ;
			data[48339] <= 8'h10 ;
			data[48340] <= 8'h10 ;
			data[48341] <= 8'h10 ;
			data[48342] <= 8'h10 ;
			data[48343] <= 8'h10 ;
			data[48344] <= 8'h10 ;
			data[48345] <= 8'h10 ;
			data[48346] <= 8'h10 ;
			data[48347] <= 8'h10 ;
			data[48348] <= 8'h10 ;
			data[48349] <= 8'h10 ;
			data[48350] <= 8'h10 ;
			data[48351] <= 8'h10 ;
			data[48352] <= 8'h10 ;
			data[48353] <= 8'h10 ;
			data[48354] <= 8'h10 ;
			data[48355] <= 8'h10 ;
			data[48356] <= 8'h10 ;
			data[48357] <= 8'h10 ;
			data[48358] <= 8'h10 ;
			data[48359] <= 8'h10 ;
			data[48360] <= 8'h10 ;
			data[48361] <= 8'h10 ;
			data[48362] <= 8'h10 ;
			data[48363] <= 8'h10 ;
			data[48364] <= 8'h10 ;
			data[48365] <= 8'h10 ;
			data[48366] <= 8'h10 ;
			data[48367] <= 8'h10 ;
			data[48368] <= 8'h10 ;
			data[48369] <= 8'h10 ;
			data[48370] <= 8'h10 ;
			data[48371] <= 8'h10 ;
			data[48372] <= 8'h10 ;
			data[48373] <= 8'h10 ;
			data[48374] <= 8'h10 ;
			data[48375] <= 8'h10 ;
			data[48376] <= 8'h10 ;
			data[48377] <= 8'h10 ;
			data[48378] <= 8'h10 ;
			data[48379] <= 8'h10 ;
			data[48380] <= 8'h10 ;
			data[48381] <= 8'h10 ;
			data[48382] <= 8'h10 ;
			data[48383] <= 8'h10 ;
			data[48384] <= 8'h10 ;
			data[48385] <= 8'h10 ;
			data[48386] <= 8'h10 ;
			data[48387] <= 8'h10 ;
			data[48388] <= 8'h10 ;
			data[48389] <= 8'h10 ;
			data[48390] <= 8'h10 ;
			data[48391] <= 8'h10 ;
			data[48392] <= 8'h10 ;
			data[48393] <= 8'h10 ;
			data[48394] <= 8'h10 ;
			data[48395] <= 8'h10 ;
			data[48396] <= 8'h10 ;
			data[48397] <= 8'h10 ;
			data[48398] <= 8'h10 ;
			data[48399] <= 8'h10 ;
			data[48400] <= 8'h10 ;
			data[48401] <= 8'h10 ;
			data[48402] <= 8'h10 ;
			data[48403] <= 8'h10 ;
			data[48404] <= 8'h10 ;
			data[48405] <= 8'h10 ;
			data[48406] <= 8'h10 ;
			data[48407] <= 8'h10 ;
			data[48408] <= 8'h10 ;
			data[48409] <= 8'h10 ;
			data[48410] <= 8'h10 ;
			data[48411] <= 8'h10 ;
			data[48412] <= 8'h10 ;
			data[48413] <= 8'h10 ;
			data[48414] <= 8'h10 ;
			data[48415] <= 8'h10 ;
			data[48416] <= 8'h10 ;
			data[48417] <= 8'h10 ;
			data[48418] <= 8'h10 ;
			data[48419] <= 8'h10 ;
			data[48420] <= 8'h10 ;
			data[48421] <= 8'h10 ;
			data[48422] <= 8'h10 ;
			data[48423] <= 8'h10 ;
			data[48424] <= 8'h10 ;
			data[48425] <= 8'h10 ;
			data[48426] <= 8'h10 ;
			data[48427] <= 8'h10 ;
			data[48428] <= 8'h10 ;
			data[48429] <= 8'h10 ;
			data[48430] <= 8'h10 ;
			data[48431] <= 8'h10 ;
			data[48432] <= 8'h10 ;
			data[48433] <= 8'h10 ;
			data[48434] <= 8'h10 ;
			data[48435] <= 8'h10 ;
			data[48436] <= 8'h10 ;
			data[48437] <= 8'h10 ;
			data[48438] <= 8'h10 ;
			data[48439] <= 8'h10 ;
			data[48440] <= 8'h10 ;
			data[48441] <= 8'h10 ;
			data[48442] <= 8'h10 ;
			data[48443] <= 8'h10 ;
			data[48444] <= 8'h10 ;
			data[48445] <= 8'h10 ;
			data[48446] <= 8'h10 ;
			data[48447] <= 8'h10 ;
			data[48448] <= 8'h10 ;
			data[48449] <= 8'h10 ;
			data[48450] <= 8'h10 ;
			data[48451] <= 8'h10 ;
			data[48452] <= 8'h10 ;
			data[48453] <= 8'h10 ;
			data[48454] <= 8'h10 ;
			data[48455] <= 8'h10 ;
			data[48456] <= 8'h10 ;
			data[48457] <= 8'h10 ;
			data[48458] <= 8'h10 ;
			data[48459] <= 8'h10 ;
			data[48460] <= 8'h10 ;
			data[48461] <= 8'h10 ;
			data[48462] <= 8'h10 ;
			data[48463] <= 8'h10 ;
			data[48464] <= 8'h10 ;
			data[48465] <= 8'h10 ;
			data[48466] <= 8'h10 ;
			data[48467] <= 8'h10 ;
			data[48468] <= 8'h10 ;
			data[48469] <= 8'h10 ;
			data[48470] <= 8'h10 ;
			data[48471] <= 8'h10 ;
			data[48472] <= 8'h10 ;
			data[48473] <= 8'h10 ;
			data[48474] <= 8'h10 ;
			data[48475] <= 8'h10 ;
			data[48476] <= 8'h10 ;
			data[48477] <= 8'h10 ;
			data[48478] <= 8'h10 ;
			data[48479] <= 8'h10 ;
			data[48480] <= 8'h10 ;
			data[48481] <= 8'h10 ;
			data[48482] <= 8'h10 ;
			data[48483] <= 8'h10 ;
			data[48484] <= 8'h10 ;
			data[48485] <= 8'h10 ;
			data[48486] <= 8'h10 ;
			data[48487] <= 8'h10 ;
			data[48488] <= 8'h10 ;
			data[48489] <= 8'h10 ;
			data[48490] <= 8'h10 ;
			data[48491] <= 8'h10 ;
			data[48492] <= 8'h10 ;
			data[48493] <= 8'h10 ;
			data[48494] <= 8'h10 ;
			data[48495] <= 8'h10 ;
			data[48496] <= 8'h10 ;
			data[48497] <= 8'h10 ;
			data[48498] <= 8'h10 ;
			data[48499] <= 8'h10 ;
			data[48500] <= 8'h10 ;
			data[48501] <= 8'h10 ;
			data[48502] <= 8'h10 ;
			data[48503] <= 8'h10 ;
			data[48504] <= 8'h10 ;
			data[48505] <= 8'h10 ;
			data[48506] <= 8'h10 ;
			data[48507] <= 8'h10 ;
			data[48508] <= 8'h10 ;
			data[48509] <= 8'h10 ;
			data[48510] <= 8'h10 ;
			data[48511] <= 8'h10 ;
			data[48512] <= 8'h10 ;
			data[48513] <= 8'h10 ;
			data[48514] <= 8'h10 ;
			data[48515] <= 8'h10 ;
			data[48516] <= 8'h10 ;
			data[48517] <= 8'h10 ;
			data[48518] <= 8'h10 ;
			data[48519] <= 8'h10 ;
			data[48520] <= 8'h10 ;
			data[48521] <= 8'h10 ;
			data[48522] <= 8'h10 ;
			data[48523] <= 8'h10 ;
			data[48524] <= 8'h10 ;
			data[48525] <= 8'h10 ;
			data[48526] <= 8'h10 ;
			data[48527] <= 8'h10 ;
			data[48528] <= 8'h10 ;
			data[48529] <= 8'h10 ;
			data[48530] <= 8'h10 ;
			data[48531] <= 8'h10 ;
			data[48532] <= 8'h10 ;
			data[48533] <= 8'h10 ;
			data[48534] <= 8'h10 ;
			data[48535] <= 8'h10 ;
			data[48536] <= 8'h10 ;
			data[48537] <= 8'h10 ;
			data[48538] <= 8'h10 ;
			data[48539] <= 8'h10 ;
			data[48540] <= 8'h10 ;
			data[48541] <= 8'h10 ;
			data[48542] <= 8'h10 ;
			data[48543] <= 8'h10 ;
			data[48544] <= 8'h10 ;
			data[48545] <= 8'h10 ;
			data[48546] <= 8'h10 ;
			data[48547] <= 8'h10 ;
			data[48548] <= 8'h10 ;
			data[48549] <= 8'h10 ;
			data[48550] <= 8'h10 ;
			data[48551] <= 8'h10 ;
			data[48552] <= 8'h10 ;
			data[48553] <= 8'h10 ;
			data[48554] <= 8'h10 ;
			data[48555] <= 8'h10 ;
			data[48556] <= 8'h10 ;
			data[48557] <= 8'h10 ;
			data[48558] <= 8'h10 ;
			data[48559] <= 8'h10 ;
			data[48560] <= 8'h10 ;
			data[48561] <= 8'h10 ;
			data[48562] <= 8'h10 ;
			data[48563] <= 8'h10 ;
			data[48564] <= 8'h10 ;
			data[48565] <= 8'h10 ;
			data[48566] <= 8'h10 ;
			data[48567] <= 8'h10 ;
			data[48568] <= 8'h10 ;
			data[48569] <= 8'h10 ;
			data[48570] <= 8'h10 ;
			data[48571] <= 8'h10 ;
			data[48572] <= 8'h10 ;
			data[48573] <= 8'h10 ;
			data[48574] <= 8'h10 ;
			data[48575] <= 8'h10 ;
			data[48576] <= 8'h10 ;
			data[48577] <= 8'h10 ;
			data[48578] <= 8'h10 ;
			data[48579] <= 8'h10 ;
			data[48580] <= 8'h10 ;
			data[48581] <= 8'h10 ;
			data[48582] <= 8'h10 ;
			data[48583] <= 8'h10 ;
			data[48584] <= 8'h10 ;
			data[48585] <= 8'h10 ;
			data[48586] <= 8'h10 ;
			data[48587] <= 8'h10 ;
			data[48588] <= 8'h10 ;
			data[48589] <= 8'h10 ;
			data[48590] <= 8'h10 ;
			data[48591] <= 8'h10 ;
			data[48592] <= 8'h10 ;
			data[48593] <= 8'h10 ;
			data[48594] <= 8'h10 ;
			data[48595] <= 8'h10 ;
			data[48596] <= 8'h10 ;
			data[48597] <= 8'h10 ;
			data[48598] <= 8'h10 ;
			data[48599] <= 8'h10 ;
			data[48600] <= 8'h10 ;
			data[48601] <= 8'h10 ;
			data[48602] <= 8'h10 ;
			data[48603] <= 8'h10 ;
			data[48604] <= 8'h10 ;
			data[48605] <= 8'h10 ;
			data[48606] <= 8'h10 ;
			data[48607] <= 8'h10 ;
			data[48608] <= 8'h10 ;
			data[48609] <= 8'h10 ;
			data[48610] <= 8'h10 ;
			data[48611] <= 8'h10 ;
			data[48612] <= 8'h10 ;
			data[48613] <= 8'h10 ;
			data[48614] <= 8'h10 ;
			data[48615] <= 8'h10 ;
			data[48616] <= 8'h10 ;
			data[48617] <= 8'h10 ;
			data[48618] <= 8'h10 ;
			data[48619] <= 8'h10 ;
			data[48620] <= 8'h10 ;
			data[48621] <= 8'h10 ;
			data[48622] <= 8'h10 ;
			data[48623] <= 8'h10 ;
			data[48624] <= 8'h10 ;
			data[48625] <= 8'h10 ;
			data[48626] <= 8'h10 ;
			data[48627] <= 8'h10 ;
			data[48628] <= 8'h10 ;
			data[48629] <= 8'h10 ;
			data[48630] <= 8'h10 ;
			data[48631] <= 8'h10 ;
			data[48632] <= 8'h10 ;
			data[48633] <= 8'h10 ;
			data[48634] <= 8'h10 ;
			data[48635] <= 8'h10 ;
			data[48636] <= 8'h10 ;
			data[48637] <= 8'h10 ;
			data[48638] <= 8'h10 ;
			data[48639] <= 8'h10 ;
			data[48640] <= 8'h10 ;
			data[48641] <= 8'h10 ;
			data[48642] <= 8'h10 ;
			data[48643] <= 8'h10 ;
			data[48644] <= 8'h10 ;
			data[48645] <= 8'h10 ;
			data[48646] <= 8'h10 ;
			data[48647] <= 8'h10 ;
			data[48648] <= 8'h10 ;
			data[48649] <= 8'h10 ;
			data[48650] <= 8'h10 ;
			data[48651] <= 8'h10 ;
			data[48652] <= 8'h10 ;
			data[48653] <= 8'h10 ;
			data[48654] <= 8'h10 ;
			data[48655] <= 8'h10 ;
			data[48656] <= 8'h10 ;
			data[48657] <= 8'h10 ;
			data[48658] <= 8'h10 ;
			data[48659] <= 8'h10 ;
			data[48660] <= 8'h10 ;
			data[48661] <= 8'h10 ;
			data[48662] <= 8'h10 ;
			data[48663] <= 8'h10 ;
			data[48664] <= 8'h10 ;
			data[48665] <= 8'h10 ;
			data[48666] <= 8'h10 ;
			data[48667] <= 8'h10 ;
			data[48668] <= 8'h10 ;
			data[48669] <= 8'h10 ;
			data[48670] <= 8'h10 ;
			data[48671] <= 8'h10 ;
			data[48672] <= 8'h10 ;
			data[48673] <= 8'h10 ;
			data[48674] <= 8'h10 ;
			data[48675] <= 8'h10 ;
			data[48676] <= 8'h10 ;
			data[48677] <= 8'h10 ;
			data[48678] <= 8'h10 ;
			data[48679] <= 8'h10 ;
			data[48680] <= 8'h10 ;
			data[48681] <= 8'h10 ;
			data[48682] <= 8'h10 ;
			data[48683] <= 8'h10 ;
			data[48684] <= 8'h10 ;
			data[48685] <= 8'h10 ;
			data[48686] <= 8'h10 ;
			data[48687] <= 8'h10 ;
			data[48688] <= 8'h10 ;
			data[48689] <= 8'h10 ;
			data[48690] <= 8'h10 ;
			data[48691] <= 8'h10 ;
			data[48692] <= 8'h10 ;
			data[48693] <= 8'h10 ;
			data[48694] <= 8'h10 ;
			data[48695] <= 8'h10 ;
			data[48696] <= 8'h10 ;
			data[48697] <= 8'h10 ;
			data[48698] <= 8'h10 ;
			data[48699] <= 8'h10 ;
			data[48700] <= 8'h10 ;
			data[48701] <= 8'h10 ;
			data[48702] <= 8'h10 ;
			data[48703] <= 8'h10 ;
			data[48704] <= 8'h10 ;
			data[48705] <= 8'h10 ;
			data[48706] <= 8'h10 ;
			data[48707] <= 8'h10 ;
			data[48708] <= 8'h10 ;
			data[48709] <= 8'h10 ;
			data[48710] <= 8'h10 ;
			data[48711] <= 8'h10 ;
			data[48712] <= 8'h10 ;
			data[48713] <= 8'h10 ;
			data[48714] <= 8'h10 ;
			data[48715] <= 8'h10 ;
			data[48716] <= 8'h10 ;
			data[48717] <= 8'h10 ;
			data[48718] <= 8'h10 ;
			data[48719] <= 8'h10 ;
			data[48720] <= 8'h10 ;
			data[48721] <= 8'h10 ;
			data[48722] <= 8'h10 ;
			data[48723] <= 8'h10 ;
			data[48724] <= 8'h10 ;
			data[48725] <= 8'h10 ;
			data[48726] <= 8'h10 ;
			data[48727] <= 8'h10 ;
			data[48728] <= 8'h10 ;
			data[48729] <= 8'h10 ;
			data[48730] <= 8'h10 ;
			data[48731] <= 8'h10 ;
			data[48732] <= 8'h10 ;
			data[48733] <= 8'h10 ;
			data[48734] <= 8'h10 ;
			data[48735] <= 8'h10 ;
			data[48736] <= 8'h10 ;
			data[48737] <= 8'h10 ;
			data[48738] <= 8'h10 ;
			data[48739] <= 8'h10 ;
			data[48740] <= 8'h10 ;
			data[48741] <= 8'h10 ;
			data[48742] <= 8'h10 ;
			data[48743] <= 8'h10 ;
			data[48744] <= 8'h10 ;
			data[48745] <= 8'h10 ;
			data[48746] <= 8'h10 ;
			data[48747] <= 8'h10 ;
			data[48748] <= 8'h10 ;
			data[48749] <= 8'h10 ;
			data[48750] <= 8'h10 ;
			data[48751] <= 8'h10 ;
			data[48752] <= 8'h10 ;
			data[48753] <= 8'h10 ;
			data[48754] <= 8'h10 ;
			data[48755] <= 8'h10 ;
			data[48756] <= 8'h10 ;
			data[48757] <= 8'h10 ;
			data[48758] <= 8'h10 ;
			data[48759] <= 8'h10 ;
			data[48760] <= 8'h10 ;
			data[48761] <= 8'h10 ;
			data[48762] <= 8'h10 ;
			data[48763] <= 8'h10 ;
			data[48764] <= 8'h10 ;
			data[48765] <= 8'h10 ;
			data[48766] <= 8'h10 ;
			data[48767] <= 8'h10 ;
			data[48768] <= 8'h10 ;
			data[48769] <= 8'h10 ;
			data[48770] <= 8'h10 ;
			data[48771] <= 8'h10 ;
			data[48772] <= 8'h10 ;
			data[48773] <= 8'h10 ;
			data[48774] <= 8'h10 ;
			data[48775] <= 8'h10 ;
			data[48776] <= 8'h10 ;
			data[48777] <= 8'h10 ;
			data[48778] <= 8'h10 ;
			data[48779] <= 8'h10 ;
			data[48780] <= 8'h10 ;
			data[48781] <= 8'h10 ;
			data[48782] <= 8'h10 ;
			data[48783] <= 8'h10 ;
			data[48784] <= 8'h10 ;
			data[48785] <= 8'h10 ;
			data[48786] <= 8'h10 ;
			data[48787] <= 8'h10 ;
			data[48788] <= 8'h10 ;
			data[48789] <= 8'h10 ;
			data[48790] <= 8'h10 ;
			data[48791] <= 8'h10 ;
			data[48792] <= 8'h10 ;
			data[48793] <= 8'h10 ;
			data[48794] <= 8'h10 ;
			data[48795] <= 8'h10 ;
			data[48796] <= 8'h10 ;
			data[48797] <= 8'h10 ;
			data[48798] <= 8'h10 ;
			data[48799] <= 8'h10 ;
			data[48800] <= 8'h10 ;
			data[48801] <= 8'h10 ;
			data[48802] <= 8'h10 ;
			data[48803] <= 8'h10 ;
			data[48804] <= 8'h10 ;
			data[48805] <= 8'h10 ;
			data[48806] <= 8'h10 ;
			data[48807] <= 8'h10 ;
			data[48808] <= 8'h10 ;
			data[48809] <= 8'h10 ;
			data[48810] <= 8'h10 ;
			data[48811] <= 8'h10 ;
			data[48812] <= 8'h10 ;
			data[48813] <= 8'h10 ;
			data[48814] <= 8'h10 ;
			data[48815] <= 8'h10 ;
			data[48816] <= 8'h10 ;
			data[48817] <= 8'h10 ;
			data[48818] <= 8'h10 ;
			data[48819] <= 8'h10 ;
			data[48820] <= 8'h10 ;
			data[48821] <= 8'h10 ;
			data[48822] <= 8'h10 ;
			data[48823] <= 8'h10 ;
			data[48824] <= 8'h10 ;
			data[48825] <= 8'h10 ;
			data[48826] <= 8'h10 ;
			data[48827] <= 8'h10 ;
			data[48828] <= 8'h10 ;
			data[48829] <= 8'h10 ;
			data[48830] <= 8'h10 ;
			data[48831] <= 8'h10 ;
			data[48832] <= 8'h10 ;
			data[48833] <= 8'h10 ;
			data[48834] <= 8'h10 ;
			data[48835] <= 8'h10 ;
			data[48836] <= 8'h10 ;
			data[48837] <= 8'h10 ;
			data[48838] <= 8'h10 ;
			data[48839] <= 8'h10 ;
			data[48840] <= 8'h10 ;
			data[48841] <= 8'h10 ;
			data[48842] <= 8'h10 ;
			data[48843] <= 8'h10 ;
			data[48844] <= 8'h10 ;
			data[48845] <= 8'h10 ;
			data[48846] <= 8'h10 ;
			data[48847] <= 8'h10 ;
			data[48848] <= 8'h10 ;
			data[48849] <= 8'h10 ;
			data[48850] <= 8'h10 ;
			data[48851] <= 8'h10 ;
			data[48852] <= 8'h10 ;
			data[48853] <= 8'h10 ;
			data[48854] <= 8'h10 ;
			data[48855] <= 8'h10 ;
			data[48856] <= 8'h10 ;
			data[48857] <= 8'h10 ;
			data[48858] <= 8'h10 ;
			data[48859] <= 8'h10 ;
			data[48860] <= 8'h10 ;
			data[48861] <= 8'h10 ;
			data[48862] <= 8'h10 ;
			data[48863] <= 8'h10 ;
			data[48864] <= 8'h10 ;
			data[48865] <= 8'h10 ;
			data[48866] <= 8'h10 ;
			data[48867] <= 8'h10 ;
			data[48868] <= 8'h10 ;
			data[48869] <= 8'h10 ;
			data[48870] <= 8'h10 ;
			data[48871] <= 8'h10 ;
			data[48872] <= 8'h10 ;
			data[48873] <= 8'h10 ;
			data[48874] <= 8'h10 ;
			data[48875] <= 8'h10 ;
			data[48876] <= 8'h10 ;
			data[48877] <= 8'h10 ;
			data[48878] <= 8'h10 ;
			data[48879] <= 8'h10 ;
			data[48880] <= 8'h10 ;
			data[48881] <= 8'h10 ;
			data[48882] <= 8'h10 ;
			data[48883] <= 8'h10 ;
			data[48884] <= 8'h10 ;
			data[48885] <= 8'h10 ;
			data[48886] <= 8'h10 ;
			data[48887] <= 8'h10 ;
			data[48888] <= 8'h10 ;
			data[48889] <= 8'h10 ;
			data[48890] <= 8'h10 ;
			data[48891] <= 8'h10 ;
			data[48892] <= 8'h10 ;
			data[48893] <= 8'h10 ;
			data[48894] <= 8'h10 ;
			data[48895] <= 8'h10 ;
			data[48896] <= 8'h10 ;
			data[48897] <= 8'h10 ;
			data[48898] <= 8'h10 ;
			data[48899] <= 8'h10 ;
			data[48900] <= 8'h10 ;
			data[48901] <= 8'h10 ;
			data[48902] <= 8'h10 ;
			data[48903] <= 8'h10 ;
			data[48904] <= 8'h10 ;
			data[48905] <= 8'h10 ;
			data[48906] <= 8'h10 ;
			data[48907] <= 8'h10 ;
			data[48908] <= 8'h10 ;
			data[48909] <= 8'h10 ;
			data[48910] <= 8'h10 ;
			data[48911] <= 8'h10 ;
			data[48912] <= 8'h10 ;
			data[48913] <= 8'h10 ;
			data[48914] <= 8'h10 ;
			data[48915] <= 8'h10 ;
			data[48916] <= 8'h10 ;
			data[48917] <= 8'h10 ;
			data[48918] <= 8'h10 ;
			data[48919] <= 8'h10 ;
			data[48920] <= 8'h10 ;
			data[48921] <= 8'h10 ;
			data[48922] <= 8'h10 ;
			data[48923] <= 8'h10 ;
			data[48924] <= 8'h10 ;
			data[48925] <= 8'h10 ;
			data[48926] <= 8'h10 ;
			data[48927] <= 8'h10 ;
			data[48928] <= 8'h10 ;
			data[48929] <= 8'h10 ;
			data[48930] <= 8'h10 ;
			data[48931] <= 8'h10 ;
			data[48932] <= 8'h10 ;
			data[48933] <= 8'h10 ;
			data[48934] <= 8'h10 ;
			data[48935] <= 8'h10 ;
			data[48936] <= 8'h10 ;
			data[48937] <= 8'h10 ;
			data[48938] <= 8'h10 ;
			data[48939] <= 8'h10 ;
			data[48940] <= 8'h10 ;
			data[48941] <= 8'h10 ;
			data[48942] <= 8'h10 ;
			data[48943] <= 8'h10 ;
			data[48944] <= 8'h10 ;
			data[48945] <= 8'h10 ;
			data[48946] <= 8'h10 ;
			data[48947] <= 8'h10 ;
			data[48948] <= 8'h10 ;
			data[48949] <= 8'h10 ;
			data[48950] <= 8'h10 ;
			data[48951] <= 8'h10 ;
			data[48952] <= 8'h10 ;
			data[48953] <= 8'h10 ;
			data[48954] <= 8'h10 ;
			data[48955] <= 8'h10 ;
			data[48956] <= 8'h10 ;
			data[48957] <= 8'h10 ;
			data[48958] <= 8'h10 ;
			data[48959] <= 8'h10 ;
			data[48960] <= 8'h10 ;
			data[48961] <= 8'h10 ;
			data[48962] <= 8'h10 ;
			data[48963] <= 8'h10 ;
			data[48964] <= 8'h10 ;
			data[48965] <= 8'h10 ;
			data[48966] <= 8'h10 ;
			data[48967] <= 8'h10 ;
			data[48968] <= 8'h10 ;
			data[48969] <= 8'h10 ;
			data[48970] <= 8'h10 ;
			data[48971] <= 8'h10 ;
			data[48972] <= 8'h10 ;
			data[48973] <= 8'h10 ;
			data[48974] <= 8'h10 ;
			data[48975] <= 8'h10 ;
			data[48976] <= 8'h10 ;
			data[48977] <= 8'h10 ;
			data[48978] <= 8'h10 ;
			data[48979] <= 8'h10 ;
			data[48980] <= 8'h10 ;
			data[48981] <= 8'h10 ;
			data[48982] <= 8'h10 ;
			data[48983] <= 8'h10 ;
			data[48984] <= 8'h10 ;
			data[48985] <= 8'h10 ;
			data[48986] <= 8'h10 ;
			data[48987] <= 8'h10 ;
			data[48988] <= 8'h10 ;
			data[48989] <= 8'h10 ;
			data[48990] <= 8'h10 ;
			data[48991] <= 8'h10 ;
			data[48992] <= 8'h10 ;
			data[48993] <= 8'h10 ;
			data[48994] <= 8'h10 ;
			data[48995] <= 8'h10 ;
			data[48996] <= 8'h10 ;
			data[48997] <= 8'h10 ;
			data[48998] <= 8'h10 ;
			data[48999] <= 8'h10 ;
			data[49000] <= 8'h10 ;
			data[49001] <= 8'h10 ;
			data[49002] <= 8'h10 ;
			data[49003] <= 8'h10 ;
			data[49004] <= 8'h10 ;
			data[49005] <= 8'h10 ;
			data[49006] <= 8'h10 ;
			data[49007] <= 8'h10 ;
			data[49008] <= 8'h10 ;
			data[49009] <= 8'h10 ;
			data[49010] <= 8'h10 ;
			data[49011] <= 8'h10 ;
			data[49012] <= 8'h10 ;
			data[49013] <= 8'h10 ;
			data[49014] <= 8'h10 ;
			data[49015] <= 8'h10 ;
			data[49016] <= 8'h10 ;
			data[49017] <= 8'h10 ;
			data[49018] <= 8'h10 ;
			data[49019] <= 8'h10 ;
			data[49020] <= 8'h10 ;
			data[49021] <= 8'h10 ;
			data[49022] <= 8'h10 ;
			data[49023] <= 8'h10 ;
			data[49024] <= 8'h10 ;
			data[49025] <= 8'h10 ;
			data[49026] <= 8'h10 ;
			data[49027] <= 8'h10 ;
			data[49028] <= 8'h10 ;
			data[49029] <= 8'h10 ;
			data[49030] <= 8'h10 ;
			data[49031] <= 8'h10 ;
			data[49032] <= 8'h10 ;
			data[49033] <= 8'h10 ;
			data[49034] <= 8'h10 ;
			data[49035] <= 8'h10 ;
			data[49036] <= 8'h10 ;
			data[49037] <= 8'h10 ;
			data[49038] <= 8'h10 ;
			data[49039] <= 8'h10 ;
			data[49040] <= 8'h10 ;
			data[49041] <= 8'h10 ;
			data[49042] <= 8'h10 ;
			data[49043] <= 8'h10 ;
			data[49044] <= 8'h10 ;
			data[49045] <= 8'h10 ;
			data[49046] <= 8'h10 ;
			data[49047] <= 8'h10 ;
			data[49048] <= 8'h10 ;
			data[49049] <= 8'h10 ;
			data[49050] <= 8'h10 ;
			data[49051] <= 8'h10 ;
			data[49052] <= 8'h10 ;
			data[49053] <= 8'h10 ;
			data[49054] <= 8'h10 ;
			data[49055] <= 8'h10 ;
			data[49056] <= 8'h10 ;
			data[49057] <= 8'h10 ;
			data[49058] <= 8'h10 ;
			data[49059] <= 8'h10 ;
			data[49060] <= 8'h10 ;
			data[49061] <= 8'h10 ;
			data[49062] <= 8'h10 ;
			data[49063] <= 8'h10 ;
			data[49064] <= 8'h10 ;
			data[49065] <= 8'h10 ;
			data[49066] <= 8'h10 ;
			data[49067] <= 8'h10 ;
			data[49068] <= 8'h10 ;
			data[49069] <= 8'h10 ;
			data[49070] <= 8'h10 ;
			data[49071] <= 8'h10 ;
			data[49072] <= 8'h10 ;
			data[49073] <= 8'h10 ;
			data[49074] <= 8'h10 ;
			data[49075] <= 8'h10 ;
			data[49076] <= 8'h10 ;
			data[49077] <= 8'h10 ;
			data[49078] <= 8'h10 ;
			data[49079] <= 8'h10 ;
			data[49080] <= 8'h10 ;
			data[49081] <= 8'h10 ;
			data[49082] <= 8'h10 ;
			data[49083] <= 8'h10 ;
			data[49084] <= 8'h10 ;
			data[49085] <= 8'h10 ;
			data[49086] <= 8'h10 ;
			data[49087] <= 8'h10 ;
			data[49088] <= 8'h10 ;
			data[49089] <= 8'h10 ;
			data[49090] <= 8'h10 ;
			data[49091] <= 8'h10 ;
			data[49092] <= 8'h10 ;
			data[49093] <= 8'h10 ;
			data[49094] <= 8'h10 ;
			data[49095] <= 8'h10 ;
			data[49096] <= 8'h10 ;
			data[49097] <= 8'h10 ;
			data[49098] <= 8'h10 ;
			data[49099] <= 8'h10 ;
			data[49100] <= 8'h10 ;
			data[49101] <= 8'h10 ;
			data[49102] <= 8'h10 ;
			data[49103] <= 8'h10 ;
			data[49104] <= 8'h10 ;
			data[49105] <= 8'h10 ;
			data[49106] <= 8'h10 ;
			data[49107] <= 8'h10 ;
			data[49108] <= 8'h10 ;
			data[49109] <= 8'h10 ;
			data[49110] <= 8'h10 ;
			data[49111] <= 8'h10 ;
			data[49112] <= 8'h10 ;
			data[49113] <= 8'h10 ;
			data[49114] <= 8'h10 ;
			data[49115] <= 8'h10 ;
			data[49116] <= 8'h10 ;
			data[49117] <= 8'h10 ;
			data[49118] <= 8'h10 ;
			data[49119] <= 8'h10 ;
			data[49120] <= 8'h10 ;
			data[49121] <= 8'h10 ;
			data[49122] <= 8'h10 ;
			data[49123] <= 8'h10 ;
			data[49124] <= 8'h10 ;
			data[49125] <= 8'h10 ;
			data[49126] <= 8'h10 ;
			data[49127] <= 8'h10 ;
			data[49128] <= 8'h10 ;
			data[49129] <= 8'h10 ;
			data[49130] <= 8'h10 ;
			data[49131] <= 8'h10 ;
			data[49132] <= 8'h10 ;
			data[49133] <= 8'h10 ;
			data[49134] <= 8'h10 ;
			data[49135] <= 8'h10 ;
			data[49136] <= 8'h10 ;
			data[49137] <= 8'h10 ;
			data[49138] <= 8'h10 ;
			data[49139] <= 8'h10 ;
			data[49140] <= 8'h10 ;
			data[49141] <= 8'h10 ;
			data[49142] <= 8'h10 ;
			data[49143] <= 8'h10 ;
			data[49144] <= 8'h10 ;
			data[49145] <= 8'h10 ;
			data[49146] <= 8'h10 ;
			data[49147] <= 8'h10 ;
			data[49148] <= 8'h10 ;
			data[49149] <= 8'h10 ;
			data[49150] <= 8'h10 ;
			data[49151] <= 8'h10 ;
			data[49152] <= 8'h10 ;
			data[49153] <= 8'h10 ;
			data[49154] <= 8'h10 ;
			data[49155] <= 8'h10 ;
			data[49156] <= 8'h10 ;
			data[49157] <= 8'h10 ;
			data[49158] <= 8'h10 ;
			data[49159] <= 8'h10 ;
			data[49160] <= 8'h10 ;
			data[49161] <= 8'h10 ;
			data[49162] <= 8'h10 ;
			data[49163] <= 8'h10 ;
			data[49164] <= 8'h10 ;
			data[49165] <= 8'h10 ;
			data[49166] <= 8'h10 ;
			data[49167] <= 8'h10 ;
			data[49168] <= 8'h10 ;
			data[49169] <= 8'h10 ;
			data[49170] <= 8'h10 ;
			data[49171] <= 8'h10 ;
			data[49172] <= 8'h10 ;
			data[49173] <= 8'h10 ;
			data[49174] <= 8'h10 ;
			data[49175] <= 8'h10 ;
			data[49176] <= 8'h10 ;
			data[49177] <= 8'h10 ;
			data[49178] <= 8'h10 ;
			data[49179] <= 8'h10 ;
			data[49180] <= 8'h10 ;
			data[49181] <= 8'h10 ;
			data[49182] <= 8'h10 ;
			data[49183] <= 8'h10 ;
			data[49184] <= 8'h10 ;
			data[49185] <= 8'h10 ;
			data[49186] <= 8'h10 ;
			data[49187] <= 8'h10 ;
			data[49188] <= 8'h10 ;
			data[49189] <= 8'h10 ;
			data[49190] <= 8'h10 ;
			data[49191] <= 8'h10 ;
			data[49192] <= 8'h10 ;
			data[49193] <= 8'h10 ;
			data[49194] <= 8'h10 ;
			data[49195] <= 8'h10 ;
			data[49196] <= 8'h10 ;
			data[49197] <= 8'h10 ;
			data[49198] <= 8'h10 ;
			data[49199] <= 8'h10 ;
			data[49200] <= 8'h10 ;
			data[49201] <= 8'h10 ;
			data[49202] <= 8'h10 ;
			data[49203] <= 8'h10 ;
			data[49204] <= 8'h10 ;
			data[49205] <= 8'h10 ;
			data[49206] <= 8'h10 ;
			data[49207] <= 8'h10 ;
			data[49208] <= 8'h10 ;
			data[49209] <= 8'h10 ;
			data[49210] <= 8'h10 ;
			data[49211] <= 8'h10 ;
			data[49212] <= 8'h10 ;
			data[49213] <= 8'h10 ;
			data[49214] <= 8'h10 ;
			data[49215] <= 8'h10 ;
			data[49216] <= 8'h10 ;
			data[49217] <= 8'h10 ;
			data[49218] <= 8'h10 ;
			data[49219] <= 8'h10 ;
			data[49220] <= 8'h10 ;
			data[49221] <= 8'h10 ;
			data[49222] <= 8'h10 ;
			data[49223] <= 8'h10 ;
			data[49224] <= 8'h10 ;
			data[49225] <= 8'h10 ;
			data[49226] <= 8'h10 ;
			data[49227] <= 8'h10 ;
			data[49228] <= 8'h10 ;
			data[49229] <= 8'h10 ;
			data[49230] <= 8'h10 ;
			data[49231] <= 8'h10 ;
			data[49232] <= 8'h10 ;
			data[49233] <= 8'h10 ;
			data[49234] <= 8'h10 ;
			data[49235] <= 8'h10 ;
			data[49236] <= 8'h10 ;
			data[49237] <= 8'h10 ;
			data[49238] <= 8'h10 ;
			data[49239] <= 8'h10 ;
			data[49240] <= 8'h10 ;
			data[49241] <= 8'h10 ;
			data[49242] <= 8'h10 ;
			data[49243] <= 8'h10 ;
			data[49244] <= 8'h10 ;
			data[49245] <= 8'h10 ;
			data[49246] <= 8'h10 ;
			data[49247] <= 8'h10 ;
			data[49248] <= 8'h10 ;
			data[49249] <= 8'h10 ;
			data[49250] <= 8'h10 ;
			data[49251] <= 8'h10 ;
			data[49252] <= 8'h10 ;
			data[49253] <= 8'h10 ;
			data[49254] <= 8'h10 ;
			data[49255] <= 8'h10 ;
			data[49256] <= 8'h10 ;
			data[49257] <= 8'h10 ;
			data[49258] <= 8'h10 ;
			data[49259] <= 8'h10 ;
			data[49260] <= 8'h10 ;
			data[49261] <= 8'h10 ;
			data[49262] <= 8'h10 ;
			data[49263] <= 8'h10 ;
			data[49264] <= 8'h10 ;
			data[49265] <= 8'h10 ;
			data[49266] <= 8'h10 ;
			data[49267] <= 8'h10 ;
			data[49268] <= 8'h10 ;
			data[49269] <= 8'h10 ;
			data[49270] <= 8'h10 ;
			data[49271] <= 8'h10 ;
			data[49272] <= 8'h10 ;
			data[49273] <= 8'h10 ;
			data[49274] <= 8'h10 ;
			data[49275] <= 8'h10 ;
			data[49276] <= 8'h10 ;
			data[49277] <= 8'h10 ;
			data[49278] <= 8'h10 ;
			data[49279] <= 8'h10 ;
			data[49280] <= 8'h10 ;
			data[49281] <= 8'h10 ;
			data[49282] <= 8'h10 ;
			data[49283] <= 8'h10 ;
			data[49284] <= 8'h10 ;
			data[49285] <= 8'h10 ;
			data[49286] <= 8'h10 ;
			data[49287] <= 8'h10 ;
			data[49288] <= 8'h10 ;
			data[49289] <= 8'h10 ;
			data[49290] <= 8'h10 ;
			data[49291] <= 8'h10 ;
			data[49292] <= 8'h10 ;
			data[49293] <= 8'h10 ;
			data[49294] <= 8'h10 ;
			data[49295] <= 8'h10 ;
			data[49296] <= 8'h10 ;
			data[49297] <= 8'h10 ;
			data[49298] <= 8'h10 ;
			data[49299] <= 8'h10 ;
			data[49300] <= 8'h10 ;
			data[49301] <= 8'h10 ;
			data[49302] <= 8'h10 ;
			data[49303] <= 8'h10 ;
			data[49304] <= 8'h10 ;
			data[49305] <= 8'h10 ;
			data[49306] <= 8'h10 ;
			data[49307] <= 8'h10 ;
			data[49308] <= 8'h10 ;
			data[49309] <= 8'h10 ;
			data[49310] <= 8'h10 ;
			data[49311] <= 8'h10 ;
			data[49312] <= 8'h10 ;
			data[49313] <= 8'h10 ;
			data[49314] <= 8'h10 ;
			data[49315] <= 8'h10 ;
			data[49316] <= 8'h10 ;
			data[49317] <= 8'h10 ;
			data[49318] <= 8'h10 ;
			data[49319] <= 8'h10 ;
			data[49320] <= 8'h10 ;
			data[49321] <= 8'h10 ;
			data[49322] <= 8'h10 ;
			data[49323] <= 8'h10 ;
			data[49324] <= 8'h10 ;
			data[49325] <= 8'h10 ;
			data[49326] <= 8'h10 ;
			data[49327] <= 8'h10 ;
			data[49328] <= 8'h10 ;
			data[49329] <= 8'h10 ;
			data[49330] <= 8'h10 ;
			data[49331] <= 8'h10 ;
			data[49332] <= 8'h10 ;
			data[49333] <= 8'h10 ;
			data[49334] <= 8'h10 ;
			data[49335] <= 8'h10 ;
			data[49336] <= 8'h10 ;
			data[49337] <= 8'h10 ;
			data[49338] <= 8'h10 ;
			data[49339] <= 8'h10 ;
			data[49340] <= 8'h10 ;
			data[49341] <= 8'h10 ;
			data[49342] <= 8'h10 ;
			data[49343] <= 8'h10 ;
			data[49344] <= 8'h10 ;
			data[49345] <= 8'h10 ;
			data[49346] <= 8'h10 ;
			data[49347] <= 8'h10 ;
			data[49348] <= 8'h10 ;
			data[49349] <= 8'h10 ;
			data[49350] <= 8'h10 ;
			data[49351] <= 8'h10 ;
			data[49352] <= 8'h10 ;
			data[49353] <= 8'h10 ;
			data[49354] <= 8'h10 ;
			data[49355] <= 8'h10 ;
			data[49356] <= 8'h10 ;
			data[49357] <= 8'h10 ;
			data[49358] <= 8'h10 ;
			data[49359] <= 8'h10 ;
			data[49360] <= 8'h10 ;
			data[49361] <= 8'h10 ;
			data[49362] <= 8'h10 ;
			data[49363] <= 8'h10 ;
			data[49364] <= 8'h10 ;
			data[49365] <= 8'h10 ;
			data[49366] <= 8'h10 ;
			data[49367] <= 8'h10 ;
			data[49368] <= 8'h10 ;
			data[49369] <= 8'h10 ;
			data[49370] <= 8'h10 ;
			data[49371] <= 8'h10 ;
			data[49372] <= 8'h10 ;
			data[49373] <= 8'h10 ;
			data[49374] <= 8'h10 ;
			data[49375] <= 8'h10 ;
			data[49376] <= 8'h10 ;
			data[49377] <= 8'h10 ;
			data[49378] <= 8'h10 ;
			data[49379] <= 8'h10 ;
			data[49380] <= 8'h10 ;
			data[49381] <= 8'h10 ;
			data[49382] <= 8'h10 ;
			data[49383] <= 8'h10 ;
			data[49384] <= 8'h10 ;
			data[49385] <= 8'h10 ;
			data[49386] <= 8'h10 ;
			data[49387] <= 8'h10 ;
			data[49388] <= 8'h10 ;
			data[49389] <= 8'h10 ;
			data[49390] <= 8'h10 ;
			data[49391] <= 8'h10 ;
			data[49392] <= 8'h10 ;
			data[49393] <= 8'h10 ;
			data[49394] <= 8'h10 ;
			data[49395] <= 8'h10 ;
			data[49396] <= 8'h10 ;
			data[49397] <= 8'h10 ;
			data[49398] <= 8'h10 ;
			data[49399] <= 8'h10 ;
			data[49400] <= 8'h10 ;
			data[49401] <= 8'h10 ;
			data[49402] <= 8'h10 ;
			data[49403] <= 8'h10 ;
			data[49404] <= 8'h10 ;
			data[49405] <= 8'h10 ;
			data[49406] <= 8'h10 ;
			data[49407] <= 8'h10 ;
			data[49408] <= 8'h10 ;
			data[49409] <= 8'h10 ;
			data[49410] <= 8'h10 ;
			data[49411] <= 8'h10 ;
			data[49412] <= 8'h10 ;
			data[49413] <= 8'h10 ;
			data[49414] <= 8'h10 ;
			data[49415] <= 8'h10 ;
			data[49416] <= 8'h10 ;
			data[49417] <= 8'h10 ;
			data[49418] <= 8'h10 ;
			data[49419] <= 8'h10 ;
			data[49420] <= 8'h10 ;
			data[49421] <= 8'h10 ;
			data[49422] <= 8'h10 ;
			data[49423] <= 8'h10 ;
			data[49424] <= 8'h10 ;
			data[49425] <= 8'h10 ;
			data[49426] <= 8'h10 ;
			data[49427] <= 8'h10 ;
			data[49428] <= 8'h10 ;
			data[49429] <= 8'h10 ;
			data[49430] <= 8'h10 ;
			data[49431] <= 8'h10 ;
			data[49432] <= 8'h10 ;
			data[49433] <= 8'h10 ;
			data[49434] <= 8'h10 ;
			data[49435] <= 8'h10 ;
			data[49436] <= 8'h10 ;
			data[49437] <= 8'h10 ;
			data[49438] <= 8'h10 ;
			data[49439] <= 8'h10 ;
			data[49440] <= 8'h10 ;
			data[49441] <= 8'h10 ;
			data[49442] <= 8'h10 ;
			data[49443] <= 8'h10 ;
			data[49444] <= 8'h10 ;
			data[49445] <= 8'h10 ;
			data[49446] <= 8'h10 ;
			data[49447] <= 8'h10 ;
			data[49448] <= 8'h10 ;
			data[49449] <= 8'h10 ;
			data[49450] <= 8'h10 ;
			data[49451] <= 8'h10 ;
			data[49452] <= 8'h10 ;
			data[49453] <= 8'h10 ;
			data[49454] <= 8'h10 ;
			data[49455] <= 8'h10 ;
			data[49456] <= 8'h10 ;
			data[49457] <= 8'h10 ;
			data[49458] <= 8'h10 ;
			data[49459] <= 8'h10 ;
			data[49460] <= 8'h10 ;
			data[49461] <= 8'h10 ;
			data[49462] <= 8'h10 ;
			data[49463] <= 8'h10 ;
			data[49464] <= 8'h10 ;
			data[49465] <= 8'h10 ;
			data[49466] <= 8'h10 ;
			data[49467] <= 8'h10 ;
			data[49468] <= 8'h10 ;
			data[49469] <= 8'h10 ;
			data[49470] <= 8'h10 ;
			data[49471] <= 8'h10 ;
			data[49472] <= 8'h10 ;
			data[49473] <= 8'h10 ;
			data[49474] <= 8'h10 ;
			data[49475] <= 8'h10 ;
			data[49476] <= 8'h10 ;
			data[49477] <= 8'h10 ;
			data[49478] <= 8'h10 ;
			data[49479] <= 8'h10 ;
			data[49480] <= 8'h10 ;
			data[49481] <= 8'h10 ;
			data[49482] <= 8'h10 ;
			data[49483] <= 8'h10 ;
			data[49484] <= 8'h10 ;
			data[49485] <= 8'h10 ;
			data[49486] <= 8'h10 ;
			data[49487] <= 8'h10 ;
			data[49488] <= 8'h10 ;
			data[49489] <= 8'h10 ;
			data[49490] <= 8'h10 ;
			data[49491] <= 8'h10 ;
			data[49492] <= 8'h10 ;
			data[49493] <= 8'h10 ;
			data[49494] <= 8'h10 ;
			data[49495] <= 8'h10 ;
			data[49496] <= 8'h10 ;
			data[49497] <= 8'h10 ;
			data[49498] <= 8'h10 ;
			data[49499] <= 8'h10 ;
			data[49500] <= 8'h10 ;
			data[49501] <= 8'h10 ;
			data[49502] <= 8'h10 ;
			data[49503] <= 8'h10 ;
			data[49504] <= 8'h10 ;
			data[49505] <= 8'h10 ;
			data[49506] <= 8'h10 ;
			data[49507] <= 8'h10 ;
			data[49508] <= 8'h10 ;
			data[49509] <= 8'h10 ;
			data[49510] <= 8'h10 ;
			data[49511] <= 8'h10 ;
			data[49512] <= 8'h10 ;
			data[49513] <= 8'h10 ;
			data[49514] <= 8'h10 ;
			data[49515] <= 8'h10 ;
			data[49516] <= 8'h10 ;
			data[49517] <= 8'h10 ;
			data[49518] <= 8'h10 ;
			data[49519] <= 8'h10 ;
			data[49520] <= 8'h10 ;
			data[49521] <= 8'h10 ;
			data[49522] <= 8'h10 ;
			data[49523] <= 8'h10 ;
			data[49524] <= 8'h10 ;
			data[49525] <= 8'h10 ;
			data[49526] <= 8'h10 ;
			data[49527] <= 8'h10 ;
			data[49528] <= 8'h10 ;
			data[49529] <= 8'h10 ;
			data[49530] <= 8'h10 ;
			data[49531] <= 8'h10 ;
			data[49532] <= 8'h10 ;
			data[49533] <= 8'h10 ;
			data[49534] <= 8'h10 ;
			data[49535] <= 8'h10 ;
			data[49536] <= 8'h10 ;
			data[49537] <= 8'h10 ;
			data[49538] <= 8'h10 ;
			data[49539] <= 8'h10 ;
			data[49540] <= 8'h10 ;
			data[49541] <= 8'h10 ;
			data[49542] <= 8'h10 ;
			data[49543] <= 8'h10 ;
			data[49544] <= 8'h10 ;
			data[49545] <= 8'h10 ;
			data[49546] <= 8'h10 ;
			data[49547] <= 8'h10 ;
			data[49548] <= 8'h10 ;
			data[49549] <= 8'h10 ;
			data[49550] <= 8'h10 ;
			data[49551] <= 8'h10 ;
			data[49552] <= 8'h10 ;
			data[49553] <= 8'h10 ;
			data[49554] <= 8'h10 ;
			data[49555] <= 8'h10 ;
			data[49556] <= 8'h10 ;
			data[49557] <= 8'h10 ;
			data[49558] <= 8'h10 ;
			data[49559] <= 8'h10 ;
			data[49560] <= 8'h10 ;
			data[49561] <= 8'h10 ;
			data[49562] <= 8'h10 ;
			data[49563] <= 8'h10 ;
			data[49564] <= 8'h10 ;
			data[49565] <= 8'h10 ;
			data[49566] <= 8'h10 ;
			data[49567] <= 8'h10 ;
			data[49568] <= 8'h10 ;
			data[49569] <= 8'h10 ;
			data[49570] <= 8'h10 ;
			data[49571] <= 8'h10 ;
			data[49572] <= 8'h10 ;
			data[49573] <= 8'h10 ;
			data[49574] <= 8'h10 ;
			data[49575] <= 8'h10 ;
			data[49576] <= 8'h10 ;
			data[49577] <= 8'h10 ;
			data[49578] <= 8'h10 ;
			data[49579] <= 8'h10 ;
			data[49580] <= 8'h10 ;
			data[49581] <= 8'h10 ;
			data[49582] <= 8'h10 ;
			data[49583] <= 8'h10 ;
			data[49584] <= 8'h10 ;
			data[49585] <= 8'h10 ;
			data[49586] <= 8'h10 ;
			data[49587] <= 8'h10 ;
			data[49588] <= 8'h10 ;
			data[49589] <= 8'h10 ;
			data[49590] <= 8'h10 ;
			data[49591] <= 8'h10 ;
			data[49592] <= 8'h10 ;
			data[49593] <= 8'h10 ;
			data[49594] <= 8'h10 ;
			data[49595] <= 8'h10 ;
			data[49596] <= 8'h10 ;
			data[49597] <= 8'h10 ;
			data[49598] <= 8'h10 ;
			data[49599] <= 8'h10 ;
			data[49600] <= 8'h10 ;
			data[49601] <= 8'h10 ;
			data[49602] <= 8'h10 ;
			data[49603] <= 8'h10 ;
			data[49604] <= 8'h10 ;
			data[49605] <= 8'h10 ;
			data[49606] <= 8'h10 ;
			data[49607] <= 8'h10 ;
			data[49608] <= 8'h10 ;
			data[49609] <= 8'h10 ;
			data[49610] <= 8'h10 ;
			data[49611] <= 8'h10 ;
			data[49612] <= 8'h10 ;
			data[49613] <= 8'h10 ;
			data[49614] <= 8'h10 ;
			data[49615] <= 8'h10 ;
			data[49616] <= 8'h10 ;
			data[49617] <= 8'h10 ;
			data[49618] <= 8'h10 ;
			data[49619] <= 8'h10 ;
			data[49620] <= 8'h10 ;
			data[49621] <= 8'h10 ;
			data[49622] <= 8'h10 ;
			data[49623] <= 8'h10 ;
			data[49624] <= 8'h10 ;
			data[49625] <= 8'h10 ;
			data[49626] <= 8'h10 ;
			data[49627] <= 8'h10 ;
			data[49628] <= 8'h10 ;
			data[49629] <= 8'h10 ;
			data[49630] <= 8'h10 ;
			data[49631] <= 8'h10 ;
			data[49632] <= 8'h10 ;
			data[49633] <= 8'h10 ;
			data[49634] <= 8'h10 ;
			data[49635] <= 8'h10 ;
			data[49636] <= 8'h10 ;
			data[49637] <= 8'h10 ;
			data[49638] <= 8'h10 ;
			data[49639] <= 8'h10 ;
			data[49640] <= 8'h10 ;
			data[49641] <= 8'h10 ;
			data[49642] <= 8'h10 ;
			data[49643] <= 8'h10 ;
			data[49644] <= 8'h10 ;
			data[49645] <= 8'h10 ;
			data[49646] <= 8'h10 ;
			data[49647] <= 8'h10 ;
			data[49648] <= 8'h10 ;
			data[49649] <= 8'h10 ;
			data[49650] <= 8'h10 ;
			data[49651] <= 8'h10 ;
			data[49652] <= 8'h10 ;
			data[49653] <= 8'h10 ;
			data[49654] <= 8'h10 ;
			data[49655] <= 8'h10 ;
			data[49656] <= 8'h10 ;
			data[49657] <= 8'h10 ;
			data[49658] <= 8'h10 ;
			data[49659] <= 8'h10 ;
			data[49660] <= 8'h10 ;
			data[49661] <= 8'h10 ;
			data[49662] <= 8'h10 ;
			data[49663] <= 8'h10 ;
			data[49664] <= 8'h10 ;
			data[49665] <= 8'h10 ;
			data[49666] <= 8'h10 ;
			data[49667] <= 8'h10 ;
			data[49668] <= 8'h10 ;
			data[49669] <= 8'h10 ;
			data[49670] <= 8'h10 ;
			data[49671] <= 8'h10 ;
			data[49672] <= 8'h10 ;
			data[49673] <= 8'h10 ;
			data[49674] <= 8'h10 ;
			data[49675] <= 8'h10 ;
			data[49676] <= 8'h10 ;
			data[49677] <= 8'h10 ;
			data[49678] <= 8'h10 ;
			data[49679] <= 8'h10 ;
			data[49680] <= 8'h10 ;
			data[49681] <= 8'h10 ;
			data[49682] <= 8'h10 ;
			data[49683] <= 8'h10 ;
			data[49684] <= 8'h10 ;
			data[49685] <= 8'h10 ;
			data[49686] <= 8'h10 ;
			data[49687] <= 8'h10 ;
			data[49688] <= 8'h10 ;
			data[49689] <= 8'h10 ;
			data[49690] <= 8'h10 ;
			data[49691] <= 8'h10 ;
			data[49692] <= 8'h10 ;
			data[49693] <= 8'h10 ;
			data[49694] <= 8'h10 ;
			data[49695] <= 8'h10 ;
			data[49696] <= 8'h10 ;
			data[49697] <= 8'h10 ;
			data[49698] <= 8'h10 ;
			data[49699] <= 8'h10 ;
			data[49700] <= 8'h10 ;
			data[49701] <= 8'h10 ;
			data[49702] <= 8'h10 ;
			data[49703] <= 8'h10 ;
			data[49704] <= 8'h10 ;
			data[49705] <= 8'h10 ;
			data[49706] <= 8'h10 ;
			data[49707] <= 8'h10 ;
			data[49708] <= 8'h10 ;
			data[49709] <= 8'h10 ;
			data[49710] <= 8'h10 ;
			data[49711] <= 8'h10 ;
			data[49712] <= 8'h10 ;
			data[49713] <= 8'h10 ;
			data[49714] <= 8'h10 ;
			data[49715] <= 8'h10 ;
			data[49716] <= 8'h10 ;
			data[49717] <= 8'h10 ;
			data[49718] <= 8'h10 ;
			data[49719] <= 8'h10 ;
			data[49720] <= 8'h10 ;
			data[49721] <= 8'h10 ;
			data[49722] <= 8'h10 ;
			data[49723] <= 8'h10 ;
			data[49724] <= 8'h10 ;
			data[49725] <= 8'h10 ;
			data[49726] <= 8'h10 ;
			data[49727] <= 8'h10 ;
			data[49728] <= 8'h10 ;
			data[49729] <= 8'h10 ;
			data[49730] <= 8'h10 ;
			data[49731] <= 8'h10 ;
			data[49732] <= 8'h10 ;
			data[49733] <= 8'h10 ;
			data[49734] <= 8'h10 ;
			data[49735] <= 8'h10 ;
			data[49736] <= 8'h10 ;
			data[49737] <= 8'h10 ;
			data[49738] <= 8'h10 ;
			data[49739] <= 8'h10 ;
			data[49740] <= 8'h10 ;
			data[49741] <= 8'h10 ;
			data[49742] <= 8'h10 ;
			data[49743] <= 8'h10 ;
			data[49744] <= 8'h10 ;
			data[49745] <= 8'h10 ;
			data[49746] <= 8'h10 ;
			data[49747] <= 8'h10 ;
			data[49748] <= 8'h10 ;
			data[49749] <= 8'h10 ;
			data[49750] <= 8'h10 ;
			data[49751] <= 8'h10 ;
			data[49752] <= 8'h10 ;
			data[49753] <= 8'h10 ;
			data[49754] <= 8'h10 ;
			data[49755] <= 8'h10 ;
			data[49756] <= 8'h10 ;
			data[49757] <= 8'h10 ;
			data[49758] <= 8'h10 ;
			data[49759] <= 8'h10 ;
			data[49760] <= 8'h10 ;
			data[49761] <= 8'h10 ;
			data[49762] <= 8'h10 ;
			data[49763] <= 8'h10 ;
			data[49764] <= 8'h10 ;
			data[49765] <= 8'h10 ;
			data[49766] <= 8'h10 ;
			data[49767] <= 8'h10 ;
			data[49768] <= 8'h10 ;
			data[49769] <= 8'h10 ;
			data[49770] <= 8'h10 ;
			data[49771] <= 8'h10 ;
			data[49772] <= 8'h10 ;
			data[49773] <= 8'h10 ;
			data[49774] <= 8'h10 ;
			data[49775] <= 8'h10 ;
			data[49776] <= 8'h10 ;
			data[49777] <= 8'h10 ;
			data[49778] <= 8'h10 ;
			data[49779] <= 8'h10 ;
			data[49780] <= 8'h10 ;
			data[49781] <= 8'h10 ;
			data[49782] <= 8'h10 ;
			data[49783] <= 8'h10 ;
			data[49784] <= 8'h10 ;
			data[49785] <= 8'h10 ;
			data[49786] <= 8'h10 ;
			data[49787] <= 8'h10 ;
			data[49788] <= 8'h10 ;
			data[49789] <= 8'h10 ;
			data[49790] <= 8'h10 ;
			data[49791] <= 8'h10 ;
			data[49792] <= 8'h10 ;
			data[49793] <= 8'h10 ;
			data[49794] <= 8'h10 ;
			data[49795] <= 8'h10 ;
			data[49796] <= 8'h10 ;
			data[49797] <= 8'h10 ;
			data[49798] <= 8'h10 ;
			data[49799] <= 8'h10 ;
			data[49800] <= 8'h10 ;
			data[49801] <= 8'h10 ;
			data[49802] <= 8'h10 ;
			data[49803] <= 8'h10 ;
			data[49804] <= 8'h10 ;
			data[49805] <= 8'h10 ;
			data[49806] <= 8'h10 ;
			data[49807] <= 8'h10 ;
			data[49808] <= 8'h10 ;
			data[49809] <= 8'h10 ;
			data[49810] <= 8'h10 ;
			data[49811] <= 8'h10 ;
			data[49812] <= 8'h10 ;
			data[49813] <= 8'h10 ;
			data[49814] <= 8'h10 ;
			data[49815] <= 8'h10 ;
			data[49816] <= 8'h10 ;
			data[49817] <= 8'h10 ;
			data[49818] <= 8'h10 ;
			data[49819] <= 8'h10 ;
			data[49820] <= 8'h10 ;
			data[49821] <= 8'h10 ;
			data[49822] <= 8'h10 ;
			data[49823] <= 8'h10 ;
			data[49824] <= 8'h10 ;
			data[49825] <= 8'h10 ;
			data[49826] <= 8'h10 ;
			data[49827] <= 8'h10 ;
			data[49828] <= 8'h10 ;
			data[49829] <= 8'h10 ;
			data[49830] <= 8'h10 ;
			data[49831] <= 8'h10 ;
			data[49832] <= 8'h10 ;
			data[49833] <= 8'h10 ;
			data[49834] <= 8'h10 ;
			data[49835] <= 8'h10 ;
			data[49836] <= 8'h10 ;
			data[49837] <= 8'h10 ;
			data[49838] <= 8'h10 ;
			data[49839] <= 8'h10 ;
			data[49840] <= 8'h10 ;
			data[49841] <= 8'h10 ;
			data[49842] <= 8'h10 ;
			data[49843] <= 8'h10 ;
			data[49844] <= 8'h10 ;
			data[49845] <= 8'h10 ;
			data[49846] <= 8'h10 ;
			data[49847] <= 8'h10 ;
			data[49848] <= 8'h10 ;
			data[49849] <= 8'h10 ;
			data[49850] <= 8'h10 ;
			data[49851] <= 8'h10 ;
			data[49852] <= 8'h10 ;
			data[49853] <= 8'h10 ;
			data[49854] <= 8'h10 ;
			data[49855] <= 8'h10 ;
			data[49856] <= 8'h10 ;
			data[49857] <= 8'h10 ;
			data[49858] <= 8'h10 ;
			data[49859] <= 8'h10 ;
			data[49860] <= 8'h10 ;
			data[49861] <= 8'h10 ;
			data[49862] <= 8'h10 ;
			data[49863] <= 8'h10 ;
			data[49864] <= 8'h10 ;
			data[49865] <= 8'h10 ;
			data[49866] <= 8'h10 ;
			data[49867] <= 8'h10 ;
			data[49868] <= 8'h10 ;
			data[49869] <= 8'h10 ;
			data[49870] <= 8'h10 ;
			data[49871] <= 8'h10 ;
			data[49872] <= 8'h10 ;
			data[49873] <= 8'h10 ;
			data[49874] <= 8'h10 ;
			data[49875] <= 8'h10 ;
			data[49876] <= 8'h10 ;
			data[49877] <= 8'h10 ;
			data[49878] <= 8'h10 ;
			data[49879] <= 8'h10 ;
			data[49880] <= 8'h10 ;
			data[49881] <= 8'h10 ;
			data[49882] <= 8'h10 ;
			data[49883] <= 8'h10 ;
			data[49884] <= 8'h10 ;
			data[49885] <= 8'h10 ;
			data[49886] <= 8'h10 ;
			data[49887] <= 8'h10 ;
			data[49888] <= 8'h10 ;
			data[49889] <= 8'h10 ;
			data[49890] <= 8'h10 ;
			data[49891] <= 8'h10 ;
			data[49892] <= 8'h10 ;
			data[49893] <= 8'h10 ;
			data[49894] <= 8'h10 ;
			data[49895] <= 8'h10 ;
			data[49896] <= 8'h10 ;
			data[49897] <= 8'h10 ;
			data[49898] <= 8'h10 ;
			data[49899] <= 8'h10 ;
			data[49900] <= 8'h10 ;
			data[49901] <= 8'h10 ;
			data[49902] <= 8'h10 ;
			data[49903] <= 8'h10 ;
			data[49904] <= 8'h10 ;
			data[49905] <= 8'h10 ;
			data[49906] <= 8'h10 ;
			data[49907] <= 8'h10 ;
			data[49908] <= 8'h10 ;
			data[49909] <= 8'h10 ;
			data[49910] <= 8'h10 ;
			data[49911] <= 8'h10 ;
			data[49912] <= 8'h10 ;
			data[49913] <= 8'h10 ;
			data[49914] <= 8'h10 ;
			data[49915] <= 8'h10 ;
			data[49916] <= 8'h10 ;
			data[49917] <= 8'h10 ;
			data[49918] <= 8'h10 ;
			data[49919] <= 8'h10 ;
			data[49920] <= 8'h10 ;
			data[49921] <= 8'h10 ;
			data[49922] <= 8'h10 ;
			data[49923] <= 8'h10 ;
			data[49924] <= 8'h10 ;
			data[49925] <= 8'h10 ;
			data[49926] <= 8'h10 ;
			data[49927] <= 8'h10 ;
			data[49928] <= 8'h10 ;
			data[49929] <= 8'h10 ;
			data[49930] <= 8'h10 ;
			data[49931] <= 8'h10 ;
			data[49932] <= 8'h10 ;
			data[49933] <= 8'h10 ;
			data[49934] <= 8'h10 ;
			data[49935] <= 8'h10 ;
			data[49936] <= 8'h10 ;
			data[49937] <= 8'h10 ;
			data[49938] <= 8'h10 ;
			data[49939] <= 8'h10 ;
			data[49940] <= 8'h10 ;
			data[49941] <= 8'h10 ;
			data[49942] <= 8'h10 ;
			data[49943] <= 8'h10 ;
			data[49944] <= 8'h10 ;
			data[49945] <= 8'h10 ;
			data[49946] <= 8'h10 ;
			data[49947] <= 8'h10 ;
			data[49948] <= 8'h10 ;
			data[49949] <= 8'h10 ;
			data[49950] <= 8'h10 ;
			data[49951] <= 8'h10 ;
			data[49952] <= 8'h10 ;
			data[49953] <= 8'h10 ;
			data[49954] <= 8'h10 ;
			data[49955] <= 8'h10 ;
			data[49956] <= 8'h10 ;
			data[49957] <= 8'h10 ;
			data[49958] <= 8'h10 ;
			data[49959] <= 8'h10 ;
			data[49960] <= 8'h10 ;
			data[49961] <= 8'h10 ;
			data[49962] <= 8'h10 ;
			data[49963] <= 8'h10 ;
			data[49964] <= 8'h10 ;
			data[49965] <= 8'h10 ;
			data[49966] <= 8'h10 ;
			data[49967] <= 8'h10 ;
			data[49968] <= 8'h10 ;
			data[49969] <= 8'h10 ;
			data[49970] <= 8'h10 ;
			data[49971] <= 8'h10 ;
			data[49972] <= 8'h10 ;
			data[49973] <= 8'h10 ;
			data[49974] <= 8'h10 ;
			data[49975] <= 8'h10 ;
			data[49976] <= 8'h10 ;
			data[49977] <= 8'h10 ;
			data[49978] <= 8'h10 ;
			data[49979] <= 8'h10 ;
			data[49980] <= 8'h10 ;
			data[49981] <= 8'h10 ;
			data[49982] <= 8'h10 ;
			data[49983] <= 8'h10 ;
			data[49984] <= 8'h10 ;
			data[49985] <= 8'h10 ;
			data[49986] <= 8'h10 ;
			data[49987] <= 8'h10 ;
			data[49988] <= 8'h10 ;
			data[49989] <= 8'h10 ;
			data[49990] <= 8'h10 ;
			data[49991] <= 8'h10 ;
			data[49992] <= 8'h10 ;
			data[49993] <= 8'h10 ;
			data[49994] <= 8'h10 ;
			data[49995] <= 8'h10 ;
			data[49996] <= 8'h10 ;
			data[49997] <= 8'h10 ;
			data[49998] <= 8'h10 ;
			data[49999] <= 8'h10 ;
			data[50000] <= 8'h10 ;
			data[50001] <= 8'h10 ;
			data[50002] <= 8'h10 ;
			data[50003] <= 8'h10 ;
			data[50004] <= 8'h10 ;
			data[50005] <= 8'h10 ;
			data[50006] <= 8'h10 ;
			data[50007] <= 8'h10 ;
			data[50008] <= 8'h10 ;
			data[50009] <= 8'h10 ;
			data[50010] <= 8'h10 ;
			data[50011] <= 8'h10 ;
			data[50012] <= 8'h10 ;
			data[50013] <= 8'h10 ;
			data[50014] <= 8'h10 ;
			data[50015] <= 8'h10 ;
			data[50016] <= 8'h10 ;
			data[50017] <= 8'h10 ;
			data[50018] <= 8'h10 ;
			data[50019] <= 8'h10 ;
			data[50020] <= 8'h10 ;
			data[50021] <= 8'h10 ;
			data[50022] <= 8'h10 ;
			data[50023] <= 8'h10 ;
			data[50024] <= 8'h10 ;
			data[50025] <= 8'h10 ;
			data[50026] <= 8'h10 ;
			data[50027] <= 8'h10 ;
			data[50028] <= 8'h10 ;
			data[50029] <= 8'h10 ;
			data[50030] <= 8'h10 ;
			data[50031] <= 8'h10 ;
			data[50032] <= 8'h10 ;
			data[50033] <= 8'h10 ;
			data[50034] <= 8'h10 ;
			data[50035] <= 8'h10 ;
			data[50036] <= 8'h10 ;
			data[50037] <= 8'h10 ;
			data[50038] <= 8'h10 ;
			data[50039] <= 8'h10 ;
			data[50040] <= 8'h10 ;
			data[50041] <= 8'h10 ;
			data[50042] <= 8'h10 ;
			data[50043] <= 8'h10 ;
			data[50044] <= 8'h10 ;
			data[50045] <= 8'h10 ;
			data[50046] <= 8'h10 ;
			data[50047] <= 8'h10 ;
			data[50048] <= 8'h10 ;
			data[50049] <= 8'h10 ;
			data[50050] <= 8'h10 ;
			data[50051] <= 8'h10 ;
			data[50052] <= 8'h10 ;
			data[50053] <= 8'h10 ;
			data[50054] <= 8'h10 ;
			data[50055] <= 8'h10 ;
			data[50056] <= 8'h10 ;
			data[50057] <= 8'h10 ;
			data[50058] <= 8'h10 ;
			data[50059] <= 8'h10 ;
			data[50060] <= 8'h10 ;
			data[50061] <= 8'h10 ;
			data[50062] <= 8'h10 ;
			data[50063] <= 8'h10 ;
			data[50064] <= 8'h10 ;
			data[50065] <= 8'h10 ;
			data[50066] <= 8'h10 ;
			data[50067] <= 8'h10 ;
			data[50068] <= 8'h10 ;
			data[50069] <= 8'h10 ;
			data[50070] <= 8'h10 ;
			data[50071] <= 8'h10 ;
			data[50072] <= 8'h10 ;
			data[50073] <= 8'h10 ;
			data[50074] <= 8'h10 ;
			data[50075] <= 8'h10 ;
			data[50076] <= 8'h10 ;
			data[50077] <= 8'h10 ;
			data[50078] <= 8'h10 ;
			data[50079] <= 8'h10 ;
			data[50080] <= 8'h10 ;
			data[50081] <= 8'h10 ;
			data[50082] <= 8'h10 ;
			data[50083] <= 8'h10 ;
			data[50084] <= 8'h10 ;
			data[50085] <= 8'h10 ;
			data[50086] <= 8'h10 ;
			data[50087] <= 8'h10 ;
			data[50088] <= 8'h10 ;
			data[50089] <= 8'h10 ;
			data[50090] <= 8'h10 ;
			data[50091] <= 8'h10 ;
			data[50092] <= 8'h10 ;
			data[50093] <= 8'h10 ;
			data[50094] <= 8'h10 ;
			data[50095] <= 8'h10 ;
			data[50096] <= 8'h10 ;
			data[50097] <= 8'h10 ;
			data[50098] <= 8'h10 ;
			data[50099] <= 8'h10 ;
			data[50100] <= 8'h10 ;
			data[50101] <= 8'h10 ;
			data[50102] <= 8'h10 ;
			data[50103] <= 8'h10 ;
			data[50104] <= 8'h10 ;
			data[50105] <= 8'h10 ;
			data[50106] <= 8'h10 ;
			data[50107] <= 8'h10 ;
			data[50108] <= 8'h10 ;
			data[50109] <= 8'h10 ;
			data[50110] <= 8'h10 ;
			data[50111] <= 8'h10 ;
			data[50112] <= 8'h10 ;
			data[50113] <= 8'h10 ;
			data[50114] <= 8'h10 ;
			data[50115] <= 8'h10 ;
			data[50116] <= 8'h10 ;
			data[50117] <= 8'h10 ;
			data[50118] <= 8'h10 ;
			data[50119] <= 8'h10 ;
			data[50120] <= 8'h10 ;
			data[50121] <= 8'h10 ;
			data[50122] <= 8'h10 ;
			data[50123] <= 8'h10 ;
			data[50124] <= 8'h10 ;
			data[50125] <= 8'h10 ;
			data[50126] <= 8'h10 ;
			data[50127] <= 8'h10 ;
			data[50128] <= 8'h10 ;
			data[50129] <= 8'h10 ;
			data[50130] <= 8'h10 ;
			data[50131] <= 8'h10 ;
			data[50132] <= 8'h10 ;
			data[50133] <= 8'h10 ;
			data[50134] <= 8'h10 ;
			data[50135] <= 8'h10 ;
			data[50136] <= 8'h10 ;
			data[50137] <= 8'h10 ;
			data[50138] <= 8'h10 ;
			data[50139] <= 8'h10 ;
			data[50140] <= 8'h10 ;
			data[50141] <= 8'h10 ;
			data[50142] <= 8'h10 ;
			data[50143] <= 8'h10 ;
			data[50144] <= 8'h10 ;
			data[50145] <= 8'h10 ;
			data[50146] <= 8'h10 ;
			data[50147] <= 8'h10 ;
			data[50148] <= 8'h10 ;
			data[50149] <= 8'h10 ;
			data[50150] <= 8'h10 ;
			data[50151] <= 8'h10 ;
			data[50152] <= 8'h10 ;
			data[50153] <= 8'h10 ;
			data[50154] <= 8'h10 ;
			data[50155] <= 8'h10 ;
			data[50156] <= 8'h10 ;
			data[50157] <= 8'h10 ;
			data[50158] <= 8'h10 ;
			data[50159] <= 8'h10 ;
			data[50160] <= 8'h10 ;
			data[50161] <= 8'h10 ;
			data[50162] <= 8'h10 ;
			data[50163] <= 8'h10 ;
			data[50164] <= 8'h10 ;
			data[50165] <= 8'h10 ;
			data[50166] <= 8'h10 ;
			data[50167] <= 8'h10 ;
			data[50168] <= 8'h10 ;
			data[50169] <= 8'h10 ;
			data[50170] <= 8'h10 ;
			data[50171] <= 8'h10 ;
			data[50172] <= 8'h10 ;
			data[50173] <= 8'h10 ;
			data[50174] <= 8'h10 ;
			data[50175] <= 8'h10 ;
			data[50176] <= 8'h10 ;
			data[50177] <= 8'h10 ;
			data[50178] <= 8'h10 ;
			data[50179] <= 8'h10 ;
			data[50180] <= 8'h10 ;
			data[50181] <= 8'h10 ;
			data[50182] <= 8'h10 ;
			data[50183] <= 8'h10 ;
			data[50184] <= 8'h10 ;
			data[50185] <= 8'h10 ;
			data[50186] <= 8'h10 ;
			data[50187] <= 8'h10 ;
			data[50188] <= 8'h10 ;
			data[50189] <= 8'h10 ;
			data[50190] <= 8'h10 ;
			data[50191] <= 8'h10 ;
			data[50192] <= 8'h10 ;
			data[50193] <= 8'h10 ;
			data[50194] <= 8'h10 ;
			data[50195] <= 8'h10 ;
			data[50196] <= 8'h10 ;
			data[50197] <= 8'h10 ;
			data[50198] <= 8'h10 ;
			data[50199] <= 8'h10 ;
			data[50200] <= 8'h10 ;
			data[50201] <= 8'h10 ;
			data[50202] <= 8'h10 ;
			data[50203] <= 8'h10 ;
			data[50204] <= 8'h10 ;
			data[50205] <= 8'h10 ;
			data[50206] <= 8'h10 ;
			data[50207] <= 8'h10 ;
			data[50208] <= 8'h10 ;
			data[50209] <= 8'h10 ;
			data[50210] <= 8'h10 ;
			data[50211] <= 8'h10 ;
			data[50212] <= 8'h10 ;
			data[50213] <= 8'h10 ;
			data[50214] <= 8'h10 ;
			data[50215] <= 8'h10 ;
			data[50216] <= 8'h10 ;
			data[50217] <= 8'h10 ;
			data[50218] <= 8'h10 ;
			data[50219] <= 8'h10 ;
			data[50220] <= 8'h10 ;
			data[50221] <= 8'h10 ;
			data[50222] <= 8'h10 ;
			data[50223] <= 8'h10 ;
			data[50224] <= 8'h10 ;
			data[50225] <= 8'h10 ;
			data[50226] <= 8'h10 ;
			data[50227] <= 8'h10 ;
			data[50228] <= 8'h10 ;
			data[50229] <= 8'h10 ;
			data[50230] <= 8'h10 ;
			data[50231] <= 8'h10 ;
			data[50232] <= 8'h10 ;
			data[50233] <= 8'h10 ;
			data[50234] <= 8'h10 ;
			data[50235] <= 8'h10 ;
			data[50236] <= 8'h10 ;
			data[50237] <= 8'h10 ;
			data[50238] <= 8'h10 ;
			data[50239] <= 8'h10 ;
			data[50240] <= 8'h10 ;
			data[50241] <= 8'h10 ;
			data[50242] <= 8'h10 ;
			data[50243] <= 8'h10 ;
			data[50244] <= 8'h10 ;
			data[50245] <= 8'h10 ;
			data[50246] <= 8'h10 ;
			data[50247] <= 8'h10 ;
			data[50248] <= 8'h10 ;
			data[50249] <= 8'h10 ;
			data[50250] <= 8'h10 ;
			data[50251] <= 8'h10 ;
			data[50252] <= 8'h10 ;
			data[50253] <= 8'h10 ;
			data[50254] <= 8'h10 ;
			data[50255] <= 8'h10 ;
			data[50256] <= 8'h10 ;
			data[50257] <= 8'h10 ;
			data[50258] <= 8'h10 ;
			data[50259] <= 8'h10 ;
			data[50260] <= 8'h10 ;
			data[50261] <= 8'h10 ;
			data[50262] <= 8'h10 ;
			data[50263] <= 8'h10 ;
			data[50264] <= 8'h10 ;
			data[50265] <= 8'h10 ;
			data[50266] <= 8'h10 ;
			data[50267] <= 8'h10 ;
			data[50268] <= 8'h10 ;
			data[50269] <= 8'h10 ;
			data[50270] <= 8'h10 ;
			data[50271] <= 8'h10 ;
			data[50272] <= 8'h10 ;
			data[50273] <= 8'h10 ;
			data[50274] <= 8'h10 ;
			data[50275] <= 8'h10 ;
			data[50276] <= 8'h10 ;
			data[50277] <= 8'h10 ;
			data[50278] <= 8'h10 ;
			data[50279] <= 8'h10 ;
			data[50280] <= 8'h10 ;
			data[50281] <= 8'h10 ;
			data[50282] <= 8'h10 ;
			data[50283] <= 8'h10 ;
			data[50284] <= 8'h10 ;
			data[50285] <= 8'h10 ;
			data[50286] <= 8'h10 ;
			data[50287] <= 8'h10 ;
			data[50288] <= 8'h10 ;
			data[50289] <= 8'h10 ;
			data[50290] <= 8'h10 ;
			data[50291] <= 8'h10 ;
			data[50292] <= 8'h10 ;
			data[50293] <= 8'h10 ;
			data[50294] <= 8'h10 ;
			data[50295] <= 8'h10 ;
			data[50296] <= 8'h10 ;
			data[50297] <= 8'h10 ;
			data[50298] <= 8'h10 ;
			data[50299] <= 8'h10 ;
			data[50300] <= 8'h10 ;
			data[50301] <= 8'h10 ;
			data[50302] <= 8'h10 ;
			data[50303] <= 8'h10 ;
			data[50304] <= 8'h10 ;
			data[50305] <= 8'h10 ;
			data[50306] <= 8'h10 ;
			data[50307] <= 8'h10 ;
			data[50308] <= 8'h10 ;
			data[50309] <= 8'h10 ;
			data[50310] <= 8'h10 ;
			data[50311] <= 8'h10 ;
			data[50312] <= 8'h10 ;
			data[50313] <= 8'h10 ;
			data[50314] <= 8'h10 ;
			data[50315] <= 8'h10 ;
			data[50316] <= 8'h10 ;
			data[50317] <= 8'h10 ;
			data[50318] <= 8'h10 ;
			data[50319] <= 8'h10 ;
			data[50320] <= 8'h10 ;
			data[50321] <= 8'h10 ;
			data[50322] <= 8'h10 ;
			data[50323] <= 8'h10 ;
			data[50324] <= 8'h10 ;
			data[50325] <= 8'h10 ;
			data[50326] <= 8'h10 ;
			data[50327] <= 8'h10 ;
			data[50328] <= 8'h10 ;
			data[50329] <= 8'h10 ;
			data[50330] <= 8'h10 ;
			data[50331] <= 8'h10 ;
			data[50332] <= 8'h10 ;
			data[50333] <= 8'h10 ;
			data[50334] <= 8'h10 ;
			data[50335] <= 8'h10 ;
			data[50336] <= 8'h10 ;
			data[50337] <= 8'h10 ;
			data[50338] <= 8'h10 ;
			data[50339] <= 8'h10 ;
			data[50340] <= 8'h10 ;
			data[50341] <= 8'h10 ;
			data[50342] <= 8'h10 ;
			data[50343] <= 8'h10 ;
			data[50344] <= 8'h10 ;
			data[50345] <= 8'h10 ;
			data[50346] <= 8'h10 ;
			data[50347] <= 8'h10 ;
			data[50348] <= 8'h10 ;
			data[50349] <= 8'h10 ;
			data[50350] <= 8'h10 ;
			data[50351] <= 8'h10 ;
			data[50352] <= 8'h10 ;
			data[50353] <= 8'h10 ;
			data[50354] <= 8'h10 ;
			data[50355] <= 8'h10 ;
			data[50356] <= 8'h10 ;
			data[50357] <= 8'h10 ;
			data[50358] <= 8'h10 ;
			data[50359] <= 8'h10 ;
			data[50360] <= 8'h10 ;
			data[50361] <= 8'h10 ;
			data[50362] <= 8'h10 ;
			data[50363] <= 8'h10 ;
			data[50364] <= 8'h10 ;
			data[50365] <= 8'h10 ;
			data[50366] <= 8'h10 ;
			data[50367] <= 8'h10 ;
			data[50368] <= 8'h10 ;
			data[50369] <= 8'h10 ;
			data[50370] <= 8'h10 ;
			data[50371] <= 8'h10 ;
			data[50372] <= 8'h10 ;
			data[50373] <= 8'h10 ;
			data[50374] <= 8'h10 ;
			data[50375] <= 8'h10 ;
			data[50376] <= 8'h10 ;
			data[50377] <= 8'h10 ;
			data[50378] <= 8'h10 ;
			data[50379] <= 8'h10 ;
			data[50380] <= 8'h10 ;
			data[50381] <= 8'h10 ;
			data[50382] <= 8'h10 ;
			data[50383] <= 8'h10 ;
			data[50384] <= 8'h10 ;
			data[50385] <= 8'h10 ;
			data[50386] <= 8'h10 ;
			data[50387] <= 8'h10 ;
			data[50388] <= 8'h10 ;
			data[50389] <= 8'h10 ;
			data[50390] <= 8'h10 ;
			data[50391] <= 8'h10 ;
			data[50392] <= 8'h10 ;
			data[50393] <= 8'h10 ;
			data[50394] <= 8'h10 ;
			data[50395] <= 8'h10 ;
			data[50396] <= 8'h10 ;
			data[50397] <= 8'h10 ;
			data[50398] <= 8'h10 ;
			data[50399] <= 8'h10 ;
			data[50400] <= 8'h10 ;
			data[50401] <= 8'h10 ;
			data[50402] <= 8'h10 ;
			data[50403] <= 8'h10 ;
			data[50404] <= 8'h10 ;
			data[50405] <= 8'h10 ;
			data[50406] <= 8'h10 ;
			data[50407] <= 8'h10 ;
			data[50408] <= 8'h10 ;
			data[50409] <= 8'h10 ;
			data[50410] <= 8'h10 ;
			data[50411] <= 8'h10 ;
			data[50412] <= 8'h10 ;
			data[50413] <= 8'h10 ;
			data[50414] <= 8'h10 ;
			data[50415] <= 8'h10 ;
			data[50416] <= 8'h10 ;
			data[50417] <= 8'h10 ;
			data[50418] <= 8'h10 ;
			data[50419] <= 8'h10 ;
			data[50420] <= 8'h10 ;
			data[50421] <= 8'h10 ;
			data[50422] <= 8'h10 ;
			data[50423] <= 8'h10 ;
			data[50424] <= 8'h10 ;
			data[50425] <= 8'h10 ;
			data[50426] <= 8'h10 ;
			data[50427] <= 8'h10 ;
			data[50428] <= 8'h10 ;
			data[50429] <= 8'h10 ;
			data[50430] <= 8'h10 ;
			data[50431] <= 8'h10 ;
			data[50432] <= 8'h10 ;
			data[50433] <= 8'h10 ;
			data[50434] <= 8'h10 ;
			data[50435] <= 8'h10 ;
			data[50436] <= 8'h10 ;
			data[50437] <= 8'h10 ;
			data[50438] <= 8'h10 ;
			data[50439] <= 8'h10 ;
			data[50440] <= 8'h10 ;
			data[50441] <= 8'h10 ;
			data[50442] <= 8'h10 ;
			data[50443] <= 8'h10 ;
			data[50444] <= 8'h10 ;
			data[50445] <= 8'h10 ;
			data[50446] <= 8'h10 ;
			data[50447] <= 8'h10 ;
			data[50448] <= 8'h10 ;
			data[50449] <= 8'h10 ;
			data[50450] <= 8'h10 ;
			data[50451] <= 8'h10 ;
			data[50452] <= 8'h10 ;
			data[50453] <= 8'h10 ;
			data[50454] <= 8'h10 ;
			data[50455] <= 8'h10 ;
			data[50456] <= 8'h10 ;
			data[50457] <= 8'h10 ;
			data[50458] <= 8'h10 ;
			data[50459] <= 8'h10 ;
			data[50460] <= 8'h10 ;
			data[50461] <= 8'h10 ;
			data[50462] <= 8'h10 ;
			data[50463] <= 8'h10 ;
			data[50464] <= 8'h10 ;
			data[50465] <= 8'h10 ;
			data[50466] <= 8'h10 ;
			data[50467] <= 8'h10 ;
			data[50468] <= 8'h10 ;
			data[50469] <= 8'h10 ;
			data[50470] <= 8'h10 ;
			data[50471] <= 8'h10 ;
			data[50472] <= 8'h10 ;
			data[50473] <= 8'h10 ;
			data[50474] <= 8'h10 ;
			data[50475] <= 8'h10 ;
			data[50476] <= 8'h10 ;
			data[50477] <= 8'h10 ;
			data[50478] <= 8'h10 ;
			data[50479] <= 8'h10 ;
			data[50480] <= 8'h10 ;
			data[50481] <= 8'h10 ;
			data[50482] <= 8'h10 ;
			data[50483] <= 8'h10 ;
			data[50484] <= 8'h10 ;
			data[50485] <= 8'h10 ;
			data[50486] <= 8'h10 ;
			data[50487] <= 8'h10 ;
			data[50488] <= 8'h10 ;
			data[50489] <= 8'h10 ;
			data[50490] <= 8'h10 ;
			data[50491] <= 8'h10 ;
			data[50492] <= 8'h10 ;
			data[50493] <= 8'h10 ;
			data[50494] <= 8'h10 ;
			data[50495] <= 8'h10 ;
			data[50496] <= 8'h10 ;
			data[50497] <= 8'h10 ;
			data[50498] <= 8'h10 ;
			data[50499] <= 8'h10 ;
			data[50500] <= 8'h10 ;
			data[50501] <= 8'h10 ;
			data[50502] <= 8'h10 ;
			data[50503] <= 8'h10 ;
			data[50504] <= 8'h10 ;
			data[50505] <= 8'h10 ;
			data[50506] <= 8'h10 ;
			data[50507] <= 8'h10 ;
			data[50508] <= 8'h10 ;
			data[50509] <= 8'h10 ;
			data[50510] <= 8'h10 ;
			data[50511] <= 8'h10 ;
			data[50512] <= 8'h10 ;
			data[50513] <= 8'h10 ;
			data[50514] <= 8'h10 ;
			data[50515] <= 8'h10 ;
			data[50516] <= 8'h10 ;
			data[50517] <= 8'h10 ;
			data[50518] <= 8'h10 ;
			data[50519] <= 8'h10 ;
			data[50520] <= 8'h10 ;
			data[50521] <= 8'h10 ;
			data[50522] <= 8'h10 ;
			data[50523] <= 8'h10 ;
			data[50524] <= 8'h10 ;
			data[50525] <= 8'h10 ;
			data[50526] <= 8'h10 ;
			data[50527] <= 8'h10 ;
			data[50528] <= 8'h10 ;
			data[50529] <= 8'h10 ;
			data[50530] <= 8'h10 ;
			data[50531] <= 8'h10 ;
			data[50532] <= 8'h10 ;
			data[50533] <= 8'h10 ;
			data[50534] <= 8'h10 ;
			data[50535] <= 8'h10 ;
			data[50536] <= 8'h10 ;
			data[50537] <= 8'h10 ;
			data[50538] <= 8'h10 ;
			data[50539] <= 8'h10 ;
			data[50540] <= 8'h10 ;
			data[50541] <= 8'h10 ;
			data[50542] <= 8'h10 ;
			data[50543] <= 8'h10 ;
			data[50544] <= 8'h10 ;
			data[50545] <= 8'h10 ;
			data[50546] <= 8'h10 ;
			data[50547] <= 8'h10 ;
			data[50548] <= 8'h10 ;
			data[50549] <= 8'h10 ;
			data[50550] <= 8'h10 ;
			data[50551] <= 8'h10 ;
			data[50552] <= 8'h10 ;
			data[50553] <= 8'h10 ;
			data[50554] <= 8'h10 ;
			data[50555] <= 8'h10 ;
			data[50556] <= 8'h10 ;
			data[50557] <= 8'h10 ;
			data[50558] <= 8'h10 ;
			data[50559] <= 8'h10 ;
			data[50560] <= 8'h10 ;
			data[50561] <= 8'h10 ;
			data[50562] <= 8'h10 ;
			data[50563] <= 8'h10 ;
			data[50564] <= 8'h10 ;
			data[50565] <= 8'h10 ;
			data[50566] <= 8'h10 ;
			data[50567] <= 8'h10 ;
			data[50568] <= 8'h10 ;
			data[50569] <= 8'h10 ;
			data[50570] <= 8'h10 ;
			data[50571] <= 8'h10 ;
			data[50572] <= 8'h10 ;
			data[50573] <= 8'h10 ;
			data[50574] <= 8'h10 ;
			data[50575] <= 8'h10 ;
			data[50576] <= 8'h10 ;
			data[50577] <= 8'h10 ;
			data[50578] <= 8'h10 ;
			data[50579] <= 8'h10 ;
			data[50580] <= 8'h10 ;
			data[50581] <= 8'h10 ;
			data[50582] <= 8'h10 ;
			data[50583] <= 8'h10 ;
			data[50584] <= 8'h10 ;
			data[50585] <= 8'h10 ;
			data[50586] <= 8'h10 ;
			data[50587] <= 8'h10 ;
			data[50588] <= 8'h10 ;
			data[50589] <= 8'h10 ;
			data[50590] <= 8'h10 ;
			data[50591] <= 8'h10 ;
			data[50592] <= 8'h10 ;
			data[50593] <= 8'h10 ;
			data[50594] <= 8'h10 ;
			data[50595] <= 8'h10 ;
			data[50596] <= 8'h10 ;
			data[50597] <= 8'h10 ;
			data[50598] <= 8'h10 ;
			data[50599] <= 8'h10 ;
			data[50600] <= 8'h10 ;
			data[50601] <= 8'h10 ;
			data[50602] <= 8'h10 ;
			data[50603] <= 8'h10 ;
			data[50604] <= 8'h10 ;
			data[50605] <= 8'h10 ;
			data[50606] <= 8'h10 ;
			data[50607] <= 8'h10 ;
			data[50608] <= 8'h10 ;
			data[50609] <= 8'h10 ;
			data[50610] <= 8'h10 ;
			data[50611] <= 8'h10 ;
			data[50612] <= 8'h10 ;
			data[50613] <= 8'h10 ;
			data[50614] <= 8'h10 ;
			data[50615] <= 8'h10 ;
			data[50616] <= 8'h10 ;
			data[50617] <= 8'h10 ;
			data[50618] <= 8'h10 ;
			data[50619] <= 8'h10 ;
			data[50620] <= 8'h10 ;
			data[50621] <= 8'h10 ;
			data[50622] <= 8'h10 ;
			data[50623] <= 8'h10 ;
			data[50624] <= 8'h10 ;
			data[50625] <= 8'h10 ;
			data[50626] <= 8'h10 ;
			data[50627] <= 8'h10 ;
			data[50628] <= 8'h10 ;
			data[50629] <= 8'h10 ;
			data[50630] <= 8'h10 ;
			data[50631] <= 8'h10 ;
			data[50632] <= 8'h10 ;
			data[50633] <= 8'h10 ;
			data[50634] <= 8'h10 ;
			data[50635] <= 8'h10 ;
			data[50636] <= 8'h10 ;
			data[50637] <= 8'h10 ;
			data[50638] <= 8'h10 ;
			data[50639] <= 8'h10 ;
			data[50640] <= 8'h10 ;
			data[50641] <= 8'h10 ;
			data[50642] <= 8'h10 ;
			data[50643] <= 8'h10 ;
			data[50644] <= 8'h10 ;
			data[50645] <= 8'h10 ;
			data[50646] <= 8'h10 ;
			data[50647] <= 8'h10 ;
			data[50648] <= 8'h10 ;
			data[50649] <= 8'h10 ;
			data[50650] <= 8'h10 ;
			data[50651] <= 8'h10 ;
			data[50652] <= 8'h10 ;
			data[50653] <= 8'h10 ;
			data[50654] <= 8'h10 ;
			data[50655] <= 8'h10 ;
			data[50656] <= 8'h10 ;
			data[50657] <= 8'h10 ;
			data[50658] <= 8'h10 ;
			data[50659] <= 8'h10 ;
			data[50660] <= 8'h10 ;
			data[50661] <= 8'h10 ;
			data[50662] <= 8'h10 ;
			data[50663] <= 8'h10 ;
			data[50664] <= 8'h10 ;
			data[50665] <= 8'h10 ;
			data[50666] <= 8'h10 ;
			data[50667] <= 8'h10 ;
			data[50668] <= 8'h10 ;
			data[50669] <= 8'h10 ;
			data[50670] <= 8'h10 ;
			data[50671] <= 8'h10 ;
			data[50672] <= 8'h10 ;
			data[50673] <= 8'h10 ;
			data[50674] <= 8'h10 ;
			data[50675] <= 8'h10 ;
			data[50676] <= 8'h10 ;
			data[50677] <= 8'h10 ;
			data[50678] <= 8'h10 ;
			data[50679] <= 8'h10 ;
			data[50680] <= 8'h10 ;
			data[50681] <= 8'h10 ;
			data[50682] <= 8'h10 ;
			data[50683] <= 8'h10 ;
			data[50684] <= 8'h10 ;
			data[50685] <= 8'h10 ;
			data[50686] <= 8'h10 ;
			data[50687] <= 8'h10 ;
			data[50688] <= 8'h10 ;
			data[50689] <= 8'h10 ;
			data[50690] <= 8'h10 ;
			data[50691] <= 8'h10 ;
			data[50692] <= 8'h10 ;
			data[50693] <= 8'h10 ;
			data[50694] <= 8'h10 ;
			data[50695] <= 8'h10 ;
			data[50696] <= 8'h10 ;
			data[50697] <= 8'h10 ;
			data[50698] <= 8'h10 ;
			data[50699] <= 8'h10 ;
			data[50700] <= 8'h10 ;
			data[50701] <= 8'h10 ;
			data[50702] <= 8'h10 ;
			data[50703] <= 8'h10 ;
			data[50704] <= 8'h10 ;
			data[50705] <= 8'h10 ;
			data[50706] <= 8'h10 ;
			data[50707] <= 8'h10 ;
			data[50708] <= 8'h10 ;
			data[50709] <= 8'h10 ;
			data[50710] <= 8'h10 ;
			data[50711] <= 8'h10 ;
			data[50712] <= 8'h10 ;
			data[50713] <= 8'h10 ;
			data[50714] <= 8'h10 ;
			data[50715] <= 8'h10 ;
			data[50716] <= 8'h10 ;
			data[50717] <= 8'h10 ;
			data[50718] <= 8'h10 ;
			data[50719] <= 8'h10 ;
			data[50720] <= 8'h10 ;
			data[50721] <= 8'h10 ;
			data[50722] <= 8'h10 ;
			data[50723] <= 8'h10 ;
			data[50724] <= 8'h10 ;
			data[50725] <= 8'h10 ;
			data[50726] <= 8'h10 ;
			data[50727] <= 8'h10 ;
			data[50728] <= 8'h10 ;
			data[50729] <= 8'h10 ;
			data[50730] <= 8'h10 ;
			data[50731] <= 8'h10 ;
			data[50732] <= 8'h10 ;
			data[50733] <= 8'h10 ;
			data[50734] <= 8'h10 ;
			data[50735] <= 8'h10 ;
			data[50736] <= 8'h10 ;
			data[50737] <= 8'h10 ;
			data[50738] <= 8'h10 ;
			data[50739] <= 8'h10 ;
			data[50740] <= 8'h10 ;
			data[50741] <= 8'h10 ;
			data[50742] <= 8'h10 ;
			data[50743] <= 8'h10 ;
			data[50744] <= 8'h10 ;
			data[50745] <= 8'h10 ;
			data[50746] <= 8'h10 ;
			data[50747] <= 8'h10 ;
			data[50748] <= 8'h10 ;
			data[50749] <= 8'h10 ;
			data[50750] <= 8'h10 ;
			data[50751] <= 8'h10 ;
			data[50752] <= 8'h10 ;
			data[50753] <= 8'h10 ;
			data[50754] <= 8'h10 ;
			data[50755] <= 8'h10 ;
			data[50756] <= 8'h10 ;
			data[50757] <= 8'h10 ;
			data[50758] <= 8'h10 ;
			data[50759] <= 8'h10 ;
			data[50760] <= 8'h10 ;
			data[50761] <= 8'h10 ;
			data[50762] <= 8'h10 ;
			data[50763] <= 8'h10 ;
			data[50764] <= 8'h10 ;
			data[50765] <= 8'h10 ;
			data[50766] <= 8'h10 ;
			data[50767] <= 8'h10 ;
			data[50768] <= 8'h10 ;
			data[50769] <= 8'h10 ;
			data[50770] <= 8'h10 ;
			data[50771] <= 8'h10 ;
			data[50772] <= 8'h10 ;
			data[50773] <= 8'h10 ;
			data[50774] <= 8'h10 ;
			data[50775] <= 8'h10 ;
			data[50776] <= 8'h10 ;
			data[50777] <= 8'h10 ;
			data[50778] <= 8'h10 ;
			data[50779] <= 8'h10 ;
			data[50780] <= 8'h10 ;
			data[50781] <= 8'h10 ;
			data[50782] <= 8'h10 ;
			data[50783] <= 8'h10 ;
			data[50784] <= 8'h10 ;
			data[50785] <= 8'h10 ;
			data[50786] <= 8'h10 ;
			data[50787] <= 8'h10 ;
			data[50788] <= 8'h10 ;
			data[50789] <= 8'h10 ;
			data[50790] <= 8'h10 ;
			data[50791] <= 8'h10 ;
			data[50792] <= 8'h10 ;
			data[50793] <= 8'h10 ;
			data[50794] <= 8'h10 ;
			data[50795] <= 8'h10 ;
			data[50796] <= 8'h10 ;
			data[50797] <= 8'h10 ;
			data[50798] <= 8'h10 ;
			data[50799] <= 8'h10 ;
			data[50800] <= 8'h10 ;
			data[50801] <= 8'h10 ;
			data[50802] <= 8'h10 ;
			data[50803] <= 8'h10 ;
			data[50804] <= 8'h10 ;
			data[50805] <= 8'h10 ;
			data[50806] <= 8'h10 ;
			data[50807] <= 8'h10 ;
			data[50808] <= 8'h10 ;
			data[50809] <= 8'h10 ;
			data[50810] <= 8'h10 ;
			data[50811] <= 8'h10 ;
			data[50812] <= 8'h10 ;
			data[50813] <= 8'h10 ;
			data[50814] <= 8'h10 ;
			data[50815] <= 8'h10 ;
			data[50816] <= 8'h10 ;
			data[50817] <= 8'h10 ;
			data[50818] <= 8'h10 ;
			data[50819] <= 8'h10 ;
			data[50820] <= 8'h10 ;
			data[50821] <= 8'h10 ;
			data[50822] <= 8'h10 ;
			data[50823] <= 8'h10 ;
			data[50824] <= 8'h10 ;
			data[50825] <= 8'h10 ;
			data[50826] <= 8'h10 ;
			data[50827] <= 8'h10 ;
			data[50828] <= 8'h10 ;
			data[50829] <= 8'h10 ;
			data[50830] <= 8'h10 ;
			data[50831] <= 8'h10 ;
			data[50832] <= 8'h10 ;
			data[50833] <= 8'h10 ;
			data[50834] <= 8'h10 ;
			data[50835] <= 8'h10 ;
			data[50836] <= 8'h10 ;
			data[50837] <= 8'h10 ;
			data[50838] <= 8'h10 ;
			data[50839] <= 8'h10 ;
			data[50840] <= 8'h10 ;
			data[50841] <= 8'h10 ;
			data[50842] <= 8'h10 ;
			data[50843] <= 8'h10 ;
			data[50844] <= 8'h10 ;
			data[50845] <= 8'h10 ;
			data[50846] <= 8'h10 ;
			data[50847] <= 8'h10 ;
			data[50848] <= 8'h10 ;
			data[50849] <= 8'h10 ;
			data[50850] <= 8'h10 ;
			data[50851] <= 8'h10 ;
			data[50852] <= 8'h10 ;
			data[50853] <= 8'h10 ;
			data[50854] <= 8'h10 ;
			data[50855] <= 8'h10 ;
			data[50856] <= 8'h10 ;
			data[50857] <= 8'h10 ;
			data[50858] <= 8'h10 ;
			data[50859] <= 8'h10 ;
			data[50860] <= 8'h10 ;
			data[50861] <= 8'h10 ;
			data[50862] <= 8'h10 ;
			data[50863] <= 8'h10 ;
			data[50864] <= 8'h10 ;
			data[50865] <= 8'h10 ;
			data[50866] <= 8'h10 ;
			data[50867] <= 8'h10 ;
			data[50868] <= 8'h10 ;
			data[50869] <= 8'h10 ;
			data[50870] <= 8'h10 ;
			data[50871] <= 8'h10 ;
			data[50872] <= 8'h10 ;
			data[50873] <= 8'h10 ;
			data[50874] <= 8'h10 ;
			data[50875] <= 8'h10 ;
			data[50876] <= 8'h10 ;
			data[50877] <= 8'h10 ;
			data[50878] <= 8'h10 ;
			data[50879] <= 8'h10 ;
			data[50880] <= 8'h10 ;
			data[50881] <= 8'h10 ;
			data[50882] <= 8'h10 ;
			data[50883] <= 8'h10 ;
			data[50884] <= 8'h10 ;
			data[50885] <= 8'h10 ;
			data[50886] <= 8'h10 ;
			data[50887] <= 8'h10 ;
			data[50888] <= 8'h10 ;
			data[50889] <= 8'h10 ;
			data[50890] <= 8'h10 ;
			data[50891] <= 8'h10 ;
			data[50892] <= 8'h10 ;
			data[50893] <= 8'h10 ;
			data[50894] <= 8'h10 ;
			data[50895] <= 8'h10 ;
			data[50896] <= 8'h10 ;
			data[50897] <= 8'h10 ;
			data[50898] <= 8'h10 ;
			data[50899] <= 8'h10 ;
			data[50900] <= 8'h10 ;
			data[50901] <= 8'h10 ;
			data[50902] <= 8'h10 ;
			data[50903] <= 8'h10 ;
			data[50904] <= 8'h10 ;
			data[50905] <= 8'h10 ;
			data[50906] <= 8'h10 ;
			data[50907] <= 8'h10 ;
			data[50908] <= 8'h10 ;
			data[50909] <= 8'h10 ;
			data[50910] <= 8'h10 ;
			data[50911] <= 8'h10 ;
			data[50912] <= 8'h10 ;
			data[50913] <= 8'h10 ;
			data[50914] <= 8'h10 ;
			data[50915] <= 8'h10 ;
			data[50916] <= 8'h10 ;
			data[50917] <= 8'h10 ;
			data[50918] <= 8'h10 ;
			data[50919] <= 8'h10 ;
			data[50920] <= 8'h10 ;
			data[50921] <= 8'h10 ;
			data[50922] <= 8'h10 ;
			data[50923] <= 8'h10 ;
			data[50924] <= 8'h10 ;
			data[50925] <= 8'h10 ;
			data[50926] <= 8'h10 ;
			data[50927] <= 8'h10 ;
			data[50928] <= 8'h10 ;
			data[50929] <= 8'h10 ;
			data[50930] <= 8'h10 ;
			data[50931] <= 8'h10 ;
			data[50932] <= 8'h10 ;
			data[50933] <= 8'h10 ;
			data[50934] <= 8'h10 ;
			data[50935] <= 8'h10 ;
			data[50936] <= 8'h10 ;
			data[50937] <= 8'h10 ;
			data[50938] <= 8'h10 ;
			data[50939] <= 8'h10 ;
			data[50940] <= 8'h10 ;
			data[50941] <= 8'h10 ;
			data[50942] <= 8'h10 ;
			data[50943] <= 8'h10 ;
			data[50944] <= 8'h10 ;
			data[50945] <= 8'h10 ;
			data[50946] <= 8'h10 ;
			data[50947] <= 8'h10 ;
			data[50948] <= 8'h10 ;
			data[50949] <= 8'h10 ;
			data[50950] <= 8'h10 ;
			data[50951] <= 8'h10 ;
			data[50952] <= 8'h10 ;
			data[50953] <= 8'h10 ;
			data[50954] <= 8'h10 ;
			data[50955] <= 8'h10 ;
			data[50956] <= 8'h10 ;
			data[50957] <= 8'h10 ;
			data[50958] <= 8'h10 ;
			data[50959] <= 8'h10 ;
			data[50960] <= 8'h10 ;
			data[50961] <= 8'h10 ;
			data[50962] <= 8'h10 ;
			data[50963] <= 8'h10 ;
			data[50964] <= 8'h10 ;
			data[50965] <= 8'h10 ;
			data[50966] <= 8'h10 ;
			data[50967] <= 8'h10 ;
			data[50968] <= 8'h10 ;
			data[50969] <= 8'h10 ;
			data[50970] <= 8'h10 ;
			data[50971] <= 8'h10 ;
			data[50972] <= 8'h10 ;
			data[50973] <= 8'h10 ;
			data[50974] <= 8'h10 ;
			data[50975] <= 8'h10 ;
			data[50976] <= 8'h10 ;
			data[50977] <= 8'h10 ;
			data[50978] <= 8'h10 ;
			data[50979] <= 8'h10 ;
			data[50980] <= 8'h10 ;
			data[50981] <= 8'h10 ;
			data[50982] <= 8'h10 ;
			data[50983] <= 8'h10 ;
			data[50984] <= 8'h10 ;
			data[50985] <= 8'h10 ;
			data[50986] <= 8'h10 ;
			data[50987] <= 8'h10 ;
			data[50988] <= 8'h10 ;
			data[50989] <= 8'h10 ;
			data[50990] <= 8'h10 ;
			data[50991] <= 8'h10 ;
			data[50992] <= 8'h10 ;
			data[50993] <= 8'h10 ;
			data[50994] <= 8'h10 ;
			data[50995] <= 8'h10 ;
			data[50996] <= 8'h10 ;
			data[50997] <= 8'h10 ;
			data[50998] <= 8'h10 ;
			data[50999] <= 8'h10 ;
			data[51000] <= 8'h10 ;
			data[51001] <= 8'h10 ;
			data[51002] <= 8'h10 ;
			data[51003] <= 8'h10 ;
			data[51004] <= 8'h10 ;
			data[51005] <= 8'h10 ;
			data[51006] <= 8'h10 ;
			data[51007] <= 8'h10 ;
			data[51008] <= 8'h10 ;
			data[51009] <= 8'h10 ;
			data[51010] <= 8'h10 ;
			data[51011] <= 8'h10 ;
			data[51012] <= 8'h10 ;
			data[51013] <= 8'h10 ;
			data[51014] <= 8'h10 ;
			data[51015] <= 8'h10 ;
			data[51016] <= 8'h10 ;
			data[51017] <= 8'h10 ;
			data[51018] <= 8'h10 ;
			data[51019] <= 8'h10 ;
			data[51020] <= 8'h10 ;
			data[51021] <= 8'h10 ;
			data[51022] <= 8'h10 ;
			data[51023] <= 8'h10 ;
			data[51024] <= 8'h10 ;
			data[51025] <= 8'h10 ;
			data[51026] <= 8'h10 ;
			data[51027] <= 8'h10 ;
			data[51028] <= 8'h10 ;
			data[51029] <= 8'h10 ;
			data[51030] <= 8'h10 ;
			data[51031] <= 8'h10 ;
			data[51032] <= 8'h10 ;
			data[51033] <= 8'h10 ;
			data[51034] <= 8'h10 ;
			data[51035] <= 8'h10 ;
			data[51036] <= 8'h10 ;
			data[51037] <= 8'h10 ;
			data[51038] <= 8'h10 ;
			data[51039] <= 8'h10 ;
			data[51040] <= 8'h10 ;
			data[51041] <= 8'h10 ;
			data[51042] <= 8'h10 ;
			data[51043] <= 8'h10 ;
			data[51044] <= 8'h10 ;
			data[51045] <= 8'h10 ;
			data[51046] <= 8'h10 ;
			data[51047] <= 8'h10 ;
			data[51048] <= 8'h10 ;
			data[51049] <= 8'h10 ;
			data[51050] <= 8'h10 ;
			data[51051] <= 8'h10 ;
			data[51052] <= 8'h10 ;
			data[51053] <= 8'h10 ;
			data[51054] <= 8'h10 ;
			data[51055] <= 8'h10 ;
			data[51056] <= 8'h10 ;
			data[51057] <= 8'h10 ;
			data[51058] <= 8'h10 ;
			data[51059] <= 8'h10 ;
			data[51060] <= 8'h10 ;
			data[51061] <= 8'h10 ;
			data[51062] <= 8'h10 ;
			data[51063] <= 8'h10 ;
			data[51064] <= 8'h10 ;
			data[51065] <= 8'h10 ;
			data[51066] <= 8'h10 ;
			data[51067] <= 8'h10 ;
			data[51068] <= 8'h10 ;
			data[51069] <= 8'h10 ;
			data[51070] <= 8'h10 ;
			data[51071] <= 8'h10 ;
			data[51072] <= 8'h10 ;
			data[51073] <= 8'h10 ;
			data[51074] <= 8'h10 ;
			data[51075] <= 8'h10 ;
			data[51076] <= 8'h10 ;
			data[51077] <= 8'h10 ;
			data[51078] <= 8'h10 ;
			data[51079] <= 8'h10 ;
			data[51080] <= 8'h10 ;
			data[51081] <= 8'h10 ;
			data[51082] <= 8'h10 ;
			data[51083] <= 8'h10 ;
			data[51084] <= 8'h10 ;
			data[51085] <= 8'h10 ;
			data[51086] <= 8'h10 ;
			data[51087] <= 8'h10 ;
			data[51088] <= 8'h10 ;
			data[51089] <= 8'h10 ;
			data[51090] <= 8'h10 ;
			data[51091] <= 8'h10 ;
			data[51092] <= 8'h10 ;
			data[51093] <= 8'h10 ;
			data[51094] <= 8'h10 ;
			data[51095] <= 8'h10 ;
			data[51096] <= 8'h10 ;
			data[51097] <= 8'h10 ;
			data[51098] <= 8'h10 ;
			data[51099] <= 8'h10 ;
			data[51100] <= 8'h10 ;
			data[51101] <= 8'h10 ;
			data[51102] <= 8'h10 ;
			data[51103] <= 8'h10 ;
			data[51104] <= 8'h10 ;
			data[51105] <= 8'h10 ;
			data[51106] <= 8'h10 ;
			data[51107] <= 8'h10 ;
			data[51108] <= 8'h10 ;
			data[51109] <= 8'h10 ;
			data[51110] <= 8'h10 ;
			data[51111] <= 8'h10 ;
			data[51112] <= 8'h10 ;
			data[51113] <= 8'h10 ;
			data[51114] <= 8'h10 ;
			data[51115] <= 8'h10 ;
			data[51116] <= 8'h10 ;
			data[51117] <= 8'h10 ;
			data[51118] <= 8'h10 ;
			data[51119] <= 8'h10 ;
			data[51120] <= 8'h10 ;
			data[51121] <= 8'h10 ;
			data[51122] <= 8'h10 ;
			data[51123] <= 8'h10 ;
			data[51124] <= 8'h10 ;
			data[51125] <= 8'h10 ;
			data[51126] <= 8'h10 ;
			data[51127] <= 8'h10 ;
			data[51128] <= 8'h10 ;
			data[51129] <= 8'h10 ;
			data[51130] <= 8'h10 ;
			data[51131] <= 8'h10 ;
			data[51132] <= 8'h10 ;
			data[51133] <= 8'h10 ;
			data[51134] <= 8'h10 ;
			data[51135] <= 8'h10 ;
			data[51136] <= 8'h10 ;
			data[51137] <= 8'h10 ;
			data[51138] <= 8'h10 ;
			data[51139] <= 8'h10 ;
			data[51140] <= 8'h10 ;
			data[51141] <= 8'h10 ;
			data[51142] <= 8'h10 ;
			data[51143] <= 8'h10 ;
			data[51144] <= 8'h10 ;
			data[51145] <= 8'h10 ;
			data[51146] <= 8'h10 ;
			data[51147] <= 8'h10 ;
			data[51148] <= 8'h10 ;
			data[51149] <= 8'h10 ;
			data[51150] <= 8'h10 ;
			data[51151] <= 8'h10 ;
			data[51152] <= 8'h10 ;
			data[51153] <= 8'h10 ;
			data[51154] <= 8'h10 ;
			data[51155] <= 8'h10 ;
			data[51156] <= 8'h10 ;
			data[51157] <= 8'h10 ;
			data[51158] <= 8'h10 ;
			data[51159] <= 8'h10 ;
			data[51160] <= 8'h10 ;
			data[51161] <= 8'h10 ;
			data[51162] <= 8'h10 ;
			data[51163] <= 8'h10 ;
			data[51164] <= 8'h10 ;
			data[51165] <= 8'h10 ;
			data[51166] <= 8'h10 ;
			data[51167] <= 8'h10 ;
			data[51168] <= 8'h10 ;
			data[51169] <= 8'h10 ;
			data[51170] <= 8'h10 ;
			data[51171] <= 8'h10 ;
			data[51172] <= 8'h10 ;
			data[51173] <= 8'h10 ;
			data[51174] <= 8'h10 ;
			data[51175] <= 8'h10 ;
			data[51176] <= 8'h10 ;
			data[51177] <= 8'h10 ;
			data[51178] <= 8'h10 ;
			data[51179] <= 8'h10 ;
			data[51180] <= 8'h10 ;
			data[51181] <= 8'h10 ;
			data[51182] <= 8'h10 ;
			data[51183] <= 8'h10 ;
			data[51184] <= 8'h10 ;
			data[51185] <= 8'h10 ;
			data[51186] <= 8'h10 ;
			data[51187] <= 8'h10 ;
			data[51188] <= 8'h10 ;
			data[51189] <= 8'h10 ;
			data[51190] <= 8'h10 ;
			data[51191] <= 8'h10 ;
			data[51192] <= 8'h10 ;
			data[51193] <= 8'h10 ;
			data[51194] <= 8'h10 ;
			data[51195] <= 8'h10 ;
			data[51196] <= 8'h10 ;
			data[51197] <= 8'h10 ;
			data[51198] <= 8'h10 ;
			data[51199] <= 8'h10 ;
			data[51200] <= 8'h10 ;
			data[51201] <= 8'h10 ;
			data[51202] <= 8'h10 ;
			data[51203] <= 8'h10 ;
			data[51204] <= 8'h10 ;
			data[51205] <= 8'h10 ;
			data[51206] <= 8'h10 ;
			data[51207] <= 8'h10 ;
			data[51208] <= 8'h10 ;
			data[51209] <= 8'h10 ;
			data[51210] <= 8'h10 ;
			data[51211] <= 8'h10 ;
			data[51212] <= 8'h10 ;
			data[51213] <= 8'h10 ;
			data[51214] <= 8'h10 ;
			data[51215] <= 8'h10 ;
			data[51216] <= 8'h10 ;
			data[51217] <= 8'h10 ;
			data[51218] <= 8'h10 ;
			data[51219] <= 8'h10 ;
			data[51220] <= 8'h10 ;
			data[51221] <= 8'h10 ;
			data[51222] <= 8'h10 ;
			data[51223] <= 8'h10 ;
			data[51224] <= 8'h10 ;
			data[51225] <= 8'h10 ;
			data[51226] <= 8'h10 ;
			data[51227] <= 8'h10 ;
			data[51228] <= 8'h10 ;
			data[51229] <= 8'h10 ;
			data[51230] <= 8'h10 ;
			data[51231] <= 8'h10 ;
			data[51232] <= 8'h10 ;
			data[51233] <= 8'h10 ;
			data[51234] <= 8'h10 ;
			data[51235] <= 8'h10 ;
			data[51236] <= 8'h10 ;
			data[51237] <= 8'h10 ;
			data[51238] <= 8'h10 ;
			data[51239] <= 8'h10 ;
			data[51240] <= 8'h10 ;
			data[51241] <= 8'h10 ;
			data[51242] <= 8'h10 ;
			data[51243] <= 8'h10 ;
			data[51244] <= 8'h10 ;
			data[51245] <= 8'h10 ;
			data[51246] <= 8'h10 ;
			data[51247] <= 8'h10 ;
			data[51248] <= 8'h10 ;
			data[51249] <= 8'h10 ;
			data[51250] <= 8'h10 ;
			data[51251] <= 8'h10 ;
			data[51252] <= 8'h10 ;
			data[51253] <= 8'h10 ;
			data[51254] <= 8'h10 ;
			data[51255] <= 8'h10 ;
			data[51256] <= 8'h10 ;
			data[51257] <= 8'h10 ;
			data[51258] <= 8'h10 ;
			data[51259] <= 8'h10 ;
			data[51260] <= 8'h10 ;
			data[51261] <= 8'h10 ;
			data[51262] <= 8'h10 ;
			data[51263] <= 8'h10 ;
			data[51264] <= 8'h10 ;
			data[51265] <= 8'h10 ;
			data[51266] <= 8'h10 ;
			data[51267] <= 8'h10 ;
			data[51268] <= 8'h10 ;
			data[51269] <= 8'h10 ;
			data[51270] <= 8'h10 ;
			data[51271] <= 8'h10 ;
			data[51272] <= 8'h10 ;
			data[51273] <= 8'h10 ;
			data[51274] <= 8'h10 ;
			data[51275] <= 8'h10 ;
			data[51276] <= 8'h10 ;
			data[51277] <= 8'h10 ;
			data[51278] <= 8'h10 ;
			data[51279] <= 8'h10 ;
			data[51280] <= 8'h10 ;
			data[51281] <= 8'h10 ;
			data[51282] <= 8'h10 ;
			data[51283] <= 8'h10 ;
			data[51284] <= 8'h10 ;
			data[51285] <= 8'h10 ;
			data[51286] <= 8'h10 ;
			data[51287] <= 8'h10 ;
			data[51288] <= 8'h10 ;
			data[51289] <= 8'h10 ;
			data[51290] <= 8'h10 ;
			data[51291] <= 8'h10 ;
			data[51292] <= 8'h10 ;
			data[51293] <= 8'h10 ;
			data[51294] <= 8'h10 ;
			data[51295] <= 8'h10 ;
			data[51296] <= 8'h10 ;
			data[51297] <= 8'h10 ;
			data[51298] <= 8'h10 ;
			data[51299] <= 8'h10 ;
			data[51300] <= 8'h10 ;
			data[51301] <= 8'h10 ;
			data[51302] <= 8'h10 ;
			data[51303] <= 8'h10 ;
			data[51304] <= 8'h10 ;
			data[51305] <= 8'h10 ;
			data[51306] <= 8'h10 ;
			data[51307] <= 8'h10 ;
			data[51308] <= 8'h10 ;
			data[51309] <= 8'h10 ;
			data[51310] <= 8'h10 ;
			data[51311] <= 8'h10 ;
			data[51312] <= 8'h10 ;
			data[51313] <= 8'h10 ;
			data[51314] <= 8'h10 ;
			data[51315] <= 8'h10 ;
			data[51316] <= 8'h10 ;
			data[51317] <= 8'h10 ;
			data[51318] <= 8'h10 ;
			data[51319] <= 8'h10 ;
			data[51320] <= 8'h10 ;
			data[51321] <= 8'h10 ;
			data[51322] <= 8'h10 ;
			data[51323] <= 8'h10 ;
			data[51324] <= 8'h10 ;
			data[51325] <= 8'h10 ;
			data[51326] <= 8'h10 ;
			data[51327] <= 8'h10 ;
			data[51328] <= 8'h10 ;
			data[51329] <= 8'h10 ;
			data[51330] <= 8'h10 ;
			data[51331] <= 8'h10 ;
			data[51332] <= 8'h10 ;
			data[51333] <= 8'h10 ;
			data[51334] <= 8'h10 ;
			data[51335] <= 8'h10 ;
			data[51336] <= 8'h10 ;
			data[51337] <= 8'h10 ;
			data[51338] <= 8'h10 ;
			data[51339] <= 8'h10 ;
			data[51340] <= 8'h10 ;
			data[51341] <= 8'h10 ;
			data[51342] <= 8'h10 ;
			data[51343] <= 8'h10 ;
			data[51344] <= 8'h10 ;
			data[51345] <= 8'h10 ;
			data[51346] <= 8'h10 ;
			data[51347] <= 8'h10 ;
			data[51348] <= 8'h10 ;
			data[51349] <= 8'h10 ;
			data[51350] <= 8'h10 ;
			data[51351] <= 8'h10 ;
			data[51352] <= 8'h10 ;
			data[51353] <= 8'h10 ;
			data[51354] <= 8'h10 ;
			data[51355] <= 8'h10 ;
			data[51356] <= 8'h10 ;
			data[51357] <= 8'h10 ;
			data[51358] <= 8'h10 ;
			data[51359] <= 8'h10 ;
			data[51360] <= 8'h10 ;
			data[51361] <= 8'h10 ;
			data[51362] <= 8'h10 ;
			data[51363] <= 8'h10 ;
			data[51364] <= 8'h10 ;
			data[51365] <= 8'h10 ;
			data[51366] <= 8'h10 ;
			data[51367] <= 8'h10 ;
			data[51368] <= 8'h10 ;
			data[51369] <= 8'h10 ;
			data[51370] <= 8'h10 ;
			data[51371] <= 8'h10 ;
			data[51372] <= 8'h10 ;
			data[51373] <= 8'h10 ;
			data[51374] <= 8'h10 ;
			data[51375] <= 8'h10 ;
			data[51376] <= 8'h10 ;
			data[51377] <= 8'h10 ;
			data[51378] <= 8'h10 ;
			data[51379] <= 8'h10 ;
			data[51380] <= 8'h10 ;
			data[51381] <= 8'h10 ;
			data[51382] <= 8'h10 ;
			data[51383] <= 8'h10 ;
			data[51384] <= 8'h10 ;
			data[51385] <= 8'h10 ;
			data[51386] <= 8'h10 ;
			data[51387] <= 8'h10 ;
			data[51388] <= 8'h10 ;
			data[51389] <= 8'h10 ;
			data[51390] <= 8'h10 ;
			data[51391] <= 8'h10 ;
			data[51392] <= 8'h10 ;
			data[51393] <= 8'h10 ;
			data[51394] <= 8'h10 ;
			data[51395] <= 8'h10 ;
			data[51396] <= 8'h10 ;
			data[51397] <= 8'h10 ;
			data[51398] <= 8'h10 ;
			data[51399] <= 8'h10 ;
			data[51400] <= 8'h10 ;
			data[51401] <= 8'h10 ;
			data[51402] <= 8'h10 ;
			data[51403] <= 8'h10 ;
			data[51404] <= 8'h10 ;
			data[51405] <= 8'h10 ;
			data[51406] <= 8'h10 ;
			data[51407] <= 8'h10 ;
			data[51408] <= 8'h10 ;
			data[51409] <= 8'h10 ;
			data[51410] <= 8'h10 ;
			data[51411] <= 8'h10 ;
			data[51412] <= 8'h10 ;
			data[51413] <= 8'h10 ;
			data[51414] <= 8'h10 ;
			data[51415] <= 8'h10 ;
			data[51416] <= 8'h10 ;
			data[51417] <= 8'h10 ;
			data[51418] <= 8'h10 ;
			data[51419] <= 8'h10 ;
			data[51420] <= 8'h10 ;
			data[51421] <= 8'h10 ;
			data[51422] <= 8'h10 ;
			data[51423] <= 8'h10 ;
			data[51424] <= 8'h10 ;
			data[51425] <= 8'h10 ;
			data[51426] <= 8'h10 ;
			data[51427] <= 8'h10 ;
			data[51428] <= 8'h10 ;
			data[51429] <= 8'h10 ;
			data[51430] <= 8'h10 ;
			data[51431] <= 8'h10 ;
			data[51432] <= 8'h10 ;
			data[51433] <= 8'h10 ;
			data[51434] <= 8'h10 ;
			data[51435] <= 8'h10 ;
			data[51436] <= 8'h10 ;
			data[51437] <= 8'h10 ;
			data[51438] <= 8'h10 ;
			data[51439] <= 8'h10 ;
			data[51440] <= 8'h10 ;
			data[51441] <= 8'h10 ;
			data[51442] <= 8'h10 ;
			data[51443] <= 8'h10 ;
			data[51444] <= 8'h10 ;
			data[51445] <= 8'h10 ;
			data[51446] <= 8'h10 ;
			data[51447] <= 8'h10 ;
			data[51448] <= 8'h10 ;
			data[51449] <= 8'h10 ;
			data[51450] <= 8'h10 ;
			data[51451] <= 8'h10 ;
			data[51452] <= 8'h10 ;
			data[51453] <= 8'h10 ;
			data[51454] <= 8'h10 ;
			data[51455] <= 8'h10 ;
			data[51456] <= 8'h10 ;
			data[51457] <= 8'h10 ;
			data[51458] <= 8'h10 ;
			data[51459] <= 8'h10 ;
			data[51460] <= 8'h10 ;
			data[51461] <= 8'h10 ;
			data[51462] <= 8'h10 ;
			data[51463] <= 8'h10 ;
			data[51464] <= 8'h10 ;
			data[51465] <= 8'h10 ;
			data[51466] <= 8'h10 ;
			data[51467] <= 8'h10 ;
			data[51468] <= 8'h10 ;
			data[51469] <= 8'h10 ;
			data[51470] <= 8'h10 ;
			data[51471] <= 8'h10 ;
			data[51472] <= 8'h10 ;
			data[51473] <= 8'h10 ;
			data[51474] <= 8'h10 ;
			data[51475] <= 8'h10 ;
			data[51476] <= 8'h10 ;
			data[51477] <= 8'h10 ;
			data[51478] <= 8'h10 ;
			data[51479] <= 8'h10 ;
			data[51480] <= 8'h10 ;
			data[51481] <= 8'h10 ;
			data[51482] <= 8'h10 ;
			data[51483] <= 8'h10 ;
			data[51484] <= 8'h10 ;
			data[51485] <= 8'h10 ;
			data[51486] <= 8'h10 ;
			data[51487] <= 8'h10 ;
			data[51488] <= 8'h10 ;
			data[51489] <= 8'h10 ;
			data[51490] <= 8'h10 ;
			data[51491] <= 8'h10 ;
			data[51492] <= 8'h10 ;
			data[51493] <= 8'h10 ;
			data[51494] <= 8'h10 ;
			data[51495] <= 8'h10 ;
			data[51496] <= 8'h10 ;
			data[51497] <= 8'h10 ;
			data[51498] <= 8'h10 ;
			data[51499] <= 8'h10 ;
			data[51500] <= 8'h10 ;
			data[51501] <= 8'h10 ;
			data[51502] <= 8'h10 ;
			data[51503] <= 8'h10 ;
			data[51504] <= 8'h10 ;
			data[51505] <= 8'h10 ;
			data[51506] <= 8'h10 ;
			data[51507] <= 8'h10 ;
			data[51508] <= 8'h10 ;
			data[51509] <= 8'h10 ;
			data[51510] <= 8'h10 ;
			data[51511] <= 8'h10 ;
			data[51512] <= 8'h10 ;
			data[51513] <= 8'h10 ;
			data[51514] <= 8'h10 ;
			data[51515] <= 8'h10 ;
			data[51516] <= 8'h10 ;
			data[51517] <= 8'h10 ;
			data[51518] <= 8'h10 ;
			data[51519] <= 8'h10 ;
			data[51520] <= 8'h10 ;
			data[51521] <= 8'h10 ;
			data[51522] <= 8'h10 ;
			data[51523] <= 8'h10 ;
			data[51524] <= 8'h10 ;
			data[51525] <= 8'h10 ;
			data[51526] <= 8'h10 ;
			data[51527] <= 8'h10 ;
			data[51528] <= 8'h10 ;
			data[51529] <= 8'h10 ;
			data[51530] <= 8'h10 ;
			data[51531] <= 8'h10 ;
			data[51532] <= 8'h10 ;
			data[51533] <= 8'h10 ;
			data[51534] <= 8'h10 ;
			data[51535] <= 8'h10 ;
			data[51536] <= 8'h10 ;
			data[51537] <= 8'h10 ;
			data[51538] <= 8'h10 ;
			data[51539] <= 8'h10 ;
			data[51540] <= 8'h10 ;
			data[51541] <= 8'h10 ;
			data[51542] <= 8'h10 ;
			data[51543] <= 8'h10 ;
			data[51544] <= 8'h10 ;
			data[51545] <= 8'h10 ;
			data[51546] <= 8'h10 ;
			data[51547] <= 8'h10 ;
			data[51548] <= 8'h10 ;
			data[51549] <= 8'h10 ;
			data[51550] <= 8'h10 ;
			data[51551] <= 8'h10 ;
			data[51552] <= 8'h10 ;
			data[51553] <= 8'h10 ;
			data[51554] <= 8'h10 ;
			data[51555] <= 8'h10 ;
			data[51556] <= 8'h10 ;
			data[51557] <= 8'h10 ;
			data[51558] <= 8'h10 ;
			data[51559] <= 8'h10 ;
			data[51560] <= 8'h10 ;
			data[51561] <= 8'h10 ;
			data[51562] <= 8'h10 ;
			data[51563] <= 8'h10 ;
			data[51564] <= 8'h10 ;
			data[51565] <= 8'h10 ;
			data[51566] <= 8'h10 ;
			data[51567] <= 8'h10 ;
			data[51568] <= 8'h10 ;
			data[51569] <= 8'h10 ;
			data[51570] <= 8'h10 ;
			data[51571] <= 8'h10 ;
			data[51572] <= 8'h10 ;
			data[51573] <= 8'h10 ;
			data[51574] <= 8'h10 ;
			data[51575] <= 8'h10 ;
			data[51576] <= 8'h10 ;
			data[51577] <= 8'h10 ;
			data[51578] <= 8'h10 ;
			data[51579] <= 8'h10 ;
			data[51580] <= 8'h10 ;
			data[51581] <= 8'h10 ;
			data[51582] <= 8'h10 ;
			data[51583] <= 8'h10 ;
			data[51584] <= 8'h10 ;
			data[51585] <= 8'h10 ;
			data[51586] <= 8'h10 ;
			data[51587] <= 8'h10 ;
			data[51588] <= 8'h10 ;
			data[51589] <= 8'h10 ;
			data[51590] <= 8'h10 ;
			data[51591] <= 8'h10 ;
			data[51592] <= 8'h10 ;
			data[51593] <= 8'h10 ;
			data[51594] <= 8'h10 ;
			data[51595] <= 8'h10 ;
			data[51596] <= 8'h10 ;
			data[51597] <= 8'h10 ;
			data[51598] <= 8'h10 ;
			data[51599] <= 8'h10 ;
			data[51600] <= 8'h10 ;
			data[51601] <= 8'h10 ;
			data[51602] <= 8'h10 ;
			data[51603] <= 8'h10 ;
			data[51604] <= 8'h10 ;
			data[51605] <= 8'h10 ;
			data[51606] <= 8'h10 ;
			data[51607] <= 8'h10 ;
			data[51608] <= 8'h10 ;
			data[51609] <= 8'h10 ;
			data[51610] <= 8'h10 ;
			data[51611] <= 8'h10 ;
			data[51612] <= 8'h10 ;
			data[51613] <= 8'h10 ;
			data[51614] <= 8'h10 ;
			data[51615] <= 8'h10 ;
			data[51616] <= 8'h10 ;
			data[51617] <= 8'h10 ;
			data[51618] <= 8'h10 ;
			data[51619] <= 8'h10 ;
			data[51620] <= 8'h10 ;
			data[51621] <= 8'h10 ;
			data[51622] <= 8'h10 ;
			data[51623] <= 8'h10 ;
			data[51624] <= 8'h10 ;
			data[51625] <= 8'h10 ;
			data[51626] <= 8'h10 ;
			data[51627] <= 8'h10 ;
			data[51628] <= 8'h10 ;
			data[51629] <= 8'h10 ;
			data[51630] <= 8'h10 ;
			data[51631] <= 8'h10 ;
			data[51632] <= 8'h10 ;
			data[51633] <= 8'h10 ;
			data[51634] <= 8'h10 ;
			data[51635] <= 8'h10 ;
			data[51636] <= 8'h10 ;
			data[51637] <= 8'h10 ;
			data[51638] <= 8'h10 ;
			data[51639] <= 8'h10 ;
			data[51640] <= 8'h10 ;
			data[51641] <= 8'h10 ;
			data[51642] <= 8'h10 ;
			data[51643] <= 8'h10 ;
			data[51644] <= 8'h10 ;
			data[51645] <= 8'h10 ;
			data[51646] <= 8'h10 ;
			data[51647] <= 8'h10 ;
			data[51648] <= 8'h10 ;
			data[51649] <= 8'h10 ;
			data[51650] <= 8'h10 ;
			data[51651] <= 8'h10 ;
			data[51652] <= 8'h10 ;
			data[51653] <= 8'h10 ;
			data[51654] <= 8'h10 ;
			data[51655] <= 8'h10 ;
			data[51656] <= 8'h10 ;
			data[51657] <= 8'h10 ;
			data[51658] <= 8'h10 ;
			data[51659] <= 8'h10 ;
			data[51660] <= 8'h10 ;
			data[51661] <= 8'h10 ;
			data[51662] <= 8'h10 ;
			data[51663] <= 8'h10 ;
			data[51664] <= 8'h10 ;
			data[51665] <= 8'h10 ;
			data[51666] <= 8'h10 ;
			data[51667] <= 8'h10 ;
			data[51668] <= 8'h10 ;
			data[51669] <= 8'h10 ;
			data[51670] <= 8'h10 ;
			data[51671] <= 8'h10 ;
			data[51672] <= 8'h10 ;
			data[51673] <= 8'h10 ;
			data[51674] <= 8'h10 ;
			data[51675] <= 8'h10 ;
			data[51676] <= 8'h10 ;
			data[51677] <= 8'h10 ;
			data[51678] <= 8'h10 ;
			data[51679] <= 8'h10 ;
			data[51680] <= 8'h10 ;
			data[51681] <= 8'h10 ;
			data[51682] <= 8'h10 ;
			data[51683] <= 8'h10 ;
			data[51684] <= 8'h10 ;
			data[51685] <= 8'h10 ;
			data[51686] <= 8'h10 ;
			data[51687] <= 8'h10 ;
			data[51688] <= 8'h10 ;
			data[51689] <= 8'h10 ;
			data[51690] <= 8'h10 ;
			data[51691] <= 8'h10 ;
			data[51692] <= 8'h10 ;
			data[51693] <= 8'h10 ;
			data[51694] <= 8'h10 ;
			data[51695] <= 8'h10 ;
			data[51696] <= 8'h10 ;
			data[51697] <= 8'h10 ;
			data[51698] <= 8'h10 ;
			data[51699] <= 8'h10 ;
			data[51700] <= 8'h10 ;
			data[51701] <= 8'h10 ;
			data[51702] <= 8'h10 ;
			data[51703] <= 8'h10 ;
			data[51704] <= 8'h10 ;
			data[51705] <= 8'h10 ;
			data[51706] <= 8'h10 ;
			data[51707] <= 8'h10 ;
			data[51708] <= 8'h10 ;
			data[51709] <= 8'h10 ;
			data[51710] <= 8'h10 ;
			data[51711] <= 8'h10 ;
			data[51712] <= 8'h10 ;
			data[51713] <= 8'h10 ;
			data[51714] <= 8'h10 ;
			data[51715] <= 8'h10 ;
			data[51716] <= 8'h10 ;
			data[51717] <= 8'h10 ;
			data[51718] <= 8'h10 ;
			data[51719] <= 8'h10 ;
			data[51720] <= 8'h10 ;
			data[51721] <= 8'h10 ;
			data[51722] <= 8'h10 ;
			data[51723] <= 8'h10 ;
			data[51724] <= 8'h10 ;
			data[51725] <= 8'h10 ;
			data[51726] <= 8'h10 ;
			data[51727] <= 8'h10 ;
			data[51728] <= 8'h10 ;
			data[51729] <= 8'h10 ;
			data[51730] <= 8'h10 ;
			data[51731] <= 8'h10 ;
			data[51732] <= 8'h10 ;
			data[51733] <= 8'h10 ;
			data[51734] <= 8'h10 ;
			data[51735] <= 8'h10 ;
			data[51736] <= 8'h10 ;
			data[51737] <= 8'h10 ;
			data[51738] <= 8'h10 ;
			data[51739] <= 8'h10 ;
			data[51740] <= 8'h10 ;
			data[51741] <= 8'h10 ;
			data[51742] <= 8'h10 ;
			data[51743] <= 8'h10 ;
			data[51744] <= 8'h10 ;
			data[51745] <= 8'h10 ;
			data[51746] <= 8'h10 ;
			data[51747] <= 8'h10 ;
			data[51748] <= 8'h10 ;
			data[51749] <= 8'h10 ;
			data[51750] <= 8'h10 ;
			data[51751] <= 8'h10 ;
			data[51752] <= 8'h10 ;
			data[51753] <= 8'h10 ;
			data[51754] <= 8'h10 ;
			data[51755] <= 8'h10 ;
			data[51756] <= 8'h10 ;
			data[51757] <= 8'h10 ;
			data[51758] <= 8'h10 ;
			data[51759] <= 8'h10 ;
			data[51760] <= 8'h10 ;
			data[51761] <= 8'h10 ;
			data[51762] <= 8'h10 ;
			data[51763] <= 8'h10 ;
			data[51764] <= 8'h10 ;
			data[51765] <= 8'h10 ;
			data[51766] <= 8'h10 ;
			data[51767] <= 8'h10 ;
			data[51768] <= 8'h10 ;
			data[51769] <= 8'h10 ;
			data[51770] <= 8'h10 ;
			data[51771] <= 8'h10 ;
			data[51772] <= 8'h10 ;
			data[51773] <= 8'h10 ;
			data[51774] <= 8'h10 ;
			data[51775] <= 8'h10 ;
			data[51776] <= 8'h10 ;
			data[51777] <= 8'h10 ;
			data[51778] <= 8'h10 ;
			data[51779] <= 8'h10 ;
			data[51780] <= 8'h10 ;
			data[51781] <= 8'h10 ;
			data[51782] <= 8'h10 ;
			data[51783] <= 8'h10 ;
			data[51784] <= 8'h10 ;
			data[51785] <= 8'h10 ;
			data[51786] <= 8'h10 ;
			data[51787] <= 8'h10 ;
			data[51788] <= 8'h10 ;
			data[51789] <= 8'h10 ;
			data[51790] <= 8'h10 ;
			data[51791] <= 8'h10 ;
			data[51792] <= 8'h10 ;
			data[51793] <= 8'h10 ;
			data[51794] <= 8'h10 ;
			data[51795] <= 8'h10 ;
			data[51796] <= 8'h10 ;
			data[51797] <= 8'h10 ;
			data[51798] <= 8'h10 ;
			data[51799] <= 8'h10 ;
			data[51800] <= 8'h10 ;
			data[51801] <= 8'h10 ;
			data[51802] <= 8'h10 ;
			data[51803] <= 8'h10 ;
			data[51804] <= 8'h10 ;
			data[51805] <= 8'h10 ;
			data[51806] <= 8'h10 ;
			data[51807] <= 8'h10 ;
			data[51808] <= 8'h10 ;
			data[51809] <= 8'h10 ;
			data[51810] <= 8'h10 ;
			data[51811] <= 8'h10 ;
			data[51812] <= 8'h10 ;
			data[51813] <= 8'h10 ;
			data[51814] <= 8'h10 ;
			data[51815] <= 8'h10 ;
			data[51816] <= 8'h10 ;
			data[51817] <= 8'h10 ;
			data[51818] <= 8'h10 ;
			data[51819] <= 8'h10 ;
			data[51820] <= 8'h10 ;
			data[51821] <= 8'h10 ;
			data[51822] <= 8'h10 ;
			data[51823] <= 8'h10 ;
			data[51824] <= 8'h10 ;
			data[51825] <= 8'h10 ;
			data[51826] <= 8'h10 ;
			data[51827] <= 8'h10 ;
			data[51828] <= 8'h10 ;
			data[51829] <= 8'h10 ;
			data[51830] <= 8'h10 ;
			data[51831] <= 8'h10 ;
			data[51832] <= 8'h10 ;
			data[51833] <= 8'h10 ;
			data[51834] <= 8'h10 ;
			data[51835] <= 8'h10 ;
			data[51836] <= 8'h10 ;
			data[51837] <= 8'h10 ;
			data[51838] <= 8'h10 ;
			data[51839] <= 8'h10 ;
			data[51840] <= 8'h10 ;
			data[51841] <= 8'h10 ;
			data[51842] <= 8'h10 ;
			data[51843] <= 8'h10 ;
			data[51844] <= 8'h10 ;
			data[51845] <= 8'h10 ;
			data[51846] <= 8'h10 ;
			data[51847] <= 8'h10 ;
			data[51848] <= 8'h10 ;
			data[51849] <= 8'h10 ;
			data[51850] <= 8'h10 ;
			data[51851] <= 8'h10 ;
			data[51852] <= 8'h10 ;
			data[51853] <= 8'h10 ;
			data[51854] <= 8'h10 ;
			data[51855] <= 8'h10 ;
			data[51856] <= 8'h10 ;
			data[51857] <= 8'h10 ;
			data[51858] <= 8'h10 ;
			data[51859] <= 8'h10 ;
			data[51860] <= 8'h10 ;
			data[51861] <= 8'h10 ;
			data[51862] <= 8'h10 ;
			data[51863] <= 8'h10 ;
			data[51864] <= 8'h10 ;
			data[51865] <= 8'h10 ;
			data[51866] <= 8'h10 ;
			data[51867] <= 8'h10 ;
			data[51868] <= 8'h10 ;
			data[51869] <= 8'h10 ;
			data[51870] <= 8'h10 ;
			data[51871] <= 8'h10 ;
			data[51872] <= 8'h10 ;
			data[51873] <= 8'h10 ;
			data[51874] <= 8'h10 ;
			data[51875] <= 8'h10 ;
			data[51876] <= 8'h10 ;
			data[51877] <= 8'h10 ;
			data[51878] <= 8'h10 ;
			data[51879] <= 8'h10 ;
			data[51880] <= 8'h10 ;
			data[51881] <= 8'h10 ;
			data[51882] <= 8'h10 ;
			data[51883] <= 8'h10 ;
			data[51884] <= 8'h10 ;
			data[51885] <= 8'h10 ;
			data[51886] <= 8'h10 ;
			data[51887] <= 8'h10 ;
			data[51888] <= 8'h10 ;
			data[51889] <= 8'h10 ;
			data[51890] <= 8'h10 ;
			data[51891] <= 8'h10 ;
			data[51892] <= 8'h10 ;
			data[51893] <= 8'h10 ;
			data[51894] <= 8'h10 ;
			data[51895] <= 8'h10 ;
			data[51896] <= 8'h10 ;
			data[51897] <= 8'h10 ;
			data[51898] <= 8'h10 ;
			data[51899] <= 8'h10 ;
			data[51900] <= 8'h10 ;
			data[51901] <= 8'h10 ;
			data[51902] <= 8'h10 ;
			data[51903] <= 8'h10 ;
			data[51904] <= 8'h10 ;
			data[51905] <= 8'h10 ;
			data[51906] <= 8'h10 ;
			data[51907] <= 8'h10 ;
			data[51908] <= 8'h10 ;
			data[51909] <= 8'h10 ;
			data[51910] <= 8'h10 ;
			data[51911] <= 8'h10 ;
			data[51912] <= 8'h10 ;
			data[51913] <= 8'h10 ;
			data[51914] <= 8'h10 ;
			data[51915] <= 8'h10 ;
			data[51916] <= 8'h10 ;
			data[51917] <= 8'h10 ;
			data[51918] <= 8'h10 ;
			data[51919] <= 8'h10 ;
			data[51920] <= 8'h10 ;
			data[51921] <= 8'h10 ;
			data[51922] <= 8'h10 ;
			data[51923] <= 8'h10 ;
			data[51924] <= 8'h10 ;
			data[51925] <= 8'h10 ;
			data[51926] <= 8'h10 ;
			data[51927] <= 8'h10 ;
			data[51928] <= 8'h10 ;
			data[51929] <= 8'h10 ;
			data[51930] <= 8'h10 ;
			data[51931] <= 8'h10 ;
			data[51932] <= 8'h10 ;
			data[51933] <= 8'h10 ;
			data[51934] <= 8'h10 ;
			data[51935] <= 8'h10 ;
			data[51936] <= 8'h10 ;
			data[51937] <= 8'h10 ;
			data[51938] <= 8'h10 ;
			data[51939] <= 8'h10 ;
			data[51940] <= 8'h10 ;
			data[51941] <= 8'h10 ;
			data[51942] <= 8'h10 ;
			data[51943] <= 8'h10 ;
			data[51944] <= 8'h10 ;
			data[51945] <= 8'h10 ;
			data[51946] <= 8'h10 ;
			data[51947] <= 8'h10 ;
			data[51948] <= 8'h10 ;
			data[51949] <= 8'h10 ;
			data[51950] <= 8'h10 ;
			data[51951] <= 8'h10 ;
			data[51952] <= 8'h10 ;
			data[51953] <= 8'h10 ;
			data[51954] <= 8'h10 ;
			data[51955] <= 8'h10 ;
			data[51956] <= 8'h10 ;
			data[51957] <= 8'h10 ;
			data[51958] <= 8'h10 ;
			data[51959] <= 8'h10 ;
			data[51960] <= 8'h10 ;
			data[51961] <= 8'h10 ;
			data[51962] <= 8'h10 ;
			data[51963] <= 8'h10 ;
			data[51964] <= 8'h10 ;
			data[51965] <= 8'h10 ;
			data[51966] <= 8'h10 ;
			data[51967] <= 8'h10 ;
			data[51968] <= 8'h10 ;
			data[51969] <= 8'h10 ;
			data[51970] <= 8'h10 ;
			data[51971] <= 8'h10 ;
			data[51972] <= 8'h10 ;
			data[51973] <= 8'h10 ;
			data[51974] <= 8'h10 ;
			data[51975] <= 8'h10 ;
			data[51976] <= 8'h10 ;
			data[51977] <= 8'h10 ;
			data[51978] <= 8'h10 ;
			data[51979] <= 8'h10 ;
			data[51980] <= 8'h10 ;
			data[51981] <= 8'h10 ;
			data[51982] <= 8'h10 ;
			data[51983] <= 8'h10 ;
			data[51984] <= 8'h10 ;
			data[51985] <= 8'h10 ;
			data[51986] <= 8'h10 ;
			data[51987] <= 8'h10 ;
			data[51988] <= 8'h10 ;
			data[51989] <= 8'h10 ;
			data[51990] <= 8'h10 ;
			data[51991] <= 8'h10 ;
			data[51992] <= 8'h10 ;
			data[51993] <= 8'h10 ;
			data[51994] <= 8'h10 ;
			data[51995] <= 8'h10 ;
			data[51996] <= 8'h10 ;
			data[51997] <= 8'h10 ;
			data[51998] <= 8'h10 ;
			data[51999] <= 8'h10 ;
			data[52000] <= 8'h10 ;
			data[52001] <= 8'h10 ;
			data[52002] <= 8'h10 ;
			data[52003] <= 8'h10 ;
			data[52004] <= 8'h10 ;
			data[52005] <= 8'h10 ;
			data[52006] <= 8'h10 ;
			data[52007] <= 8'h10 ;
			data[52008] <= 8'h10 ;
			data[52009] <= 8'h10 ;
			data[52010] <= 8'h10 ;
			data[52011] <= 8'h10 ;
			data[52012] <= 8'h10 ;
			data[52013] <= 8'h10 ;
			data[52014] <= 8'h10 ;
			data[52015] <= 8'h10 ;
			data[52016] <= 8'h10 ;
			data[52017] <= 8'h10 ;
			data[52018] <= 8'h10 ;
			data[52019] <= 8'h10 ;
			data[52020] <= 8'h10 ;
			data[52021] <= 8'h10 ;
			data[52022] <= 8'h10 ;
			data[52023] <= 8'h10 ;
			data[52024] <= 8'h10 ;
			data[52025] <= 8'h10 ;
			data[52026] <= 8'h10 ;
			data[52027] <= 8'h10 ;
			data[52028] <= 8'h10 ;
			data[52029] <= 8'h10 ;
			data[52030] <= 8'h10 ;
			data[52031] <= 8'h10 ;
			data[52032] <= 8'h10 ;
			data[52033] <= 8'h10 ;
			data[52034] <= 8'h10 ;
			data[52035] <= 8'h10 ;
			data[52036] <= 8'h10 ;
			data[52037] <= 8'h10 ;
			data[52038] <= 8'h10 ;
			data[52039] <= 8'h10 ;
			data[52040] <= 8'h10 ;
			data[52041] <= 8'h10 ;
			data[52042] <= 8'h10 ;
			data[52043] <= 8'h10 ;
			data[52044] <= 8'h10 ;
			data[52045] <= 8'h10 ;
			data[52046] <= 8'h10 ;
			data[52047] <= 8'h10 ;
			data[52048] <= 8'h10 ;
			data[52049] <= 8'h10 ;
			data[52050] <= 8'h10 ;
			data[52051] <= 8'h10 ;
			data[52052] <= 8'h10 ;
			data[52053] <= 8'h10 ;
			data[52054] <= 8'h10 ;
			data[52055] <= 8'h10 ;
			data[52056] <= 8'h10 ;
			data[52057] <= 8'h10 ;
			data[52058] <= 8'h10 ;
			data[52059] <= 8'h10 ;
			data[52060] <= 8'h10 ;
			data[52061] <= 8'h10 ;
			data[52062] <= 8'h10 ;
			data[52063] <= 8'h10 ;
			data[52064] <= 8'h10 ;
			data[52065] <= 8'h10 ;
			data[52066] <= 8'h10 ;
			data[52067] <= 8'h10 ;
			data[52068] <= 8'h10 ;
			data[52069] <= 8'h10 ;
			data[52070] <= 8'h10 ;
			data[52071] <= 8'h10 ;
			data[52072] <= 8'h10 ;
			data[52073] <= 8'h10 ;
			data[52074] <= 8'h10 ;
			data[52075] <= 8'h10 ;
			data[52076] <= 8'h10 ;
			data[52077] <= 8'h10 ;
			data[52078] <= 8'h10 ;
			data[52079] <= 8'h10 ;
			data[52080] <= 8'h10 ;
			data[52081] <= 8'h10 ;
			data[52082] <= 8'h10 ;
			data[52083] <= 8'h10 ;
			data[52084] <= 8'h10 ;
			data[52085] <= 8'h10 ;
			data[52086] <= 8'h10 ;
			data[52087] <= 8'h10 ;
			data[52088] <= 8'h10 ;
			data[52089] <= 8'h10 ;
			data[52090] <= 8'h10 ;
			data[52091] <= 8'h10 ;
			data[52092] <= 8'h10 ;
			data[52093] <= 8'h10 ;
			data[52094] <= 8'h10 ;
			data[52095] <= 8'h10 ;
			data[52096] <= 8'h10 ;
			data[52097] <= 8'h10 ;
			data[52098] <= 8'h10 ;
			data[52099] <= 8'h10 ;
			data[52100] <= 8'h10 ;
			data[52101] <= 8'h10 ;
			data[52102] <= 8'h10 ;
			data[52103] <= 8'h10 ;
			data[52104] <= 8'h10 ;
			data[52105] <= 8'h10 ;
			data[52106] <= 8'h10 ;
			data[52107] <= 8'h10 ;
			data[52108] <= 8'h10 ;
			data[52109] <= 8'h10 ;
			data[52110] <= 8'h10 ;
			data[52111] <= 8'h10 ;
			data[52112] <= 8'h10 ;
			data[52113] <= 8'h10 ;
			data[52114] <= 8'h10 ;
			data[52115] <= 8'h10 ;
			data[52116] <= 8'h10 ;
			data[52117] <= 8'h10 ;
			data[52118] <= 8'h10 ;
			data[52119] <= 8'h10 ;
			data[52120] <= 8'h10 ;
			data[52121] <= 8'h10 ;
			data[52122] <= 8'h10 ;
			data[52123] <= 8'h10 ;
			data[52124] <= 8'h10 ;
			data[52125] <= 8'h10 ;
			data[52126] <= 8'h10 ;
			data[52127] <= 8'h10 ;
			data[52128] <= 8'h10 ;
			data[52129] <= 8'h10 ;
			data[52130] <= 8'h10 ;
			data[52131] <= 8'h10 ;
			data[52132] <= 8'h10 ;
			data[52133] <= 8'h10 ;
			data[52134] <= 8'h10 ;
			data[52135] <= 8'h10 ;
			data[52136] <= 8'h10 ;
			data[52137] <= 8'h10 ;
			data[52138] <= 8'h10 ;
			data[52139] <= 8'h10 ;
			data[52140] <= 8'h10 ;
			data[52141] <= 8'h10 ;
			data[52142] <= 8'h10 ;
			data[52143] <= 8'h10 ;
			data[52144] <= 8'h10 ;
			data[52145] <= 8'h10 ;
			data[52146] <= 8'h10 ;
			data[52147] <= 8'h10 ;
			data[52148] <= 8'h10 ;
			data[52149] <= 8'h10 ;
			data[52150] <= 8'h10 ;
			data[52151] <= 8'h10 ;
			data[52152] <= 8'h10 ;
			data[52153] <= 8'h10 ;
			data[52154] <= 8'h10 ;
			data[52155] <= 8'h10 ;
			data[52156] <= 8'h10 ;
			data[52157] <= 8'h10 ;
			data[52158] <= 8'h10 ;
			data[52159] <= 8'h10 ;
			data[52160] <= 8'h10 ;
			data[52161] <= 8'h10 ;
			data[52162] <= 8'h10 ;
			data[52163] <= 8'h10 ;
			data[52164] <= 8'h10 ;
			data[52165] <= 8'h10 ;
			data[52166] <= 8'h10 ;
			data[52167] <= 8'h10 ;
			data[52168] <= 8'h10 ;
			data[52169] <= 8'h10 ;
			data[52170] <= 8'h10 ;
			data[52171] <= 8'h10 ;
			data[52172] <= 8'h10 ;
			data[52173] <= 8'h10 ;
			data[52174] <= 8'h10 ;
			data[52175] <= 8'h10 ;
			data[52176] <= 8'h10 ;
			data[52177] <= 8'h10 ;
			data[52178] <= 8'h10 ;
			data[52179] <= 8'h10 ;
			data[52180] <= 8'h10 ;
			data[52181] <= 8'h10 ;
			data[52182] <= 8'h10 ;
			data[52183] <= 8'h10 ;
			data[52184] <= 8'h10 ;
			data[52185] <= 8'h10 ;
			data[52186] <= 8'h10 ;
			data[52187] <= 8'h10 ;
			data[52188] <= 8'h10 ;
			data[52189] <= 8'h10 ;
			data[52190] <= 8'h10 ;
			data[52191] <= 8'h10 ;
			data[52192] <= 8'h10 ;
			data[52193] <= 8'h10 ;
			data[52194] <= 8'h10 ;
			data[52195] <= 8'h10 ;
			data[52196] <= 8'h10 ;
			data[52197] <= 8'h10 ;
			data[52198] <= 8'h10 ;
			data[52199] <= 8'h10 ;
			data[52200] <= 8'h10 ;
			data[52201] <= 8'h10 ;
			data[52202] <= 8'h10 ;
			data[52203] <= 8'h10 ;
			data[52204] <= 8'h10 ;
			data[52205] <= 8'h10 ;
			data[52206] <= 8'h10 ;
			data[52207] <= 8'h10 ;
			data[52208] <= 8'h10 ;
			data[52209] <= 8'h10 ;
			data[52210] <= 8'h10 ;
			data[52211] <= 8'h10 ;
			data[52212] <= 8'h10 ;
			data[52213] <= 8'h10 ;
			data[52214] <= 8'h10 ;
			data[52215] <= 8'h10 ;
			data[52216] <= 8'h10 ;
			data[52217] <= 8'h10 ;
			data[52218] <= 8'h10 ;
			data[52219] <= 8'h10 ;
			data[52220] <= 8'h10 ;
			data[52221] <= 8'h10 ;
			data[52222] <= 8'h10 ;
			data[52223] <= 8'h10 ;
			data[52224] <= 8'h10 ;
			data[52225] <= 8'h10 ;
			data[52226] <= 8'h10 ;
			data[52227] <= 8'h10 ;
			data[52228] <= 8'h10 ;
			data[52229] <= 8'h10 ;
			data[52230] <= 8'h10 ;
			data[52231] <= 8'h10 ;
			data[52232] <= 8'h10 ;
			data[52233] <= 8'h10 ;
			data[52234] <= 8'h10 ;
			data[52235] <= 8'h10 ;
			data[52236] <= 8'h10 ;
			data[52237] <= 8'h10 ;
			data[52238] <= 8'h10 ;
			data[52239] <= 8'h10 ;
			data[52240] <= 8'h10 ;
			data[52241] <= 8'h10 ;
			data[52242] <= 8'h10 ;
			data[52243] <= 8'h10 ;
			data[52244] <= 8'h10 ;
			data[52245] <= 8'h10 ;
			data[52246] <= 8'h10 ;
			data[52247] <= 8'h10 ;
			data[52248] <= 8'h10 ;
			data[52249] <= 8'h10 ;
			data[52250] <= 8'h10 ;
			data[52251] <= 8'h10 ;
			data[52252] <= 8'h10 ;
			data[52253] <= 8'h10 ;
			data[52254] <= 8'h10 ;
			data[52255] <= 8'h10 ;
			data[52256] <= 8'h10 ;
			data[52257] <= 8'h10 ;
			data[52258] <= 8'h10 ;
			data[52259] <= 8'h10 ;
			data[52260] <= 8'h10 ;
			data[52261] <= 8'h10 ;
			data[52262] <= 8'h10 ;
			data[52263] <= 8'h10 ;
			data[52264] <= 8'h10 ;
			data[52265] <= 8'h10 ;
			data[52266] <= 8'h10 ;
			data[52267] <= 8'h10 ;
			data[52268] <= 8'h10 ;
			data[52269] <= 8'h10 ;
			data[52270] <= 8'h10 ;
			data[52271] <= 8'h10 ;
			data[52272] <= 8'h10 ;
			data[52273] <= 8'h10 ;
			data[52274] <= 8'h10 ;
			data[52275] <= 8'h10 ;
			data[52276] <= 8'h10 ;
			data[52277] <= 8'h10 ;
			data[52278] <= 8'h10 ;
			data[52279] <= 8'h10 ;
			data[52280] <= 8'h10 ;
			data[52281] <= 8'h10 ;
			data[52282] <= 8'h10 ;
			data[52283] <= 8'h10 ;
			data[52284] <= 8'h10 ;
			data[52285] <= 8'h10 ;
			data[52286] <= 8'h10 ;
			data[52287] <= 8'h10 ;
			data[52288] <= 8'h10 ;
			data[52289] <= 8'h10 ;
			data[52290] <= 8'h10 ;
			data[52291] <= 8'h10 ;
			data[52292] <= 8'h10 ;
			data[52293] <= 8'h10 ;
			data[52294] <= 8'h10 ;
			data[52295] <= 8'h10 ;
			data[52296] <= 8'h10 ;
			data[52297] <= 8'h10 ;
			data[52298] <= 8'h10 ;
			data[52299] <= 8'h10 ;
			data[52300] <= 8'h10 ;
			data[52301] <= 8'h10 ;
			data[52302] <= 8'h10 ;
			data[52303] <= 8'h10 ;
			data[52304] <= 8'h10 ;
			data[52305] <= 8'h10 ;
			data[52306] <= 8'h10 ;
			data[52307] <= 8'h10 ;
			data[52308] <= 8'h10 ;
			data[52309] <= 8'h10 ;
			data[52310] <= 8'h10 ;
			data[52311] <= 8'h10 ;
			data[52312] <= 8'h10 ;
			data[52313] <= 8'h10 ;
			data[52314] <= 8'h10 ;
			data[52315] <= 8'h10 ;
			data[52316] <= 8'h10 ;
			data[52317] <= 8'h10 ;
			data[52318] <= 8'h10 ;
			data[52319] <= 8'h10 ;
			data[52320] <= 8'h10 ;
			data[52321] <= 8'h10 ;
			data[52322] <= 8'h10 ;
			data[52323] <= 8'h10 ;
			data[52324] <= 8'h10 ;
			data[52325] <= 8'h10 ;
			data[52326] <= 8'h10 ;
			data[52327] <= 8'h10 ;
			data[52328] <= 8'h10 ;
			data[52329] <= 8'h10 ;
			data[52330] <= 8'h10 ;
			data[52331] <= 8'h10 ;
			data[52332] <= 8'h10 ;
			data[52333] <= 8'h10 ;
			data[52334] <= 8'h10 ;
			data[52335] <= 8'h10 ;
			data[52336] <= 8'h10 ;
			data[52337] <= 8'h10 ;
			data[52338] <= 8'h10 ;
			data[52339] <= 8'h10 ;
			data[52340] <= 8'h10 ;
			data[52341] <= 8'h10 ;
			data[52342] <= 8'h10 ;
			data[52343] <= 8'h10 ;
			data[52344] <= 8'h10 ;
			data[52345] <= 8'h10 ;
			data[52346] <= 8'h10 ;
			data[52347] <= 8'h10 ;
			data[52348] <= 8'h10 ;
			data[52349] <= 8'h10 ;
			data[52350] <= 8'h10 ;
			data[52351] <= 8'h10 ;
			data[52352] <= 8'h10 ;
			data[52353] <= 8'h10 ;
			data[52354] <= 8'h10 ;
			data[52355] <= 8'h10 ;
			data[52356] <= 8'h10 ;
			data[52357] <= 8'h10 ;
			data[52358] <= 8'h10 ;
			data[52359] <= 8'h10 ;
			data[52360] <= 8'h10 ;
			data[52361] <= 8'h10 ;
			data[52362] <= 8'h10 ;
			data[52363] <= 8'h10 ;
			data[52364] <= 8'h10 ;
			data[52365] <= 8'h10 ;
			data[52366] <= 8'h10 ;
			data[52367] <= 8'h10 ;
			data[52368] <= 8'h10 ;
			data[52369] <= 8'h10 ;
			data[52370] <= 8'h10 ;
			data[52371] <= 8'h10 ;
			data[52372] <= 8'h10 ;
			data[52373] <= 8'h10 ;
			data[52374] <= 8'h10 ;
			data[52375] <= 8'h10 ;
			data[52376] <= 8'h10 ;
			data[52377] <= 8'h10 ;
			data[52378] <= 8'h10 ;
			data[52379] <= 8'h10 ;
			data[52380] <= 8'h10 ;
			data[52381] <= 8'h10 ;
			data[52382] <= 8'h10 ;
			data[52383] <= 8'h10 ;
			data[52384] <= 8'h10 ;
			data[52385] <= 8'h10 ;
			data[52386] <= 8'h10 ;
			data[52387] <= 8'h10 ;
			data[52388] <= 8'h10 ;
			data[52389] <= 8'h10 ;
			data[52390] <= 8'h10 ;
			data[52391] <= 8'h10 ;
			data[52392] <= 8'h10 ;
			data[52393] <= 8'h10 ;
			data[52394] <= 8'h10 ;
			data[52395] <= 8'h10 ;
			data[52396] <= 8'h10 ;
			data[52397] <= 8'h10 ;
			data[52398] <= 8'h10 ;
			data[52399] <= 8'h10 ;
			data[52400] <= 8'h10 ;
			data[52401] <= 8'h10 ;
			data[52402] <= 8'h10 ;
			data[52403] <= 8'h10 ;
			data[52404] <= 8'h10 ;
			data[52405] <= 8'h10 ;
			data[52406] <= 8'h10 ;
			data[52407] <= 8'h10 ;
			data[52408] <= 8'h10 ;
			data[52409] <= 8'h10 ;
			data[52410] <= 8'h10 ;
			data[52411] <= 8'h10 ;
			data[52412] <= 8'h10 ;
			data[52413] <= 8'h10 ;
			data[52414] <= 8'h10 ;
			data[52415] <= 8'h10 ;
			data[52416] <= 8'h10 ;
			data[52417] <= 8'h10 ;
			data[52418] <= 8'h10 ;
			data[52419] <= 8'h10 ;
			data[52420] <= 8'h10 ;
			data[52421] <= 8'h10 ;
			data[52422] <= 8'h10 ;
			data[52423] <= 8'h10 ;
			data[52424] <= 8'h10 ;
			data[52425] <= 8'h10 ;
			data[52426] <= 8'h10 ;
			data[52427] <= 8'h10 ;
			data[52428] <= 8'h10 ;
			data[52429] <= 8'h10 ;
			data[52430] <= 8'h10 ;
			data[52431] <= 8'h10 ;
			data[52432] <= 8'h10 ;
			data[52433] <= 8'h10 ;
			data[52434] <= 8'h10 ;
			data[52435] <= 8'h10 ;
			data[52436] <= 8'h10 ;
			data[52437] <= 8'h10 ;
			data[52438] <= 8'h10 ;
			data[52439] <= 8'h10 ;
			data[52440] <= 8'h10 ;
			data[52441] <= 8'h10 ;
			data[52442] <= 8'h10 ;
			data[52443] <= 8'h10 ;
			data[52444] <= 8'h10 ;
			data[52445] <= 8'h10 ;
			data[52446] <= 8'h10 ;
			data[52447] <= 8'h10 ;
			data[52448] <= 8'h10 ;
			data[52449] <= 8'h10 ;
			data[52450] <= 8'h10 ;
			data[52451] <= 8'h10 ;
			data[52452] <= 8'h10 ;
			data[52453] <= 8'h10 ;
			data[52454] <= 8'h10 ;
			data[52455] <= 8'h10 ;
			data[52456] <= 8'h10 ;
			data[52457] <= 8'h10 ;
			data[52458] <= 8'h10 ;
			data[52459] <= 8'h10 ;
			data[52460] <= 8'h10 ;
			data[52461] <= 8'h10 ;
			data[52462] <= 8'h10 ;
			data[52463] <= 8'h10 ;
			data[52464] <= 8'h10 ;
			data[52465] <= 8'h10 ;
			data[52466] <= 8'h10 ;
			data[52467] <= 8'h10 ;
			data[52468] <= 8'h10 ;
			data[52469] <= 8'h10 ;
			data[52470] <= 8'h10 ;
			data[52471] <= 8'h10 ;
			data[52472] <= 8'h10 ;
			data[52473] <= 8'h10 ;
			data[52474] <= 8'h10 ;
			data[52475] <= 8'h10 ;
			data[52476] <= 8'h10 ;
			data[52477] <= 8'h10 ;
			data[52478] <= 8'h10 ;
			data[52479] <= 8'h10 ;
			data[52480] <= 8'h10 ;
			data[52481] <= 8'h10 ;
			data[52482] <= 8'h10 ;
			data[52483] <= 8'h10 ;
			data[52484] <= 8'h10 ;
			data[52485] <= 8'h10 ;
			data[52486] <= 8'h10 ;
			data[52487] <= 8'h10 ;
			data[52488] <= 8'h10 ;
			data[52489] <= 8'h10 ;
			data[52490] <= 8'h10 ;
			data[52491] <= 8'h10 ;
			data[52492] <= 8'h10 ;
			data[52493] <= 8'h10 ;
			data[52494] <= 8'h10 ;
			data[52495] <= 8'h10 ;
			data[52496] <= 8'h10 ;
			data[52497] <= 8'h10 ;
			data[52498] <= 8'h10 ;
			data[52499] <= 8'h10 ;
			data[52500] <= 8'h10 ;
			data[52501] <= 8'h10 ;
			data[52502] <= 8'h10 ;
			data[52503] <= 8'h10 ;
			data[52504] <= 8'h10 ;
			data[52505] <= 8'h10 ;
			data[52506] <= 8'h10 ;
			data[52507] <= 8'h10 ;
			data[52508] <= 8'h10 ;
			data[52509] <= 8'h10 ;
			data[52510] <= 8'h10 ;
			data[52511] <= 8'h10 ;
			data[52512] <= 8'h10 ;
			data[52513] <= 8'h10 ;
			data[52514] <= 8'h10 ;
			data[52515] <= 8'h10 ;
			data[52516] <= 8'h10 ;
			data[52517] <= 8'h10 ;
			data[52518] <= 8'h10 ;
			data[52519] <= 8'h10 ;
			data[52520] <= 8'h10 ;
			data[52521] <= 8'h10 ;
			data[52522] <= 8'h10 ;
			data[52523] <= 8'h10 ;
			data[52524] <= 8'h10 ;
			data[52525] <= 8'h10 ;
			data[52526] <= 8'h10 ;
			data[52527] <= 8'h10 ;
			data[52528] <= 8'h10 ;
			data[52529] <= 8'h10 ;
			data[52530] <= 8'h10 ;
			data[52531] <= 8'h10 ;
			data[52532] <= 8'h10 ;
			data[52533] <= 8'h10 ;
			data[52534] <= 8'h10 ;
			data[52535] <= 8'h10 ;
			data[52536] <= 8'h10 ;
			data[52537] <= 8'h10 ;
			data[52538] <= 8'h10 ;
			data[52539] <= 8'h10 ;
			data[52540] <= 8'h10 ;
			data[52541] <= 8'h10 ;
			data[52542] <= 8'h10 ;
			data[52543] <= 8'h10 ;
			data[52544] <= 8'h10 ;
			data[52545] <= 8'h10 ;
			data[52546] <= 8'h10 ;
			data[52547] <= 8'h10 ;
			data[52548] <= 8'h10 ;
			data[52549] <= 8'h10 ;
			data[52550] <= 8'h10 ;
			data[52551] <= 8'h10 ;
			data[52552] <= 8'h10 ;
			data[52553] <= 8'h10 ;
			data[52554] <= 8'h10 ;
			data[52555] <= 8'h10 ;
			data[52556] <= 8'h10 ;
			data[52557] <= 8'h10 ;
			data[52558] <= 8'h10 ;
			data[52559] <= 8'h10 ;
			data[52560] <= 8'h10 ;
			data[52561] <= 8'h10 ;
			data[52562] <= 8'h10 ;
			data[52563] <= 8'h10 ;
			data[52564] <= 8'h10 ;
			data[52565] <= 8'h10 ;
			data[52566] <= 8'h10 ;
			data[52567] <= 8'h10 ;
			data[52568] <= 8'h10 ;
			data[52569] <= 8'h10 ;
			data[52570] <= 8'h10 ;
			data[52571] <= 8'h10 ;
			data[52572] <= 8'h10 ;
			data[52573] <= 8'h10 ;
			data[52574] <= 8'h10 ;
			data[52575] <= 8'h10 ;
			data[52576] <= 8'h10 ;
			data[52577] <= 8'h10 ;
			data[52578] <= 8'h10 ;
			data[52579] <= 8'h10 ;
			data[52580] <= 8'h10 ;
			data[52581] <= 8'h10 ;
			data[52582] <= 8'h10 ;
			data[52583] <= 8'h10 ;
			data[52584] <= 8'h10 ;
			data[52585] <= 8'h10 ;
			data[52586] <= 8'h10 ;
			data[52587] <= 8'h10 ;
			data[52588] <= 8'h10 ;
			data[52589] <= 8'h10 ;
			data[52590] <= 8'h10 ;
			data[52591] <= 8'h10 ;
			data[52592] <= 8'h10 ;
			data[52593] <= 8'h10 ;
			data[52594] <= 8'h10 ;
			data[52595] <= 8'h10 ;
			data[52596] <= 8'h10 ;
			data[52597] <= 8'h10 ;
			data[52598] <= 8'h10 ;
			data[52599] <= 8'h10 ;
			data[52600] <= 8'h10 ;
			data[52601] <= 8'h10 ;
			data[52602] <= 8'h10 ;
			data[52603] <= 8'h10 ;
			data[52604] <= 8'h10 ;
			data[52605] <= 8'h10 ;
			data[52606] <= 8'h10 ;
			data[52607] <= 8'h10 ;
			data[52608] <= 8'h10 ;
			data[52609] <= 8'h10 ;
			data[52610] <= 8'h10 ;
			data[52611] <= 8'h10 ;
			data[52612] <= 8'h10 ;
			data[52613] <= 8'h10 ;
			data[52614] <= 8'h10 ;
			data[52615] <= 8'h10 ;
			data[52616] <= 8'h10 ;
			data[52617] <= 8'h10 ;
			data[52618] <= 8'h10 ;
			data[52619] <= 8'h10 ;
			data[52620] <= 8'h10 ;
			data[52621] <= 8'h10 ;
			data[52622] <= 8'h10 ;
			data[52623] <= 8'h10 ;
			data[52624] <= 8'h10 ;
			data[52625] <= 8'h10 ;
			data[52626] <= 8'h10 ;
			data[52627] <= 8'h10 ;
			data[52628] <= 8'h10 ;
			data[52629] <= 8'h10 ;
			data[52630] <= 8'h10 ;
			data[52631] <= 8'h10 ;
			data[52632] <= 8'h10 ;
			data[52633] <= 8'h10 ;
			data[52634] <= 8'h10 ;
			data[52635] <= 8'h10 ;
			data[52636] <= 8'h10 ;
			data[52637] <= 8'h10 ;
			data[52638] <= 8'h10 ;
			data[52639] <= 8'h10 ;
			data[52640] <= 8'h10 ;
			data[52641] <= 8'h10 ;
			data[52642] <= 8'h10 ;
			data[52643] <= 8'h10 ;
			data[52644] <= 8'h10 ;
			data[52645] <= 8'h10 ;
			data[52646] <= 8'h10 ;
			data[52647] <= 8'h10 ;
			data[52648] <= 8'h10 ;
			data[52649] <= 8'h10 ;
			data[52650] <= 8'h10 ;
			data[52651] <= 8'h10 ;
			data[52652] <= 8'h10 ;
			data[52653] <= 8'h10 ;
			data[52654] <= 8'h10 ;
			data[52655] <= 8'h10 ;
			data[52656] <= 8'h10 ;
			data[52657] <= 8'h10 ;
			data[52658] <= 8'h10 ;
			data[52659] <= 8'h10 ;
			data[52660] <= 8'h10 ;
			data[52661] <= 8'h10 ;
			data[52662] <= 8'h10 ;
			data[52663] <= 8'h10 ;
			data[52664] <= 8'h10 ;
			data[52665] <= 8'h10 ;
			data[52666] <= 8'h10 ;
			data[52667] <= 8'h10 ;
			data[52668] <= 8'h10 ;
			data[52669] <= 8'h10 ;
			data[52670] <= 8'h10 ;
			data[52671] <= 8'h10 ;
			data[52672] <= 8'h10 ;
			data[52673] <= 8'h10 ;
			data[52674] <= 8'h10 ;
			data[52675] <= 8'h10 ;
			data[52676] <= 8'h10 ;
			data[52677] <= 8'h10 ;
			data[52678] <= 8'h10 ;
			data[52679] <= 8'h10 ;
			data[52680] <= 8'h10 ;
			data[52681] <= 8'h10 ;
			data[52682] <= 8'h10 ;
			data[52683] <= 8'h10 ;
			data[52684] <= 8'h10 ;
			data[52685] <= 8'h10 ;
			data[52686] <= 8'h10 ;
			data[52687] <= 8'h10 ;
			data[52688] <= 8'h10 ;
			data[52689] <= 8'h10 ;
			data[52690] <= 8'h10 ;
			data[52691] <= 8'h10 ;
			data[52692] <= 8'h10 ;
			data[52693] <= 8'h10 ;
			data[52694] <= 8'h10 ;
			data[52695] <= 8'h10 ;
			data[52696] <= 8'h10 ;
			data[52697] <= 8'h10 ;
			data[52698] <= 8'h10 ;
			data[52699] <= 8'h10 ;
			data[52700] <= 8'h10 ;
			data[52701] <= 8'h10 ;
			data[52702] <= 8'h10 ;
			data[52703] <= 8'h10 ;
			data[52704] <= 8'h10 ;
			data[52705] <= 8'h10 ;
			data[52706] <= 8'h10 ;
			data[52707] <= 8'h10 ;
			data[52708] <= 8'h10 ;
			data[52709] <= 8'h10 ;
			data[52710] <= 8'h10 ;
			data[52711] <= 8'h10 ;
			data[52712] <= 8'h10 ;
			data[52713] <= 8'h10 ;
			data[52714] <= 8'h10 ;
			data[52715] <= 8'h10 ;
			data[52716] <= 8'h10 ;
			data[52717] <= 8'h10 ;
			data[52718] <= 8'h10 ;
			data[52719] <= 8'h10 ;
			data[52720] <= 8'h10 ;
			data[52721] <= 8'h10 ;
			data[52722] <= 8'h10 ;
			data[52723] <= 8'h10 ;
			data[52724] <= 8'h10 ;
			data[52725] <= 8'h10 ;
			data[52726] <= 8'h10 ;
			data[52727] <= 8'h10 ;
			data[52728] <= 8'h10 ;
			data[52729] <= 8'h10 ;
			data[52730] <= 8'h10 ;
			data[52731] <= 8'h10 ;
			data[52732] <= 8'h10 ;
			data[52733] <= 8'h10 ;
			data[52734] <= 8'h10 ;
			data[52735] <= 8'h10 ;
			data[52736] <= 8'h10 ;
			data[52737] <= 8'h10 ;
			data[52738] <= 8'h10 ;
			data[52739] <= 8'h10 ;
			data[52740] <= 8'h10 ;
			data[52741] <= 8'h10 ;
			data[52742] <= 8'h10 ;
			data[52743] <= 8'h10 ;
			data[52744] <= 8'h10 ;
			data[52745] <= 8'h10 ;
			data[52746] <= 8'h10 ;
			data[52747] <= 8'h10 ;
			data[52748] <= 8'h10 ;
			data[52749] <= 8'h10 ;
			data[52750] <= 8'h10 ;
			data[52751] <= 8'h10 ;
			data[52752] <= 8'h10 ;
			data[52753] <= 8'h10 ;
			data[52754] <= 8'h10 ;
			data[52755] <= 8'h10 ;
			data[52756] <= 8'h10 ;
			data[52757] <= 8'h10 ;
			data[52758] <= 8'h10 ;
			data[52759] <= 8'h10 ;
			data[52760] <= 8'h10 ;
			data[52761] <= 8'h10 ;
			data[52762] <= 8'h10 ;
			data[52763] <= 8'h10 ;
			data[52764] <= 8'h10 ;
			data[52765] <= 8'h10 ;
			data[52766] <= 8'h10 ;
			data[52767] <= 8'h10 ;
			data[52768] <= 8'h10 ;
			data[52769] <= 8'h10 ;
			data[52770] <= 8'h10 ;
			data[52771] <= 8'h10 ;
			data[52772] <= 8'h10 ;
			data[52773] <= 8'h10 ;
			data[52774] <= 8'h10 ;
			data[52775] <= 8'h10 ;
			data[52776] <= 8'h10 ;
			data[52777] <= 8'h10 ;
			data[52778] <= 8'h10 ;
			data[52779] <= 8'h10 ;
			data[52780] <= 8'h10 ;
			data[52781] <= 8'h10 ;
			data[52782] <= 8'h10 ;
			data[52783] <= 8'h10 ;
			data[52784] <= 8'h10 ;
			data[52785] <= 8'h10 ;
			data[52786] <= 8'h10 ;
			data[52787] <= 8'h10 ;
			data[52788] <= 8'h10 ;
			data[52789] <= 8'h10 ;
			data[52790] <= 8'h10 ;
			data[52791] <= 8'h10 ;
			data[52792] <= 8'h10 ;
			data[52793] <= 8'h10 ;
			data[52794] <= 8'h10 ;
			data[52795] <= 8'h10 ;
			data[52796] <= 8'h10 ;
			data[52797] <= 8'h10 ;
			data[52798] <= 8'h10 ;
			data[52799] <= 8'h10 ;
			data[52800] <= 8'h10 ;
			data[52801] <= 8'h10 ;
			data[52802] <= 8'h10 ;
			data[52803] <= 8'h10 ;
			data[52804] <= 8'h10 ;
			data[52805] <= 8'h10 ;
			data[52806] <= 8'h10 ;
			data[52807] <= 8'h10 ;
			data[52808] <= 8'h10 ;
			data[52809] <= 8'h10 ;
			data[52810] <= 8'h10 ;
			data[52811] <= 8'h10 ;
			data[52812] <= 8'h10 ;
			data[52813] <= 8'h10 ;
			data[52814] <= 8'h10 ;
			data[52815] <= 8'h10 ;
			data[52816] <= 8'h10 ;
			data[52817] <= 8'h10 ;
			data[52818] <= 8'h10 ;
			data[52819] <= 8'h10 ;
			data[52820] <= 8'h10 ;
			data[52821] <= 8'h10 ;
			data[52822] <= 8'h10 ;
			data[52823] <= 8'h10 ;
			data[52824] <= 8'h10 ;
			data[52825] <= 8'h10 ;
			data[52826] <= 8'h10 ;
			data[52827] <= 8'h10 ;
			data[52828] <= 8'h10 ;
			data[52829] <= 8'h10 ;
			data[52830] <= 8'h10 ;
			data[52831] <= 8'h10 ;
			data[52832] <= 8'h10 ;
			data[52833] <= 8'h10 ;
			data[52834] <= 8'h10 ;
			data[52835] <= 8'h10 ;
			data[52836] <= 8'h10 ;
			data[52837] <= 8'h10 ;
			data[52838] <= 8'h10 ;
			data[52839] <= 8'h10 ;
			data[52840] <= 8'h10 ;
			data[52841] <= 8'h10 ;
			data[52842] <= 8'h10 ;
			data[52843] <= 8'h10 ;
			data[52844] <= 8'h10 ;
			data[52845] <= 8'h10 ;
			data[52846] <= 8'h10 ;
			data[52847] <= 8'h10 ;
			data[52848] <= 8'h10 ;
			data[52849] <= 8'h10 ;
			data[52850] <= 8'h10 ;
			data[52851] <= 8'h10 ;
			data[52852] <= 8'h10 ;
			data[52853] <= 8'h10 ;
			data[52854] <= 8'h10 ;
			data[52855] <= 8'h10 ;
			data[52856] <= 8'h10 ;
			data[52857] <= 8'h10 ;
			data[52858] <= 8'h10 ;
			data[52859] <= 8'h10 ;
			data[52860] <= 8'h10 ;
			data[52861] <= 8'h10 ;
			data[52862] <= 8'h10 ;
			data[52863] <= 8'h10 ;
			data[52864] <= 8'h10 ;
			data[52865] <= 8'h10 ;
			data[52866] <= 8'h10 ;
			data[52867] <= 8'h10 ;
			data[52868] <= 8'h10 ;
			data[52869] <= 8'h10 ;
			data[52870] <= 8'h10 ;
			data[52871] <= 8'h10 ;
			data[52872] <= 8'h10 ;
			data[52873] <= 8'h10 ;
			data[52874] <= 8'h10 ;
			data[52875] <= 8'h10 ;
			data[52876] <= 8'h10 ;
			data[52877] <= 8'h10 ;
			data[52878] <= 8'h10 ;
			data[52879] <= 8'h10 ;
			data[52880] <= 8'h10 ;
			data[52881] <= 8'h10 ;
			data[52882] <= 8'h10 ;
			data[52883] <= 8'h10 ;
			data[52884] <= 8'h10 ;
			data[52885] <= 8'h10 ;
			data[52886] <= 8'h10 ;
			data[52887] <= 8'h10 ;
			data[52888] <= 8'h10 ;
			data[52889] <= 8'h10 ;
			data[52890] <= 8'h10 ;
			data[52891] <= 8'h10 ;
			data[52892] <= 8'h10 ;
			data[52893] <= 8'h10 ;
			data[52894] <= 8'h10 ;
			data[52895] <= 8'h10 ;
			data[52896] <= 8'h10 ;
			data[52897] <= 8'h10 ;
			data[52898] <= 8'h10 ;
			data[52899] <= 8'h10 ;
			data[52900] <= 8'h10 ;
			data[52901] <= 8'h10 ;
			data[52902] <= 8'h10 ;
			data[52903] <= 8'h10 ;
			data[52904] <= 8'h10 ;
			data[52905] <= 8'h10 ;
			data[52906] <= 8'h10 ;
			data[52907] <= 8'h10 ;
			data[52908] <= 8'h10 ;
			data[52909] <= 8'h10 ;
			data[52910] <= 8'h10 ;
			data[52911] <= 8'h10 ;
			data[52912] <= 8'h10 ;
			data[52913] <= 8'h10 ;
			data[52914] <= 8'h10 ;
			data[52915] <= 8'h10 ;
			data[52916] <= 8'h10 ;
			data[52917] <= 8'h10 ;
			data[52918] <= 8'h10 ;
			data[52919] <= 8'h10 ;
			data[52920] <= 8'h10 ;
			data[52921] <= 8'h10 ;
			data[52922] <= 8'h10 ;
			data[52923] <= 8'h10 ;
			data[52924] <= 8'h10 ;
			data[52925] <= 8'h10 ;
			data[52926] <= 8'h10 ;
			data[52927] <= 8'h10 ;
			data[52928] <= 8'h10 ;
			data[52929] <= 8'h10 ;
			data[52930] <= 8'h10 ;
			data[52931] <= 8'h10 ;
			data[52932] <= 8'h10 ;
			data[52933] <= 8'h10 ;
			data[52934] <= 8'h10 ;
			data[52935] <= 8'h10 ;
			data[52936] <= 8'h10 ;
			data[52937] <= 8'h10 ;
			data[52938] <= 8'h10 ;
			data[52939] <= 8'h10 ;
			data[52940] <= 8'h10 ;
			data[52941] <= 8'h10 ;
			data[52942] <= 8'h10 ;
			data[52943] <= 8'h10 ;
			data[52944] <= 8'h10 ;
			data[52945] <= 8'h10 ;
			data[52946] <= 8'h10 ;
			data[52947] <= 8'h10 ;
			data[52948] <= 8'h10 ;
			data[52949] <= 8'h10 ;
			data[52950] <= 8'h10 ;
			data[52951] <= 8'h10 ;
			data[52952] <= 8'h10 ;
			data[52953] <= 8'h10 ;
			data[52954] <= 8'h10 ;
			data[52955] <= 8'h10 ;
			data[52956] <= 8'h10 ;
			data[52957] <= 8'h10 ;
			data[52958] <= 8'h10 ;
			data[52959] <= 8'h10 ;
			data[52960] <= 8'h10 ;
			data[52961] <= 8'h10 ;
			data[52962] <= 8'h10 ;
			data[52963] <= 8'h10 ;
			data[52964] <= 8'h10 ;
			data[52965] <= 8'h10 ;
			data[52966] <= 8'h10 ;
			data[52967] <= 8'h10 ;
			data[52968] <= 8'h10 ;
			data[52969] <= 8'h10 ;
			data[52970] <= 8'h10 ;
			data[52971] <= 8'h10 ;
			data[52972] <= 8'h10 ;
			data[52973] <= 8'h10 ;
			data[52974] <= 8'h10 ;
			data[52975] <= 8'h10 ;
			data[52976] <= 8'h10 ;
			data[52977] <= 8'h10 ;
			data[52978] <= 8'h10 ;
			data[52979] <= 8'h10 ;
			data[52980] <= 8'h10 ;
			data[52981] <= 8'h10 ;
			data[52982] <= 8'h10 ;
			data[52983] <= 8'h10 ;
			data[52984] <= 8'h10 ;
			data[52985] <= 8'h10 ;
			data[52986] <= 8'h10 ;
			data[52987] <= 8'h10 ;
			data[52988] <= 8'h10 ;
			data[52989] <= 8'h10 ;
			data[52990] <= 8'h10 ;
			data[52991] <= 8'h10 ;
			data[52992] <= 8'h10 ;
			data[52993] <= 8'h10 ;
			data[52994] <= 8'h10 ;
			data[52995] <= 8'h10 ;
			data[52996] <= 8'h10 ;
			data[52997] <= 8'h10 ;
			data[52998] <= 8'h10 ;
			data[52999] <= 8'h10 ;
			data[53000] <= 8'h10 ;
			data[53001] <= 8'h10 ;
			data[53002] <= 8'h10 ;
			data[53003] <= 8'h10 ;
			data[53004] <= 8'h10 ;
			data[53005] <= 8'h10 ;
			data[53006] <= 8'h10 ;
			data[53007] <= 8'h10 ;
			data[53008] <= 8'h10 ;
			data[53009] <= 8'h10 ;
			data[53010] <= 8'h10 ;
			data[53011] <= 8'h10 ;
			data[53012] <= 8'h10 ;
			data[53013] <= 8'h10 ;
			data[53014] <= 8'h10 ;
			data[53015] <= 8'h10 ;
			data[53016] <= 8'h10 ;
			data[53017] <= 8'h10 ;
			data[53018] <= 8'h10 ;
			data[53019] <= 8'h10 ;
			data[53020] <= 8'h10 ;
			data[53021] <= 8'h10 ;
			data[53022] <= 8'h10 ;
			data[53023] <= 8'h10 ;
			data[53024] <= 8'h10 ;
			data[53025] <= 8'h10 ;
			data[53026] <= 8'h10 ;
			data[53027] <= 8'h10 ;
			data[53028] <= 8'h10 ;
			data[53029] <= 8'h10 ;
			data[53030] <= 8'h10 ;
			data[53031] <= 8'h10 ;
			data[53032] <= 8'h10 ;
			data[53033] <= 8'h10 ;
			data[53034] <= 8'h10 ;
			data[53035] <= 8'h10 ;
			data[53036] <= 8'h10 ;
			data[53037] <= 8'h10 ;
			data[53038] <= 8'h10 ;
			data[53039] <= 8'h10 ;
			data[53040] <= 8'h10 ;
			data[53041] <= 8'h10 ;
			data[53042] <= 8'h10 ;
			data[53043] <= 8'h10 ;
			data[53044] <= 8'h10 ;
			data[53045] <= 8'h10 ;
			data[53046] <= 8'h10 ;
			data[53047] <= 8'h10 ;
			data[53048] <= 8'h10 ;
			data[53049] <= 8'h10 ;
			data[53050] <= 8'h10 ;
			data[53051] <= 8'h10 ;
			data[53052] <= 8'h10 ;
			data[53053] <= 8'h10 ;
			data[53054] <= 8'h10 ;
			data[53055] <= 8'h10 ;
			data[53056] <= 8'h10 ;
			data[53057] <= 8'h10 ;
			data[53058] <= 8'h10 ;
			data[53059] <= 8'h10 ;
			data[53060] <= 8'h10 ;
			data[53061] <= 8'h10 ;
			data[53062] <= 8'h10 ;
			data[53063] <= 8'h10 ;
			data[53064] <= 8'h10 ;
			data[53065] <= 8'h10 ;
			data[53066] <= 8'h10 ;
			data[53067] <= 8'h10 ;
			data[53068] <= 8'h10 ;
			data[53069] <= 8'h10 ;
			data[53070] <= 8'h10 ;
			data[53071] <= 8'h10 ;
			data[53072] <= 8'h10 ;
			data[53073] <= 8'h10 ;
			data[53074] <= 8'h10 ;
			data[53075] <= 8'h10 ;
			data[53076] <= 8'h10 ;
			data[53077] <= 8'h10 ;
			data[53078] <= 8'h10 ;
			data[53079] <= 8'h10 ;
			data[53080] <= 8'h10 ;
			data[53081] <= 8'h10 ;
			data[53082] <= 8'h10 ;
			data[53083] <= 8'h10 ;
			data[53084] <= 8'h10 ;
			data[53085] <= 8'h10 ;
			data[53086] <= 8'h10 ;
			data[53087] <= 8'h10 ;
			data[53088] <= 8'h10 ;
			data[53089] <= 8'h10 ;
			data[53090] <= 8'h10 ;
			data[53091] <= 8'h10 ;
			data[53092] <= 8'h10 ;
			data[53093] <= 8'h10 ;
			data[53094] <= 8'h10 ;
			data[53095] <= 8'h10 ;
			data[53096] <= 8'h10 ;
			data[53097] <= 8'h10 ;
			data[53098] <= 8'h10 ;
			data[53099] <= 8'h10 ;
			data[53100] <= 8'h10 ;
			data[53101] <= 8'h10 ;
			data[53102] <= 8'h10 ;
			data[53103] <= 8'h10 ;
			data[53104] <= 8'h10 ;
			data[53105] <= 8'h10 ;
			data[53106] <= 8'h10 ;
			data[53107] <= 8'h10 ;
			data[53108] <= 8'h10 ;
			data[53109] <= 8'h10 ;
			data[53110] <= 8'h10 ;
			data[53111] <= 8'h10 ;
			data[53112] <= 8'h10 ;
			data[53113] <= 8'h10 ;
			data[53114] <= 8'h10 ;
			data[53115] <= 8'h10 ;
			data[53116] <= 8'h10 ;
			data[53117] <= 8'h10 ;
			data[53118] <= 8'h10 ;
			data[53119] <= 8'h10 ;
			data[53120] <= 8'h10 ;
			data[53121] <= 8'h10 ;
			data[53122] <= 8'h10 ;
			data[53123] <= 8'h10 ;
			data[53124] <= 8'h10 ;
			data[53125] <= 8'h10 ;
			data[53126] <= 8'h10 ;
			data[53127] <= 8'h10 ;
			data[53128] <= 8'h10 ;
			data[53129] <= 8'h10 ;
			data[53130] <= 8'h10 ;
			data[53131] <= 8'h10 ;
			data[53132] <= 8'h10 ;
			data[53133] <= 8'h10 ;
			data[53134] <= 8'h10 ;
			data[53135] <= 8'h10 ;
			data[53136] <= 8'h10 ;
			data[53137] <= 8'h10 ;
			data[53138] <= 8'h10 ;
			data[53139] <= 8'h10 ;
			data[53140] <= 8'h10 ;
			data[53141] <= 8'h10 ;
			data[53142] <= 8'h10 ;
			data[53143] <= 8'h10 ;
			data[53144] <= 8'h10 ;
			data[53145] <= 8'h10 ;
			data[53146] <= 8'h10 ;
			data[53147] <= 8'h10 ;
			data[53148] <= 8'h10 ;
			data[53149] <= 8'h10 ;
			data[53150] <= 8'h10 ;
			data[53151] <= 8'h10 ;
			data[53152] <= 8'h10 ;
			data[53153] <= 8'h10 ;
			data[53154] <= 8'h10 ;
			data[53155] <= 8'h10 ;
			data[53156] <= 8'h10 ;
			data[53157] <= 8'h10 ;
			data[53158] <= 8'h10 ;
			data[53159] <= 8'h10 ;
			data[53160] <= 8'h10 ;
			data[53161] <= 8'h10 ;
			data[53162] <= 8'h10 ;
			data[53163] <= 8'h10 ;
			data[53164] <= 8'h10 ;
			data[53165] <= 8'h10 ;
			data[53166] <= 8'h10 ;
			data[53167] <= 8'h10 ;
			data[53168] <= 8'h10 ;
			data[53169] <= 8'h10 ;
			data[53170] <= 8'h10 ;
			data[53171] <= 8'h10 ;
			data[53172] <= 8'h10 ;
			data[53173] <= 8'h10 ;
			data[53174] <= 8'h10 ;
			data[53175] <= 8'h10 ;
			data[53176] <= 8'h10 ;
			data[53177] <= 8'h10 ;
			data[53178] <= 8'h10 ;
			data[53179] <= 8'h10 ;
			data[53180] <= 8'h10 ;
			data[53181] <= 8'h10 ;
			data[53182] <= 8'h10 ;
			data[53183] <= 8'h10 ;
			data[53184] <= 8'h10 ;
			data[53185] <= 8'h10 ;
			data[53186] <= 8'h10 ;
			data[53187] <= 8'h10 ;
			data[53188] <= 8'h10 ;
			data[53189] <= 8'h10 ;
			data[53190] <= 8'h10 ;
			data[53191] <= 8'h10 ;
			data[53192] <= 8'h10 ;
			data[53193] <= 8'h10 ;
			data[53194] <= 8'h10 ;
			data[53195] <= 8'h10 ;
			data[53196] <= 8'h10 ;
			data[53197] <= 8'h10 ;
			data[53198] <= 8'h10 ;
			data[53199] <= 8'h10 ;
			data[53200] <= 8'h10 ;
			data[53201] <= 8'h10 ;
			data[53202] <= 8'h10 ;
			data[53203] <= 8'h10 ;
			data[53204] <= 8'h10 ;
			data[53205] <= 8'h10 ;
			data[53206] <= 8'h10 ;
			data[53207] <= 8'h10 ;
			data[53208] <= 8'h10 ;
			data[53209] <= 8'h10 ;
			data[53210] <= 8'h10 ;
			data[53211] <= 8'h10 ;
			data[53212] <= 8'h10 ;
			data[53213] <= 8'h10 ;
			data[53214] <= 8'h10 ;
			data[53215] <= 8'h10 ;
			data[53216] <= 8'h10 ;
			data[53217] <= 8'h10 ;
			data[53218] <= 8'h10 ;
			data[53219] <= 8'h10 ;
			data[53220] <= 8'h10 ;
			data[53221] <= 8'h10 ;
			data[53222] <= 8'h10 ;
			data[53223] <= 8'h10 ;
			data[53224] <= 8'h10 ;
			data[53225] <= 8'h10 ;
			data[53226] <= 8'h10 ;
			data[53227] <= 8'h10 ;
			data[53228] <= 8'h10 ;
			data[53229] <= 8'h10 ;
			data[53230] <= 8'h10 ;
			data[53231] <= 8'h10 ;
			data[53232] <= 8'h10 ;
			data[53233] <= 8'h10 ;
			data[53234] <= 8'h10 ;
			data[53235] <= 8'h10 ;
			data[53236] <= 8'h10 ;
			data[53237] <= 8'h10 ;
			data[53238] <= 8'h10 ;
			data[53239] <= 8'h10 ;
			data[53240] <= 8'h10 ;
			data[53241] <= 8'h10 ;
			data[53242] <= 8'h10 ;
			data[53243] <= 8'h10 ;
			data[53244] <= 8'h10 ;
			data[53245] <= 8'h10 ;
			data[53246] <= 8'h10 ;
			data[53247] <= 8'h10 ;
			data[53248] <= 8'h10 ;
			data[53249] <= 8'h10 ;
			data[53250] <= 8'h10 ;
			data[53251] <= 8'h10 ;
			data[53252] <= 8'h10 ;
			data[53253] <= 8'h10 ;
			data[53254] <= 8'h10 ;
			data[53255] <= 8'h10 ;
			data[53256] <= 8'h10 ;
			data[53257] <= 8'h10 ;
			data[53258] <= 8'h10 ;
			data[53259] <= 8'h10 ;
			data[53260] <= 8'h10 ;
			data[53261] <= 8'h10 ;
			data[53262] <= 8'h10 ;
			data[53263] <= 8'h10 ;
			data[53264] <= 8'h10 ;
			data[53265] <= 8'h10 ;
			data[53266] <= 8'h10 ;
			data[53267] <= 8'h10 ;
			data[53268] <= 8'h10 ;
			data[53269] <= 8'h10 ;
			data[53270] <= 8'h10 ;
			data[53271] <= 8'h10 ;
			data[53272] <= 8'h10 ;
			data[53273] <= 8'h10 ;
			data[53274] <= 8'h10 ;
			data[53275] <= 8'h10 ;
			data[53276] <= 8'h10 ;
			data[53277] <= 8'h10 ;
			data[53278] <= 8'h10 ;
			data[53279] <= 8'h10 ;
			data[53280] <= 8'h10 ;
			data[53281] <= 8'h10 ;
			data[53282] <= 8'h10 ;
			data[53283] <= 8'h10 ;
			data[53284] <= 8'h10 ;
			data[53285] <= 8'h10 ;
			data[53286] <= 8'h10 ;
			data[53287] <= 8'h10 ;
			data[53288] <= 8'h10 ;
			data[53289] <= 8'h10 ;
			data[53290] <= 8'h10 ;
			data[53291] <= 8'h10 ;
			data[53292] <= 8'h10 ;
			data[53293] <= 8'h10 ;
			data[53294] <= 8'h10 ;
			data[53295] <= 8'h10 ;
			data[53296] <= 8'h10 ;
			data[53297] <= 8'h10 ;
			data[53298] <= 8'h10 ;
			data[53299] <= 8'h10 ;
			data[53300] <= 8'h10 ;
			data[53301] <= 8'h10 ;
			data[53302] <= 8'h10 ;
			data[53303] <= 8'h10 ;
			data[53304] <= 8'h10 ;
			data[53305] <= 8'h10 ;
			data[53306] <= 8'h10 ;
			data[53307] <= 8'h10 ;
			data[53308] <= 8'h10 ;
			data[53309] <= 8'h10 ;
			data[53310] <= 8'h10 ;
			data[53311] <= 8'h10 ;
			data[53312] <= 8'h10 ;
			data[53313] <= 8'h10 ;
			data[53314] <= 8'h10 ;
			data[53315] <= 8'h10 ;
			data[53316] <= 8'h10 ;
			data[53317] <= 8'h10 ;
			data[53318] <= 8'h10 ;
			data[53319] <= 8'h10 ;
			data[53320] <= 8'h10 ;
			data[53321] <= 8'h10 ;
			data[53322] <= 8'h10 ;
			data[53323] <= 8'h10 ;
			data[53324] <= 8'h10 ;
			data[53325] <= 8'h10 ;
			data[53326] <= 8'h10 ;
			data[53327] <= 8'h10 ;
			data[53328] <= 8'h10 ;
			data[53329] <= 8'h10 ;
			data[53330] <= 8'h10 ;
			data[53331] <= 8'h10 ;
			data[53332] <= 8'h10 ;
			data[53333] <= 8'h10 ;
			data[53334] <= 8'h10 ;
			data[53335] <= 8'h10 ;
			data[53336] <= 8'h10 ;
			data[53337] <= 8'h10 ;
			data[53338] <= 8'h10 ;
			data[53339] <= 8'h10 ;
			data[53340] <= 8'h10 ;
			data[53341] <= 8'h10 ;
			data[53342] <= 8'h10 ;
			data[53343] <= 8'h10 ;
			data[53344] <= 8'h10 ;
			data[53345] <= 8'h10 ;
			data[53346] <= 8'h10 ;
			data[53347] <= 8'h10 ;
			data[53348] <= 8'h10 ;
			data[53349] <= 8'h10 ;
			data[53350] <= 8'h10 ;
			data[53351] <= 8'h10 ;
			data[53352] <= 8'h10 ;
			data[53353] <= 8'h10 ;
			data[53354] <= 8'h10 ;
			data[53355] <= 8'h10 ;
			data[53356] <= 8'h10 ;
			data[53357] <= 8'h10 ;
			data[53358] <= 8'h10 ;
			data[53359] <= 8'h10 ;
			data[53360] <= 8'h10 ;
			data[53361] <= 8'h10 ;
			data[53362] <= 8'h10 ;
			data[53363] <= 8'h10 ;
			data[53364] <= 8'h10 ;
			data[53365] <= 8'h10 ;
			data[53366] <= 8'h10 ;
			data[53367] <= 8'h10 ;
			data[53368] <= 8'h10 ;
			data[53369] <= 8'h10 ;
			data[53370] <= 8'h10 ;
			data[53371] <= 8'h10 ;
			data[53372] <= 8'h10 ;
			data[53373] <= 8'h10 ;
			data[53374] <= 8'h10 ;
			data[53375] <= 8'h10 ;
			data[53376] <= 8'h10 ;
			data[53377] <= 8'h10 ;
			data[53378] <= 8'h10 ;
			data[53379] <= 8'h10 ;
			data[53380] <= 8'h10 ;
			data[53381] <= 8'h10 ;
			data[53382] <= 8'h10 ;
			data[53383] <= 8'h10 ;
			data[53384] <= 8'h10 ;
			data[53385] <= 8'h10 ;
			data[53386] <= 8'h10 ;
			data[53387] <= 8'h10 ;
			data[53388] <= 8'h10 ;
			data[53389] <= 8'h10 ;
			data[53390] <= 8'h10 ;
			data[53391] <= 8'h10 ;
			data[53392] <= 8'h10 ;
			data[53393] <= 8'h10 ;
			data[53394] <= 8'h10 ;
			data[53395] <= 8'h10 ;
			data[53396] <= 8'h10 ;
			data[53397] <= 8'h10 ;
			data[53398] <= 8'h10 ;
			data[53399] <= 8'h10 ;
			data[53400] <= 8'h10 ;
			data[53401] <= 8'h10 ;
			data[53402] <= 8'h10 ;
			data[53403] <= 8'h10 ;
			data[53404] <= 8'h10 ;
			data[53405] <= 8'h10 ;
			data[53406] <= 8'h10 ;
			data[53407] <= 8'h10 ;
			data[53408] <= 8'h10 ;
			data[53409] <= 8'h10 ;
			data[53410] <= 8'h10 ;
			data[53411] <= 8'h10 ;
			data[53412] <= 8'h10 ;
			data[53413] <= 8'h10 ;
			data[53414] <= 8'h10 ;
			data[53415] <= 8'h10 ;
			data[53416] <= 8'h10 ;
			data[53417] <= 8'h10 ;
			data[53418] <= 8'h10 ;
			data[53419] <= 8'h10 ;
			data[53420] <= 8'h10 ;
			data[53421] <= 8'h10 ;
			data[53422] <= 8'h10 ;
			data[53423] <= 8'h10 ;
			data[53424] <= 8'h10 ;
			data[53425] <= 8'h10 ;
			data[53426] <= 8'h10 ;
			data[53427] <= 8'h10 ;
			data[53428] <= 8'h10 ;
			data[53429] <= 8'h10 ;
			data[53430] <= 8'h10 ;
			data[53431] <= 8'h10 ;
			data[53432] <= 8'h10 ;
			data[53433] <= 8'h10 ;
			data[53434] <= 8'h10 ;
			data[53435] <= 8'h10 ;
			data[53436] <= 8'h10 ;
			data[53437] <= 8'h10 ;
			data[53438] <= 8'h10 ;
			data[53439] <= 8'h10 ;
			data[53440] <= 8'h10 ;
			data[53441] <= 8'h10 ;
			data[53442] <= 8'h10 ;
			data[53443] <= 8'h10 ;
			data[53444] <= 8'h10 ;
			data[53445] <= 8'h10 ;
			data[53446] <= 8'h10 ;
			data[53447] <= 8'h10 ;
			data[53448] <= 8'h10 ;
			data[53449] <= 8'h10 ;
			data[53450] <= 8'h10 ;
			data[53451] <= 8'h10 ;
			data[53452] <= 8'h10 ;
			data[53453] <= 8'h10 ;
			data[53454] <= 8'h10 ;
			data[53455] <= 8'h10 ;
			data[53456] <= 8'h10 ;
			data[53457] <= 8'h10 ;
			data[53458] <= 8'h10 ;
			data[53459] <= 8'h10 ;
			data[53460] <= 8'h10 ;
			data[53461] <= 8'h10 ;
			data[53462] <= 8'h10 ;
			data[53463] <= 8'h10 ;
			data[53464] <= 8'h10 ;
			data[53465] <= 8'h10 ;
			data[53466] <= 8'h10 ;
			data[53467] <= 8'h10 ;
			data[53468] <= 8'h10 ;
			data[53469] <= 8'h10 ;
			data[53470] <= 8'h10 ;
			data[53471] <= 8'h10 ;
			data[53472] <= 8'h10 ;
			data[53473] <= 8'h10 ;
			data[53474] <= 8'h10 ;
			data[53475] <= 8'h10 ;
			data[53476] <= 8'h10 ;
			data[53477] <= 8'h10 ;
			data[53478] <= 8'h10 ;
			data[53479] <= 8'h10 ;
			data[53480] <= 8'h10 ;
			data[53481] <= 8'h10 ;
			data[53482] <= 8'h10 ;
			data[53483] <= 8'h10 ;
			data[53484] <= 8'h10 ;
			data[53485] <= 8'h10 ;
			data[53486] <= 8'h10 ;
			data[53487] <= 8'h10 ;
			data[53488] <= 8'h10 ;
			data[53489] <= 8'h10 ;
			data[53490] <= 8'h10 ;
			data[53491] <= 8'h10 ;
			data[53492] <= 8'h10 ;
			data[53493] <= 8'h10 ;
			data[53494] <= 8'h10 ;
			data[53495] <= 8'h10 ;
			data[53496] <= 8'h10 ;
			data[53497] <= 8'h10 ;
			data[53498] <= 8'h10 ;
			data[53499] <= 8'h10 ;
			data[53500] <= 8'h10 ;
			data[53501] <= 8'h10 ;
			data[53502] <= 8'h10 ;
			data[53503] <= 8'h10 ;
			data[53504] <= 8'h10 ;
			data[53505] <= 8'h10 ;
			data[53506] <= 8'h10 ;
			data[53507] <= 8'h10 ;
			data[53508] <= 8'h10 ;
			data[53509] <= 8'h10 ;
			data[53510] <= 8'h10 ;
			data[53511] <= 8'h10 ;
			data[53512] <= 8'h10 ;
			data[53513] <= 8'h10 ;
			data[53514] <= 8'h10 ;
			data[53515] <= 8'h10 ;
			data[53516] <= 8'h10 ;
			data[53517] <= 8'h10 ;
			data[53518] <= 8'h10 ;
			data[53519] <= 8'h10 ;
			data[53520] <= 8'h10 ;
			data[53521] <= 8'h10 ;
			data[53522] <= 8'h10 ;
			data[53523] <= 8'h10 ;
			data[53524] <= 8'h10 ;
			data[53525] <= 8'h10 ;
			data[53526] <= 8'h10 ;
			data[53527] <= 8'h10 ;
			data[53528] <= 8'h10 ;
			data[53529] <= 8'h10 ;
			data[53530] <= 8'h10 ;
			data[53531] <= 8'h10 ;
			data[53532] <= 8'h10 ;
			data[53533] <= 8'h10 ;
			data[53534] <= 8'h10 ;
			data[53535] <= 8'h10 ;
			data[53536] <= 8'h10 ;
			data[53537] <= 8'h10 ;
			data[53538] <= 8'h10 ;
			data[53539] <= 8'h10 ;
			data[53540] <= 8'h10 ;
			data[53541] <= 8'h10 ;
			data[53542] <= 8'h10 ;
			data[53543] <= 8'h10 ;
			data[53544] <= 8'h10 ;
			data[53545] <= 8'h10 ;
			data[53546] <= 8'h10 ;
			data[53547] <= 8'h10 ;
			data[53548] <= 8'h10 ;
			data[53549] <= 8'h10 ;
			data[53550] <= 8'h10 ;
			data[53551] <= 8'h10 ;
			data[53552] <= 8'h10 ;
			data[53553] <= 8'h10 ;
			data[53554] <= 8'h10 ;
			data[53555] <= 8'h10 ;
			data[53556] <= 8'h10 ;
			data[53557] <= 8'h10 ;
			data[53558] <= 8'h10 ;
			data[53559] <= 8'h10 ;
			data[53560] <= 8'h10 ;
			data[53561] <= 8'h10 ;
			data[53562] <= 8'h10 ;
			data[53563] <= 8'h10 ;
			data[53564] <= 8'h10 ;
			data[53565] <= 8'h10 ;
			data[53566] <= 8'h10 ;
			data[53567] <= 8'h10 ;
			data[53568] <= 8'h10 ;
			data[53569] <= 8'h10 ;
			data[53570] <= 8'h10 ;
			data[53571] <= 8'h10 ;
			data[53572] <= 8'h10 ;
			data[53573] <= 8'h10 ;
			data[53574] <= 8'h10 ;
			data[53575] <= 8'h10 ;
			data[53576] <= 8'h10 ;
			data[53577] <= 8'h10 ;
			data[53578] <= 8'h10 ;
			data[53579] <= 8'h10 ;
			data[53580] <= 8'h10 ;
			data[53581] <= 8'h10 ;
			data[53582] <= 8'h10 ;
			data[53583] <= 8'h10 ;
			data[53584] <= 8'h10 ;
			data[53585] <= 8'h10 ;
			data[53586] <= 8'h10 ;
			data[53587] <= 8'h10 ;
			data[53588] <= 8'h10 ;
			data[53589] <= 8'h10 ;
			data[53590] <= 8'h10 ;
			data[53591] <= 8'h10 ;
			data[53592] <= 8'h10 ;
			data[53593] <= 8'h10 ;
			data[53594] <= 8'h10 ;
			data[53595] <= 8'h10 ;
			data[53596] <= 8'h10 ;
			data[53597] <= 8'h10 ;
			data[53598] <= 8'h10 ;
			data[53599] <= 8'h10 ;
			data[53600] <= 8'h10 ;
			data[53601] <= 8'h10 ;
			data[53602] <= 8'h10 ;
			data[53603] <= 8'h10 ;
			data[53604] <= 8'h10 ;
			data[53605] <= 8'h10 ;
			data[53606] <= 8'h10 ;
			data[53607] <= 8'h10 ;
			data[53608] <= 8'h10 ;
			data[53609] <= 8'h10 ;
			data[53610] <= 8'h10 ;
			data[53611] <= 8'h10 ;
			data[53612] <= 8'h10 ;
			data[53613] <= 8'h10 ;
			data[53614] <= 8'h10 ;
			data[53615] <= 8'h10 ;
			data[53616] <= 8'h10 ;
			data[53617] <= 8'h10 ;
			data[53618] <= 8'h10 ;
			data[53619] <= 8'h10 ;
			data[53620] <= 8'h10 ;
			data[53621] <= 8'h10 ;
			data[53622] <= 8'h10 ;
			data[53623] <= 8'h10 ;
			data[53624] <= 8'h10 ;
			data[53625] <= 8'h10 ;
			data[53626] <= 8'h10 ;
			data[53627] <= 8'h10 ;
			data[53628] <= 8'h10 ;
			data[53629] <= 8'h10 ;
			data[53630] <= 8'h10 ;
			data[53631] <= 8'h10 ;
			data[53632] <= 8'h10 ;
			data[53633] <= 8'h10 ;
			data[53634] <= 8'h10 ;
			data[53635] <= 8'h10 ;
			data[53636] <= 8'h10 ;
			data[53637] <= 8'h10 ;
			data[53638] <= 8'h10 ;
			data[53639] <= 8'h10 ;
			data[53640] <= 8'h10 ;
			data[53641] <= 8'h10 ;
			data[53642] <= 8'h10 ;
			data[53643] <= 8'h10 ;
			data[53644] <= 8'h10 ;
			data[53645] <= 8'h10 ;
			data[53646] <= 8'h10 ;
			data[53647] <= 8'h10 ;
			data[53648] <= 8'h10 ;
			data[53649] <= 8'h10 ;
			data[53650] <= 8'h10 ;
			data[53651] <= 8'h10 ;
			data[53652] <= 8'h10 ;
			data[53653] <= 8'h10 ;
			data[53654] <= 8'h10 ;
			data[53655] <= 8'h10 ;
			data[53656] <= 8'h10 ;
			data[53657] <= 8'h10 ;
			data[53658] <= 8'h10 ;
			data[53659] <= 8'h10 ;
			data[53660] <= 8'h10 ;
			data[53661] <= 8'h10 ;
			data[53662] <= 8'h10 ;
			data[53663] <= 8'h10 ;
			data[53664] <= 8'h10 ;
			data[53665] <= 8'h10 ;
			data[53666] <= 8'h10 ;
			data[53667] <= 8'h10 ;
			data[53668] <= 8'h10 ;
			data[53669] <= 8'h10 ;
			data[53670] <= 8'h10 ;
			data[53671] <= 8'h10 ;
			data[53672] <= 8'h10 ;
			data[53673] <= 8'h10 ;
			data[53674] <= 8'h10 ;
			data[53675] <= 8'h10 ;
			data[53676] <= 8'h10 ;
			data[53677] <= 8'h10 ;
			data[53678] <= 8'h10 ;
			data[53679] <= 8'h10 ;
			data[53680] <= 8'h10 ;
			data[53681] <= 8'h10 ;
			data[53682] <= 8'h10 ;
			data[53683] <= 8'h10 ;
			data[53684] <= 8'h10 ;
			data[53685] <= 8'h10 ;
			data[53686] <= 8'h10 ;
			data[53687] <= 8'h10 ;
			data[53688] <= 8'h10 ;
			data[53689] <= 8'h10 ;
			data[53690] <= 8'h10 ;
			data[53691] <= 8'h10 ;
			data[53692] <= 8'h10 ;
			data[53693] <= 8'h10 ;
			data[53694] <= 8'h10 ;
			data[53695] <= 8'h10 ;
			data[53696] <= 8'h10 ;
			data[53697] <= 8'h10 ;
			data[53698] <= 8'h10 ;
			data[53699] <= 8'h10 ;
			data[53700] <= 8'h10 ;
			data[53701] <= 8'h10 ;
			data[53702] <= 8'h10 ;
			data[53703] <= 8'h10 ;
			data[53704] <= 8'h10 ;
			data[53705] <= 8'h10 ;
			data[53706] <= 8'h10 ;
			data[53707] <= 8'h10 ;
			data[53708] <= 8'h10 ;
			data[53709] <= 8'h10 ;
			data[53710] <= 8'h10 ;
			data[53711] <= 8'h10 ;
			data[53712] <= 8'h10 ;
			data[53713] <= 8'h10 ;
			data[53714] <= 8'h10 ;
			data[53715] <= 8'h10 ;
			data[53716] <= 8'h10 ;
			data[53717] <= 8'h10 ;
			data[53718] <= 8'h10 ;
			data[53719] <= 8'h10 ;
			data[53720] <= 8'h10 ;
			data[53721] <= 8'h10 ;
			data[53722] <= 8'h10 ;
			data[53723] <= 8'h10 ;
			data[53724] <= 8'h10 ;
			data[53725] <= 8'h10 ;
			data[53726] <= 8'h10 ;
			data[53727] <= 8'h10 ;
			data[53728] <= 8'h10 ;
			data[53729] <= 8'h10 ;
			data[53730] <= 8'h10 ;
			data[53731] <= 8'h10 ;
			data[53732] <= 8'h10 ;
			data[53733] <= 8'h10 ;
			data[53734] <= 8'h10 ;
			data[53735] <= 8'h10 ;
			data[53736] <= 8'h10 ;
			data[53737] <= 8'h10 ;
			data[53738] <= 8'h10 ;
			data[53739] <= 8'h10 ;
			data[53740] <= 8'h10 ;
			data[53741] <= 8'h10 ;
			data[53742] <= 8'h10 ;
			data[53743] <= 8'h10 ;
			data[53744] <= 8'h10 ;
			data[53745] <= 8'h10 ;
			data[53746] <= 8'h10 ;
			data[53747] <= 8'h10 ;
			data[53748] <= 8'h10 ;
			data[53749] <= 8'h10 ;
			data[53750] <= 8'h10 ;
			data[53751] <= 8'h10 ;
			data[53752] <= 8'h10 ;
			data[53753] <= 8'h10 ;
			data[53754] <= 8'h10 ;
			data[53755] <= 8'h10 ;
			data[53756] <= 8'h10 ;
			data[53757] <= 8'h10 ;
			data[53758] <= 8'h10 ;
			data[53759] <= 8'h10 ;
			data[53760] <= 8'h10 ;
			data[53761] <= 8'h10 ;
			data[53762] <= 8'h10 ;
			data[53763] <= 8'h10 ;
			data[53764] <= 8'h10 ;
			data[53765] <= 8'h10 ;
			data[53766] <= 8'h10 ;
			data[53767] <= 8'h10 ;
			data[53768] <= 8'h10 ;
			data[53769] <= 8'h10 ;
			data[53770] <= 8'h10 ;
			data[53771] <= 8'h10 ;
			data[53772] <= 8'h10 ;
			data[53773] <= 8'h10 ;
			data[53774] <= 8'h10 ;
			data[53775] <= 8'h10 ;
			data[53776] <= 8'h10 ;
			data[53777] <= 8'h10 ;
			data[53778] <= 8'h10 ;
			data[53779] <= 8'h10 ;
			data[53780] <= 8'h10 ;
			data[53781] <= 8'h10 ;
			data[53782] <= 8'h10 ;
			data[53783] <= 8'h10 ;
			data[53784] <= 8'h10 ;
			data[53785] <= 8'h10 ;
			data[53786] <= 8'h10 ;
			data[53787] <= 8'h10 ;
			data[53788] <= 8'h10 ;
			data[53789] <= 8'h10 ;
			data[53790] <= 8'h10 ;
			data[53791] <= 8'h10 ;
			data[53792] <= 8'h10 ;
			data[53793] <= 8'h10 ;
			data[53794] <= 8'h10 ;
			data[53795] <= 8'h10 ;
			data[53796] <= 8'h10 ;
			data[53797] <= 8'h10 ;
			data[53798] <= 8'h10 ;
			data[53799] <= 8'h10 ;
			data[53800] <= 8'h10 ;
			data[53801] <= 8'h10 ;
			data[53802] <= 8'h10 ;
			data[53803] <= 8'h10 ;
			data[53804] <= 8'h10 ;
			data[53805] <= 8'h10 ;
			data[53806] <= 8'h10 ;
			data[53807] <= 8'h10 ;
			data[53808] <= 8'h10 ;
			data[53809] <= 8'h10 ;
			data[53810] <= 8'h10 ;
			data[53811] <= 8'h10 ;
			data[53812] <= 8'h10 ;
			data[53813] <= 8'h10 ;
			data[53814] <= 8'h10 ;
			data[53815] <= 8'h10 ;
			data[53816] <= 8'h10 ;
			data[53817] <= 8'h10 ;
			data[53818] <= 8'h10 ;
			data[53819] <= 8'h10 ;
			data[53820] <= 8'h10 ;
			data[53821] <= 8'h10 ;
			data[53822] <= 8'h10 ;
			data[53823] <= 8'h10 ;
			data[53824] <= 8'h10 ;
			data[53825] <= 8'h10 ;
			data[53826] <= 8'h10 ;
			data[53827] <= 8'h10 ;
			data[53828] <= 8'h10 ;
			data[53829] <= 8'h10 ;
			data[53830] <= 8'h10 ;
			data[53831] <= 8'h10 ;
			data[53832] <= 8'h10 ;
			data[53833] <= 8'h10 ;
			data[53834] <= 8'h10 ;
			data[53835] <= 8'h10 ;
			data[53836] <= 8'h10 ;
			data[53837] <= 8'h10 ;
			data[53838] <= 8'h10 ;
			data[53839] <= 8'h10 ;
			data[53840] <= 8'h10 ;
			data[53841] <= 8'h10 ;
			data[53842] <= 8'h10 ;
			data[53843] <= 8'h10 ;
			data[53844] <= 8'h10 ;
			data[53845] <= 8'h10 ;
			data[53846] <= 8'h10 ;
			data[53847] <= 8'h10 ;
			data[53848] <= 8'h10 ;
			data[53849] <= 8'h10 ;
			data[53850] <= 8'h10 ;
			data[53851] <= 8'h10 ;
			data[53852] <= 8'h10 ;
			data[53853] <= 8'h10 ;
			data[53854] <= 8'h10 ;
			data[53855] <= 8'h10 ;
			data[53856] <= 8'h10 ;
			data[53857] <= 8'h10 ;
			data[53858] <= 8'h10 ;
			data[53859] <= 8'h10 ;
			data[53860] <= 8'h10 ;
			data[53861] <= 8'h10 ;
			data[53862] <= 8'h10 ;
			data[53863] <= 8'h10 ;
			data[53864] <= 8'h10 ;
			data[53865] <= 8'h10 ;
			data[53866] <= 8'h10 ;
			data[53867] <= 8'h10 ;
			data[53868] <= 8'h10 ;
			data[53869] <= 8'h10 ;
			data[53870] <= 8'h10 ;
			data[53871] <= 8'h10 ;
			data[53872] <= 8'h10 ;
			data[53873] <= 8'h10 ;
			data[53874] <= 8'h10 ;
			data[53875] <= 8'h10 ;
			data[53876] <= 8'h10 ;
			data[53877] <= 8'h10 ;
			data[53878] <= 8'h10 ;
			data[53879] <= 8'h10 ;
			data[53880] <= 8'h10 ;
			data[53881] <= 8'h10 ;
			data[53882] <= 8'h10 ;
			data[53883] <= 8'h10 ;
			data[53884] <= 8'h10 ;
			data[53885] <= 8'h10 ;
			data[53886] <= 8'h10 ;
			data[53887] <= 8'h10 ;
			data[53888] <= 8'h10 ;
			data[53889] <= 8'h10 ;
			data[53890] <= 8'h10 ;
			data[53891] <= 8'h10 ;
			data[53892] <= 8'h10 ;
			data[53893] <= 8'h10 ;
			data[53894] <= 8'h10 ;
			data[53895] <= 8'h10 ;
			data[53896] <= 8'h10 ;
			data[53897] <= 8'h10 ;
			data[53898] <= 8'h10 ;
			data[53899] <= 8'h10 ;
			data[53900] <= 8'h10 ;
			data[53901] <= 8'h10 ;
			data[53902] <= 8'h10 ;
			data[53903] <= 8'h10 ;
			data[53904] <= 8'h10 ;
			data[53905] <= 8'h10 ;
			data[53906] <= 8'h10 ;
			data[53907] <= 8'h10 ;
			data[53908] <= 8'h10 ;
			data[53909] <= 8'h10 ;
			data[53910] <= 8'h10 ;
			data[53911] <= 8'h10 ;
			data[53912] <= 8'h10 ;
			data[53913] <= 8'h10 ;
			data[53914] <= 8'h10 ;
			data[53915] <= 8'h10 ;
			data[53916] <= 8'h10 ;
			data[53917] <= 8'h10 ;
			data[53918] <= 8'h10 ;
			data[53919] <= 8'h10 ;
			data[53920] <= 8'h10 ;
			data[53921] <= 8'h10 ;
			data[53922] <= 8'h10 ;
			data[53923] <= 8'h10 ;
			data[53924] <= 8'h10 ;
			data[53925] <= 8'h10 ;
			data[53926] <= 8'h10 ;
			data[53927] <= 8'h10 ;
			data[53928] <= 8'h10 ;
			data[53929] <= 8'h10 ;
			data[53930] <= 8'h10 ;
			data[53931] <= 8'h10 ;
			data[53932] <= 8'h10 ;
			data[53933] <= 8'h10 ;
			data[53934] <= 8'h10 ;
			data[53935] <= 8'h10 ;
			data[53936] <= 8'h10 ;
			data[53937] <= 8'h10 ;
			data[53938] <= 8'h10 ;
			data[53939] <= 8'h10 ;
			data[53940] <= 8'h10 ;
			data[53941] <= 8'h10 ;
			data[53942] <= 8'h10 ;
			data[53943] <= 8'h10 ;
			data[53944] <= 8'h10 ;
			data[53945] <= 8'h10 ;
			data[53946] <= 8'h10 ;
			data[53947] <= 8'h10 ;
			data[53948] <= 8'h10 ;
			data[53949] <= 8'h10 ;
			data[53950] <= 8'h10 ;
			data[53951] <= 8'h10 ;
			data[53952] <= 8'h10 ;
			data[53953] <= 8'h10 ;
			data[53954] <= 8'h10 ;
			data[53955] <= 8'h10 ;
			data[53956] <= 8'h10 ;
			data[53957] <= 8'h10 ;
			data[53958] <= 8'h10 ;
			data[53959] <= 8'h10 ;
			data[53960] <= 8'h10 ;
			data[53961] <= 8'h10 ;
			data[53962] <= 8'h10 ;
			data[53963] <= 8'h10 ;
			data[53964] <= 8'h10 ;
			data[53965] <= 8'h10 ;
			data[53966] <= 8'h10 ;
			data[53967] <= 8'h10 ;
			data[53968] <= 8'h10 ;
			data[53969] <= 8'h10 ;
			data[53970] <= 8'h10 ;
			data[53971] <= 8'h10 ;
			data[53972] <= 8'h10 ;
			data[53973] <= 8'h10 ;
			data[53974] <= 8'h10 ;
			data[53975] <= 8'h10 ;
			data[53976] <= 8'h10 ;
			data[53977] <= 8'h10 ;
			data[53978] <= 8'h10 ;
			data[53979] <= 8'h10 ;
			data[53980] <= 8'h10 ;
			data[53981] <= 8'h10 ;
			data[53982] <= 8'h10 ;
			data[53983] <= 8'h10 ;
			data[53984] <= 8'h10 ;
			data[53985] <= 8'h10 ;
			data[53986] <= 8'h10 ;
			data[53987] <= 8'h10 ;
			data[53988] <= 8'h10 ;
			data[53989] <= 8'h10 ;
			data[53990] <= 8'h10 ;
			data[53991] <= 8'h10 ;
			data[53992] <= 8'h10 ;
			data[53993] <= 8'h10 ;
			data[53994] <= 8'h10 ;
			data[53995] <= 8'h10 ;
			data[53996] <= 8'h10 ;
			data[53997] <= 8'h10 ;
			data[53998] <= 8'h10 ;
			data[53999] <= 8'h10 ;
			data[54000] <= 8'h10 ;
			data[54001] <= 8'h10 ;
			data[54002] <= 8'h10 ;
			data[54003] <= 8'h10 ;
			data[54004] <= 8'h10 ;
			data[54005] <= 8'h10 ;
			data[54006] <= 8'h10 ;
			data[54007] <= 8'h10 ;
			data[54008] <= 8'h10 ;
			data[54009] <= 8'h10 ;
			data[54010] <= 8'h10 ;
			data[54011] <= 8'h10 ;
			data[54012] <= 8'h10 ;
			data[54013] <= 8'h10 ;
			data[54014] <= 8'h10 ;
			data[54015] <= 8'h10 ;
			data[54016] <= 8'h10 ;
			data[54017] <= 8'h10 ;
			data[54018] <= 8'h10 ;
			data[54019] <= 8'h10 ;
			data[54020] <= 8'h10 ;
			data[54021] <= 8'h10 ;
			data[54022] <= 8'h10 ;
			data[54023] <= 8'h10 ;
			data[54024] <= 8'h10 ;
			data[54025] <= 8'h10 ;
			data[54026] <= 8'h10 ;
			data[54027] <= 8'h10 ;
			data[54028] <= 8'h10 ;
			data[54029] <= 8'h10 ;
			data[54030] <= 8'h10 ;
			data[54031] <= 8'h10 ;
			data[54032] <= 8'h10 ;
			data[54033] <= 8'h10 ;
			data[54034] <= 8'h10 ;
			data[54035] <= 8'h10 ;
			data[54036] <= 8'h10 ;
			data[54037] <= 8'h10 ;
			data[54038] <= 8'h10 ;
			data[54039] <= 8'h10 ;
			data[54040] <= 8'h10 ;
			data[54041] <= 8'h10 ;
			data[54042] <= 8'h10 ;
			data[54043] <= 8'h10 ;
			data[54044] <= 8'h10 ;
			data[54045] <= 8'h10 ;
			data[54046] <= 8'h10 ;
			data[54047] <= 8'h10 ;
			data[54048] <= 8'h10 ;
			data[54049] <= 8'h10 ;
			data[54050] <= 8'h10 ;
			data[54051] <= 8'h10 ;
			data[54052] <= 8'h10 ;
			data[54053] <= 8'h10 ;
			data[54054] <= 8'h10 ;
			data[54055] <= 8'h10 ;
			data[54056] <= 8'h10 ;
			data[54057] <= 8'h10 ;
			data[54058] <= 8'h10 ;
			data[54059] <= 8'h10 ;
			data[54060] <= 8'h10 ;
			data[54061] <= 8'h10 ;
			data[54062] <= 8'h10 ;
			data[54063] <= 8'h10 ;
			data[54064] <= 8'h10 ;
			data[54065] <= 8'h10 ;
			data[54066] <= 8'h10 ;
			data[54067] <= 8'h10 ;
			data[54068] <= 8'h10 ;
			data[54069] <= 8'h10 ;
			data[54070] <= 8'h10 ;
			data[54071] <= 8'h10 ;
			data[54072] <= 8'h10 ;
			data[54073] <= 8'h10 ;
			data[54074] <= 8'h10 ;
			data[54075] <= 8'h10 ;
			data[54076] <= 8'h10 ;
			data[54077] <= 8'h10 ;
			data[54078] <= 8'h10 ;
			data[54079] <= 8'h10 ;
			data[54080] <= 8'h10 ;
			data[54081] <= 8'h10 ;
			data[54082] <= 8'h10 ;
			data[54083] <= 8'h10 ;
			data[54084] <= 8'h10 ;
			data[54085] <= 8'h10 ;
			data[54086] <= 8'h10 ;
			data[54087] <= 8'h10 ;
			data[54088] <= 8'h10 ;
			data[54089] <= 8'h10 ;
			data[54090] <= 8'h10 ;
			data[54091] <= 8'h10 ;
			data[54092] <= 8'h10 ;
			data[54093] <= 8'h10 ;
			data[54094] <= 8'h10 ;
			data[54095] <= 8'h10 ;
			data[54096] <= 8'h10 ;
			data[54097] <= 8'h10 ;
			data[54098] <= 8'h10 ;
			data[54099] <= 8'h10 ;
			data[54100] <= 8'h10 ;
			data[54101] <= 8'h10 ;
			data[54102] <= 8'h10 ;
			data[54103] <= 8'h10 ;
			data[54104] <= 8'h10 ;
			data[54105] <= 8'h10 ;
			data[54106] <= 8'h10 ;
			data[54107] <= 8'h10 ;
			data[54108] <= 8'h10 ;
			data[54109] <= 8'h10 ;
			data[54110] <= 8'h10 ;
			data[54111] <= 8'h10 ;
			data[54112] <= 8'h10 ;
			data[54113] <= 8'h10 ;
			data[54114] <= 8'h10 ;
			data[54115] <= 8'h10 ;
			data[54116] <= 8'h10 ;
			data[54117] <= 8'h10 ;
			data[54118] <= 8'h10 ;
			data[54119] <= 8'h10 ;
			data[54120] <= 8'h10 ;
			data[54121] <= 8'h10 ;
			data[54122] <= 8'h10 ;
			data[54123] <= 8'h10 ;
			data[54124] <= 8'h10 ;
			data[54125] <= 8'h10 ;
			data[54126] <= 8'h10 ;
			data[54127] <= 8'h10 ;
			data[54128] <= 8'h10 ;
			data[54129] <= 8'h10 ;
			data[54130] <= 8'h10 ;
			data[54131] <= 8'h10 ;
			data[54132] <= 8'h10 ;
			data[54133] <= 8'h10 ;
			data[54134] <= 8'h10 ;
			data[54135] <= 8'h10 ;
			data[54136] <= 8'h10 ;
			data[54137] <= 8'h10 ;
			data[54138] <= 8'h10 ;
			data[54139] <= 8'h10 ;
			data[54140] <= 8'h10 ;
			data[54141] <= 8'h10 ;
			data[54142] <= 8'h10 ;
			data[54143] <= 8'h10 ;
			data[54144] <= 8'h10 ;
			data[54145] <= 8'h10 ;
			data[54146] <= 8'h10 ;
			data[54147] <= 8'h10 ;
			data[54148] <= 8'h10 ;
			data[54149] <= 8'h10 ;
			data[54150] <= 8'h10 ;
			data[54151] <= 8'h10 ;
			data[54152] <= 8'h10 ;
			data[54153] <= 8'h10 ;
			data[54154] <= 8'h10 ;
			data[54155] <= 8'h10 ;
			data[54156] <= 8'h10 ;
			data[54157] <= 8'h10 ;
			data[54158] <= 8'h10 ;
			data[54159] <= 8'h10 ;
			data[54160] <= 8'h10 ;
			data[54161] <= 8'h10 ;
			data[54162] <= 8'h10 ;
			data[54163] <= 8'h10 ;
			data[54164] <= 8'h10 ;
			data[54165] <= 8'h10 ;
			data[54166] <= 8'h10 ;
			data[54167] <= 8'h10 ;
			data[54168] <= 8'h10 ;
			data[54169] <= 8'h10 ;
			data[54170] <= 8'h10 ;
			data[54171] <= 8'h10 ;
			data[54172] <= 8'h10 ;
			data[54173] <= 8'h10 ;
			data[54174] <= 8'h10 ;
			data[54175] <= 8'h10 ;
			data[54176] <= 8'h10 ;
			data[54177] <= 8'h10 ;
			data[54178] <= 8'h10 ;
			data[54179] <= 8'h10 ;
			data[54180] <= 8'h10 ;
			data[54181] <= 8'h10 ;
			data[54182] <= 8'h10 ;
			data[54183] <= 8'h10 ;
			data[54184] <= 8'h10 ;
			data[54185] <= 8'h10 ;
			data[54186] <= 8'h10 ;
			data[54187] <= 8'h10 ;
			data[54188] <= 8'h10 ;
			data[54189] <= 8'h10 ;
			data[54190] <= 8'h10 ;
			data[54191] <= 8'h10 ;
			data[54192] <= 8'h10 ;
			data[54193] <= 8'h10 ;
			data[54194] <= 8'h10 ;
			data[54195] <= 8'h10 ;
			data[54196] <= 8'h10 ;
			data[54197] <= 8'h10 ;
			data[54198] <= 8'h10 ;
			data[54199] <= 8'h10 ;
			data[54200] <= 8'h10 ;
			data[54201] <= 8'h10 ;
			data[54202] <= 8'h10 ;
			data[54203] <= 8'h10 ;
			data[54204] <= 8'h10 ;
			data[54205] <= 8'h10 ;
			data[54206] <= 8'h10 ;
			data[54207] <= 8'h10 ;
			data[54208] <= 8'h10 ;
			data[54209] <= 8'h10 ;
			data[54210] <= 8'h10 ;
			data[54211] <= 8'h10 ;
			data[54212] <= 8'h10 ;
			data[54213] <= 8'h10 ;
			data[54214] <= 8'h10 ;
			data[54215] <= 8'h10 ;
			data[54216] <= 8'h10 ;
			data[54217] <= 8'h10 ;
			data[54218] <= 8'h10 ;
			data[54219] <= 8'h10 ;
			data[54220] <= 8'h10 ;
			data[54221] <= 8'h10 ;
			data[54222] <= 8'h10 ;
			data[54223] <= 8'h10 ;
			data[54224] <= 8'h10 ;
			data[54225] <= 8'h10 ;
			data[54226] <= 8'h10 ;
			data[54227] <= 8'h10 ;
			data[54228] <= 8'h10 ;
			data[54229] <= 8'h10 ;
			data[54230] <= 8'h10 ;
			data[54231] <= 8'h10 ;
			data[54232] <= 8'h10 ;
			data[54233] <= 8'h10 ;
			data[54234] <= 8'h10 ;
			data[54235] <= 8'h10 ;
			data[54236] <= 8'h10 ;
			data[54237] <= 8'h10 ;
			data[54238] <= 8'h10 ;
			data[54239] <= 8'h10 ;
			data[54240] <= 8'h10 ;
			data[54241] <= 8'h10 ;
			data[54242] <= 8'h10 ;
			data[54243] <= 8'h10 ;
			data[54244] <= 8'h10 ;
			data[54245] <= 8'h10 ;
			data[54246] <= 8'h10 ;
			data[54247] <= 8'h10 ;
			data[54248] <= 8'h10 ;
			data[54249] <= 8'h10 ;
			data[54250] <= 8'h10 ;
			data[54251] <= 8'h10 ;
			data[54252] <= 8'h10 ;
			data[54253] <= 8'h10 ;
			data[54254] <= 8'h10 ;
			data[54255] <= 8'h10 ;
			data[54256] <= 8'h10 ;
			data[54257] <= 8'h10 ;
			data[54258] <= 8'h10 ;
			data[54259] <= 8'h10 ;
			data[54260] <= 8'h10 ;
			data[54261] <= 8'h10 ;
			data[54262] <= 8'h10 ;
			data[54263] <= 8'h10 ;
			data[54264] <= 8'h10 ;
			data[54265] <= 8'h10 ;
			data[54266] <= 8'h10 ;
			data[54267] <= 8'h10 ;
			data[54268] <= 8'h10 ;
			data[54269] <= 8'h10 ;
			data[54270] <= 8'h10 ;
			data[54271] <= 8'h10 ;
			data[54272] <= 8'h10 ;
			data[54273] <= 8'h10 ;
			data[54274] <= 8'h10 ;
			data[54275] <= 8'h10 ;
			data[54276] <= 8'h10 ;
			data[54277] <= 8'h10 ;
			data[54278] <= 8'h10 ;
			data[54279] <= 8'h10 ;
			data[54280] <= 8'h10 ;
			data[54281] <= 8'h10 ;
			data[54282] <= 8'h10 ;
			data[54283] <= 8'h10 ;
			data[54284] <= 8'h10 ;
			data[54285] <= 8'h10 ;
			data[54286] <= 8'h10 ;
			data[54287] <= 8'h10 ;
			data[54288] <= 8'h10 ;
			data[54289] <= 8'h10 ;
			data[54290] <= 8'h10 ;
			data[54291] <= 8'h10 ;
			data[54292] <= 8'h10 ;
			data[54293] <= 8'h10 ;
			data[54294] <= 8'h10 ;
			data[54295] <= 8'h10 ;
			data[54296] <= 8'h10 ;
			data[54297] <= 8'h10 ;
			data[54298] <= 8'h10 ;
			data[54299] <= 8'h10 ;
			data[54300] <= 8'h10 ;
			data[54301] <= 8'h10 ;
			data[54302] <= 8'h10 ;
			data[54303] <= 8'h10 ;
			data[54304] <= 8'h10 ;
			data[54305] <= 8'h10 ;
			data[54306] <= 8'h10 ;
			data[54307] <= 8'h10 ;
			data[54308] <= 8'h10 ;
			data[54309] <= 8'h10 ;
			data[54310] <= 8'h10 ;
			data[54311] <= 8'h10 ;
			data[54312] <= 8'h10 ;
			data[54313] <= 8'h10 ;
			data[54314] <= 8'h10 ;
			data[54315] <= 8'h10 ;
			data[54316] <= 8'h10 ;
			data[54317] <= 8'h10 ;
			data[54318] <= 8'h10 ;
			data[54319] <= 8'h10 ;
			data[54320] <= 8'h10 ;
			data[54321] <= 8'h10 ;
			data[54322] <= 8'h10 ;
			data[54323] <= 8'h10 ;
			data[54324] <= 8'h10 ;
			data[54325] <= 8'h10 ;
			data[54326] <= 8'h10 ;
			data[54327] <= 8'h10 ;
			data[54328] <= 8'h10 ;
			data[54329] <= 8'h10 ;
			data[54330] <= 8'h10 ;
			data[54331] <= 8'h10 ;
			data[54332] <= 8'h10 ;
			data[54333] <= 8'h10 ;
			data[54334] <= 8'h10 ;
			data[54335] <= 8'h10 ;
			data[54336] <= 8'h10 ;
			data[54337] <= 8'h10 ;
			data[54338] <= 8'h10 ;
			data[54339] <= 8'h10 ;
			data[54340] <= 8'h10 ;
			data[54341] <= 8'h10 ;
			data[54342] <= 8'h10 ;
			data[54343] <= 8'h10 ;
			data[54344] <= 8'h10 ;
			data[54345] <= 8'h10 ;
			data[54346] <= 8'h10 ;
			data[54347] <= 8'h10 ;
			data[54348] <= 8'h10 ;
			data[54349] <= 8'h10 ;
			data[54350] <= 8'h10 ;
			data[54351] <= 8'h10 ;
			data[54352] <= 8'h10 ;
			data[54353] <= 8'h10 ;
			data[54354] <= 8'h10 ;
			data[54355] <= 8'h10 ;
			data[54356] <= 8'h10 ;
			data[54357] <= 8'h10 ;
			data[54358] <= 8'h10 ;
			data[54359] <= 8'h10 ;
			data[54360] <= 8'h10 ;
			data[54361] <= 8'h10 ;
			data[54362] <= 8'h10 ;
			data[54363] <= 8'h10 ;
			data[54364] <= 8'h10 ;
			data[54365] <= 8'h10 ;
			data[54366] <= 8'h10 ;
			data[54367] <= 8'h10 ;
			data[54368] <= 8'h10 ;
			data[54369] <= 8'h10 ;
			data[54370] <= 8'h10 ;
			data[54371] <= 8'h10 ;
			data[54372] <= 8'h10 ;
			data[54373] <= 8'h10 ;
			data[54374] <= 8'h10 ;
			data[54375] <= 8'h10 ;
			data[54376] <= 8'h10 ;
			data[54377] <= 8'h10 ;
			data[54378] <= 8'h10 ;
			data[54379] <= 8'h10 ;
			data[54380] <= 8'h10 ;
			data[54381] <= 8'h10 ;
			data[54382] <= 8'h10 ;
			data[54383] <= 8'h10 ;
			data[54384] <= 8'h10 ;
			data[54385] <= 8'h10 ;
			data[54386] <= 8'h10 ;
			data[54387] <= 8'h10 ;
			data[54388] <= 8'h10 ;
			data[54389] <= 8'h10 ;
			data[54390] <= 8'h10 ;
			data[54391] <= 8'h10 ;
			data[54392] <= 8'h10 ;
			data[54393] <= 8'h10 ;
			data[54394] <= 8'h10 ;
			data[54395] <= 8'h10 ;
			data[54396] <= 8'h10 ;
			data[54397] <= 8'h10 ;
			data[54398] <= 8'h10 ;
			data[54399] <= 8'h10 ;
			data[54400] <= 8'h10 ;
			data[54401] <= 8'h10 ;
			data[54402] <= 8'h10 ;
			data[54403] <= 8'h10 ;
			data[54404] <= 8'h10 ;
			data[54405] <= 8'h10 ;
			data[54406] <= 8'h10 ;
			data[54407] <= 8'h10 ;
			data[54408] <= 8'h10 ;
			data[54409] <= 8'h10 ;
			data[54410] <= 8'h10 ;
			data[54411] <= 8'h10 ;
			data[54412] <= 8'h10 ;
			data[54413] <= 8'h10 ;
			data[54414] <= 8'h10 ;
			data[54415] <= 8'h10 ;
			data[54416] <= 8'h10 ;
			data[54417] <= 8'h10 ;
			data[54418] <= 8'h10 ;
			data[54419] <= 8'h10 ;
			data[54420] <= 8'h10 ;
			data[54421] <= 8'h10 ;
			data[54422] <= 8'h10 ;
			data[54423] <= 8'h10 ;
			data[54424] <= 8'h10 ;
			data[54425] <= 8'h10 ;
			data[54426] <= 8'h10 ;
			data[54427] <= 8'h10 ;
			data[54428] <= 8'h10 ;
			data[54429] <= 8'h10 ;
			data[54430] <= 8'h10 ;
			data[54431] <= 8'h10 ;
			data[54432] <= 8'h10 ;
			data[54433] <= 8'h10 ;
			data[54434] <= 8'h10 ;
			data[54435] <= 8'h10 ;
			data[54436] <= 8'h10 ;
			data[54437] <= 8'h10 ;
			data[54438] <= 8'h10 ;
			data[54439] <= 8'h10 ;
			data[54440] <= 8'h10 ;
			data[54441] <= 8'h10 ;
			data[54442] <= 8'h10 ;
			data[54443] <= 8'h10 ;
			data[54444] <= 8'h10 ;
			data[54445] <= 8'h10 ;
			data[54446] <= 8'h10 ;
			data[54447] <= 8'h10 ;
			data[54448] <= 8'h10 ;
			data[54449] <= 8'h10 ;
			data[54450] <= 8'h10 ;
			data[54451] <= 8'h10 ;
			data[54452] <= 8'h10 ;
			data[54453] <= 8'h10 ;
			data[54454] <= 8'h10 ;
			data[54455] <= 8'h10 ;
			data[54456] <= 8'h10 ;
			data[54457] <= 8'h10 ;
			data[54458] <= 8'h10 ;
			data[54459] <= 8'h10 ;
			data[54460] <= 8'h10 ;
			data[54461] <= 8'h10 ;
			data[54462] <= 8'h10 ;
			data[54463] <= 8'h10 ;
			data[54464] <= 8'h10 ;
			data[54465] <= 8'h10 ;
			data[54466] <= 8'h10 ;
			data[54467] <= 8'h10 ;
			data[54468] <= 8'h10 ;
			data[54469] <= 8'h10 ;
			data[54470] <= 8'h10 ;
			data[54471] <= 8'h10 ;
			data[54472] <= 8'h10 ;
			data[54473] <= 8'h10 ;
			data[54474] <= 8'h10 ;
			data[54475] <= 8'h10 ;
			data[54476] <= 8'h10 ;
			data[54477] <= 8'h10 ;
			data[54478] <= 8'h10 ;
			data[54479] <= 8'h10 ;
			data[54480] <= 8'h10 ;
			data[54481] <= 8'h10 ;
			data[54482] <= 8'h10 ;
			data[54483] <= 8'h10 ;
			data[54484] <= 8'h10 ;
			data[54485] <= 8'h10 ;
			data[54486] <= 8'h10 ;
			data[54487] <= 8'h10 ;
			data[54488] <= 8'h10 ;
			data[54489] <= 8'h10 ;
			data[54490] <= 8'h10 ;
			data[54491] <= 8'h10 ;
			data[54492] <= 8'h10 ;
			data[54493] <= 8'h10 ;
			data[54494] <= 8'h10 ;
			data[54495] <= 8'h10 ;
			data[54496] <= 8'h10 ;
			data[54497] <= 8'h10 ;
			data[54498] <= 8'h10 ;
			data[54499] <= 8'h10 ;
			data[54500] <= 8'h10 ;
			data[54501] <= 8'h10 ;
			data[54502] <= 8'h10 ;
			data[54503] <= 8'h10 ;
			data[54504] <= 8'h10 ;
			data[54505] <= 8'h10 ;
			data[54506] <= 8'h10 ;
			data[54507] <= 8'h10 ;
			data[54508] <= 8'h10 ;
			data[54509] <= 8'h10 ;
			data[54510] <= 8'h10 ;
			data[54511] <= 8'h10 ;
			data[54512] <= 8'h10 ;
			data[54513] <= 8'h10 ;
			data[54514] <= 8'h10 ;
			data[54515] <= 8'h10 ;
			data[54516] <= 8'h10 ;
			data[54517] <= 8'h10 ;
			data[54518] <= 8'h10 ;
			data[54519] <= 8'h10 ;
			data[54520] <= 8'h10 ;
			data[54521] <= 8'h10 ;
			data[54522] <= 8'h10 ;
			data[54523] <= 8'h10 ;
			data[54524] <= 8'h10 ;
			data[54525] <= 8'h10 ;
			data[54526] <= 8'h10 ;
			data[54527] <= 8'h10 ;
			data[54528] <= 8'h10 ;
			data[54529] <= 8'h10 ;
			data[54530] <= 8'h10 ;
			data[54531] <= 8'h10 ;
			data[54532] <= 8'h10 ;
			data[54533] <= 8'h10 ;
			data[54534] <= 8'h10 ;
			data[54535] <= 8'h10 ;
			data[54536] <= 8'h10 ;
			data[54537] <= 8'h10 ;
			data[54538] <= 8'h10 ;
			data[54539] <= 8'h10 ;
			data[54540] <= 8'h10 ;
			data[54541] <= 8'h10 ;
			data[54542] <= 8'h10 ;
			data[54543] <= 8'h10 ;
			data[54544] <= 8'h10 ;
			data[54545] <= 8'h10 ;
			data[54546] <= 8'h10 ;
			data[54547] <= 8'h10 ;
			data[54548] <= 8'h10 ;
			data[54549] <= 8'h10 ;
			data[54550] <= 8'h10 ;
			data[54551] <= 8'h10 ;
			data[54552] <= 8'h10 ;
			data[54553] <= 8'h10 ;
			data[54554] <= 8'h10 ;
			data[54555] <= 8'h10 ;
			data[54556] <= 8'h10 ;
			data[54557] <= 8'h10 ;
			data[54558] <= 8'h10 ;
			data[54559] <= 8'h10 ;
			data[54560] <= 8'h10 ;
			data[54561] <= 8'h10 ;
			data[54562] <= 8'h10 ;
			data[54563] <= 8'h10 ;
			data[54564] <= 8'h10 ;
			data[54565] <= 8'h10 ;
			data[54566] <= 8'h10 ;
			data[54567] <= 8'h10 ;
			data[54568] <= 8'h10 ;
			data[54569] <= 8'h10 ;
			data[54570] <= 8'h10 ;
			data[54571] <= 8'h10 ;
			data[54572] <= 8'h10 ;
			data[54573] <= 8'h10 ;
			data[54574] <= 8'h10 ;
			data[54575] <= 8'h10 ;
			data[54576] <= 8'h10 ;
			data[54577] <= 8'h10 ;
			data[54578] <= 8'h10 ;
			data[54579] <= 8'h10 ;
			data[54580] <= 8'h10 ;
			data[54581] <= 8'h10 ;
			data[54582] <= 8'h10 ;
			data[54583] <= 8'h10 ;
			data[54584] <= 8'h10 ;
			data[54585] <= 8'h10 ;
			data[54586] <= 8'h10 ;
			data[54587] <= 8'h10 ;
			data[54588] <= 8'h10 ;
			data[54589] <= 8'h10 ;
			data[54590] <= 8'h10 ;
			data[54591] <= 8'h10 ;
			data[54592] <= 8'h10 ;
			data[54593] <= 8'h10 ;
			data[54594] <= 8'h10 ;
			data[54595] <= 8'h10 ;
			data[54596] <= 8'h10 ;
			data[54597] <= 8'h10 ;
			data[54598] <= 8'h10 ;
			data[54599] <= 8'h10 ;
			data[54600] <= 8'h10 ;
			data[54601] <= 8'h10 ;
			data[54602] <= 8'h10 ;
			data[54603] <= 8'h10 ;
			data[54604] <= 8'h10 ;
			data[54605] <= 8'h10 ;
			data[54606] <= 8'h10 ;
			data[54607] <= 8'h10 ;
			data[54608] <= 8'h10 ;
			data[54609] <= 8'h10 ;
			data[54610] <= 8'h10 ;
			data[54611] <= 8'h10 ;
			data[54612] <= 8'h10 ;
			data[54613] <= 8'h10 ;
			data[54614] <= 8'h10 ;
			data[54615] <= 8'h10 ;
			data[54616] <= 8'h10 ;
			data[54617] <= 8'h10 ;
			data[54618] <= 8'h10 ;
			data[54619] <= 8'h10 ;
			data[54620] <= 8'h10 ;
			data[54621] <= 8'h10 ;
			data[54622] <= 8'h10 ;
			data[54623] <= 8'h10 ;
			data[54624] <= 8'h10 ;
			data[54625] <= 8'h10 ;
			data[54626] <= 8'h10 ;
			data[54627] <= 8'h10 ;
			data[54628] <= 8'h10 ;
			data[54629] <= 8'h10 ;
			data[54630] <= 8'h10 ;
			data[54631] <= 8'h10 ;
			data[54632] <= 8'h10 ;
			data[54633] <= 8'h10 ;
			data[54634] <= 8'h10 ;
			data[54635] <= 8'h10 ;
			data[54636] <= 8'h10 ;
			data[54637] <= 8'h10 ;
			data[54638] <= 8'h10 ;
			data[54639] <= 8'h10 ;
			data[54640] <= 8'h10 ;
			data[54641] <= 8'h10 ;
			data[54642] <= 8'h10 ;
			data[54643] <= 8'h10 ;
			data[54644] <= 8'h10 ;
			data[54645] <= 8'h10 ;
			data[54646] <= 8'h10 ;
			data[54647] <= 8'h10 ;
			data[54648] <= 8'h10 ;
			data[54649] <= 8'h10 ;
			data[54650] <= 8'h10 ;
			data[54651] <= 8'h10 ;
			data[54652] <= 8'h10 ;
			data[54653] <= 8'h10 ;
			data[54654] <= 8'h10 ;
			data[54655] <= 8'h10 ;
			data[54656] <= 8'h10 ;
			data[54657] <= 8'h10 ;
			data[54658] <= 8'h10 ;
			data[54659] <= 8'h10 ;
			data[54660] <= 8'h10 ;
			data[54661] <= 8'h10 ;
			data[54662] <= 8'h10 ;
			data[54663] <= 8'h10 ;
			data[54664] <= 8'h10 ;
			data[54665] <= 8'h10 ;
			data[54666] <= 8'h10 ;
			data[54667] <= 8'h10 ;
			data[54668] <= 8'h10 ;
			data[54669] <= 8'h10 ;
			data[54670] <= 8'h10 ;
			data[54671] <= 8'h10 ;
			data[54672] <= 8'h10 ;
			data[54673] <= 8'h10 ;
			data[54674] <= 8'h10 ;
			data[54675] <= 8'h10 ;
			data[54676] <= 8'h10 ;
			data[54677] <= 8'h10 ;
			data[54678] <= 8'h10 ;
			data[54679] <= 8'h10 ;
			data[54680] <= 8'h10 ;
			data[54681] <= 8'h10 ;
			data[54682] <= 8'h10 ;
			data[54683] <= 8'h10 ;
			data[54684] <= 8'h10 ;
			data[54685] <= 8'h10 ;
			data[54686] <= 8'h10 ;
			data[54687] <= 8'h10 ;
			data[54688] <= 8'h10 ;
			data[54689] <= 8'h10 ;
			data[54690] <= 8'h10 ;
			data[54691] <= 8'h10 ;
			data[54692] <= 8'h10 ;
			data[54693] <= 8'h10 ;
			data[54694] <= 8'h10 ;
			data[54695] <= 8'h10 ;
			data[54696] <= 8'h10 ;
			data[54697] <= 8'h10 ;
			data[54698] <= 8'h10 ;
			data[54699] <= 8'h10 ;
			data[54700] <= 8'h10 ;
			data[54701] <= 8'h10 ;
			data[54702] <= 8'h10 ;
			data[54703] <= 8'h10 ;
			data[54704] <= 8'h10 ;
			data[54705] <= 8'h10 ;
			data[54706] <= 8'h10 ;
			data[54707] <= 8'h10 ;
			data[54708] <= 8'h10 ;
			data[54709] <= 8'h10 ;
			data[54710] <= 8'h10 ;
			data[54711] <= 8'h10 ;
			data[54712] <= 8'h10 ;
			data[54713] <= 8'h10 ;
			data[54714] <= 8'h10 ;
			data[54715] <= 8'h10 ;
			data[54716] <= 8'h10 ;
			data[54717] <= 8'h10 ;
			data[54718] <= 8'h10 ;
			data[54719] <= 8'h10 ;
			data[54720] <= 8'h10 ;
			data[54721] <= 8'h10 ;
			data[54722] <= 8'h10 ;
			data[54723] <= 8'h10 ;
			data[54724] <= 8'h10 ;
			data[54725] <= 8'h10 ;
			data[54726] <= 8'h10 ;
			data[54727] <= 8'h10 ;
			data[54728] <= 8'h10 ;
			data[54729] <= 8'h10 ;
			data[54730] <= 8'h10 ;
			data[54731] <= 8'h10 ;
			data[54732] <= 8'h10 ;
			data[54733] <= 8'h10 ;
			data[54734] <= 8'h10 ;
			data[54735] <= 8'h10 ;
			data[54736] <= 8'h10 ;
			data[54737] <= 8'h10 ;
			data[54738] <= 8'h10 ;
			data[54739] <= 8'h10 ;
			data[54740] <= 8'h10 ;
			data[54741] <= 8'h10 ;
			data[54742] <= 8'h10 ;
			data[54743] <= 8'h10 ;
			data[54744] <= 8'h10 ;
			data[54745] <= 8'h10 ;
			data[54746] <= 8'h10 ;
			data[54747] <= 8'h10 ;
			data[54748] <= 8'h10 ;
			data[54749] <= 8'h10 ;
			data[54750] <= 8'h10 ;
			data[54751] <= 8'h10 ;
			data[54752] <= 8'h10 ;
			data[54753] <= 8'h10 ;
			data[54754] <= 8'h10 ;
			data[54755] <= 8'h10 ;
			data[54756] <= 8'h10 ;
			data[54757] <= 8'h10 ;
			data[54758] <= 8'h10 ;
			data[54759] <= 8'h10 ;
			data[54760] <= 8'h10 ;
			data[54761] <= 8'h10 ;
			data[54762] <= 8'h10 ;
			data[54763] <= 8'h10 ;
			data[54764] <= 8'h10 ;
			data[54765] <= 8'h10 ;
			data[54766] <= 8'h10 ;
			data[54767] <= 8'h10 ;
			data[54768] <= 8'h10 ;
			data[54769] <= 8'h10 ;
			data[54770] <= 8'h10 ;
			data[54771] <= 8'h10 ;
			data[54772] <= 8'h10 ;
			data[54773] <= 8'h10 ;
			data[54774] <= 8'h10 ;
			data[54775] <= 8'h10 ;
			data[54776] <= 8'h10 ;
			data[54777] <= 8'h10 ;
			data[54778] <= 8'h10 ;
			data[54779] <= 8'h10 ;
			data[54780] <= 8'h10 ;
			data[54781] <= 8'h10 ;
			data[54782] <= 8'h10 ;
			data[54783] <= 8'h10 ;
			data[54784] <= 8'h10 ;
			data[54785] <= 8'h10 ;
			data[54786] <= 8'h10 ;
			data[54787] <= 8'h10 ;
			data[54788] <= 8'h10 ;
			data[54789] <= 8'h10 ;
			data[54790] <= 8'h10 ;
			data[54791] <= 8'h10 ;
			data[54792] <= 8'h10 ;
			data[54793] <= 8'h10 ;
			data[54794] <= 8'h10 ;
			data[54795] <= 8'h10 ;
			data[54796] <= 8'h10 ;
			data[54797] <= 8'h10 ;
			data[54798] <= 8'h10 ;
			data[54799] <= 8'h10 ;
			data[54800] <= 8'h10 ;
			data[54801] <= 8'h10 ;
			data[54802] <= 8'h10 ;
			data[54803] <= 8'h10 ;
			data[54804] <= 8'h10 ;
			data[54805] <= 8'h10 ;
			data[54806] <= 8'h10 ;
			data[54807] <= 8'h10 ;
			data[54808] <= 8'h10 ;
			data[54809] <= 8'h10 ;
			data[54810] <= 8'h10 ;
			data[54811] <= 8'h10 ;
			data[54812] <= 8'h10 ;
			data[54813] <= 8'h10 ;
			data[54814] <= 8'h10 ;
			data[54815] <= 8'h10 ;
			data[54816] <= 8'h10 ;
			data[54817] <= 8'h10 ;
			data[54818] <= 8'h10 ;
			data[54819] <= 8'h10 ;
			data[54820] <= 8'h10 ;
			data[54821] <= 8'h10 ;
			data[54822] <= 8'h10 ;
			data[54823] <= 8'h10 ;
			data[54824] <= 8'h10 ;
			data[54825] <= 8'h10 ;
			data[54826] <= 8'h10 ;
			data[54827] <= 8'h10 ;
			data[54828] <= 8'h10 ;
			data[54829] <= 8'h10 ;
			data[54830] <= 8'h10 ;
			data[54831] <= 8'h10 ;
			data[54832] <= 8'h10 ;
			data[54833] <= 8'h10 ;
			data[54834] <= 8'h10 ;
			data[54835] <= 8'h10 ;
			data[54836] <= 8'h10 ;
			data[54837] <= 8'h10 ;
			data[54838] <= 8'h10 ;
			data[54839] <= 8'h10 ;
			data[54840] <= 8'h10 ;
			data[54841] <= 8'h10 ;
			data[54842] <= 8'h10 ;
			data[54843] <= 8'h10 ;
			data[54844] <= 8'h10 ;
			data[54845] <= 8'h10 ;
			data[54846] <= 8'h10 ;
			data[54847] <= 8'h10 ;
			data[54848] <= 8'h10 ;
			data[54849] <= 8'h10 ;
			data[54850] <= 8'h10 ;
			data[54851] <= 8'h10 ;
			data[54852] <= 8'h10 ;
			data[54853] <= 8'h10 ;
			data[54854] <= 8'h10 ;
			data[54855] <= 8'h10 ;
			data[54856] <= 8'h10 ;
			data[54857] <= 8'h10 ;
			data[54858] <= 8'h10 ;
			data[54859] <= 8'h10 ;
			data[54860] <= 8'h10 ;
			data[54861] <= 8'h10 ;
			data[54862] <= 8'h10 ;
			data[54863] <= 8'h10 ;
			data[54864] <= 8'h10 ;
			data[54865] <= 8'h10 ;
			data[54866] <= 8'h10 ;
			data[54867] <= 8'h10 ;
			data[54868] <= 8'h10 ;
			data[54869] <= 8'h10 ;
			data[54870] <= 8'h10 ;
			data[54871] <= 8'h10 ;
			data[54872] <= 8'h10 ;
			data[54873] <= 8'h10 ;
			data[54874] <= 8'h10 ;
			data[54875] <= 8'h10 ;
			data[54876] <= 8'h10 ;
			data[54877] <= 8'h10 ;
			data[54878] <= 8'h10 ;
			data[54879] <= 8'h10 ;
			data[54880] <= 8'h10 ;
			data[54881] <= 8'h10 ;
			data[54882] <= 8'h10 ;
			data[54883] <= 8'h10 ;
			data[54884] <= 8'h10 ;
			data[54885] <= 8'h10 ;
			data[54886] <= 8'h10 ;
			data[54887] <= 8'h10 ;
			data[54888] <= 8'h10 ;
			data[54889] <= 8'h10 ;
			data[54890] <= 8'h10 ;
			data[54891] <= 8'h10 ;
			data[54892] <= 8'h10 ;
			data[54893] <= 8'h10 ;
			data[54894] <= 8'h10 ;
			data[54895] <= 8'h10 ;
			data[54896] <= 8'h10 ;
			data[54897] <= 8'h10 ;
			data[54898] <= 8'h10 ;
			data[54899] <= 8'h10 ;
			data[54900] <= 8'h10 ;
			data[54901] <= 8'h10 ;
			data[54902] <= 8'h10 ;
			data[54903] <= 8'h10 ;
			data[54904] <= 8'h10 ;
			data[54905] <= 8'h10 ;
			data[54906] <= 8'h10 ;
			data[54907] <= 8'h10 ;
			data[54908] <= 8'h10 ;
			data[54909] <= 8'h10 ;
			data[54910] <= 8'h10 ;
			data[54911] <= 8'h10 ;
			data[54912] <= 8'h10 ;
			data[54913] <= 8'h10 ;
			data[54914] <= 8'h10 ;
			data[54915] <= 8'h10 ;
			data[54916] <= 8'h10 ;
			data[54917] <= 8'h10 ;
			data[54918] <= 8'h10 ;
			data[54919] <= 8'h10 ;
			data[54920] <= 8'h10 ;
			data[54921] <= 8'h10 ;
			data[54922] <= 8'h10 ;
			data[54923] <= 8'h10 ;
			data[54924] <= 8'h10 ;
			data[54925] <= 8'h10 ;
			data[54926] <= 8'h10 ;
			data[54927] <= 8'h10 ;
			data[54928] <= 8'h10 ;
			data[54929] <= 8'h10 ;
			data[54930] <= 8'h10 ;
			data[54931] <= 8'h10 ;
			data[54932] <= 8'h10 ;
			data[54933] <= 8'h10 ;
			data[54934] <= 8'h10 ;
			data[54935] <= 8'h10 ;
			data[54936] <= 8'h10 ;
			data[54937] <= 8'h10 ;
			data[54938] <= 8'h10 ;
			data[54939] <= 8'h10 ;
			data[54940] <= 8'h10 ;
			data[54941] <= 8'h10 ;
			data[54942] <= 8'h10 ;
			data[54943] <= 8'h10 ;
			data[54944] <= 8'h10 ;
			data[54945] <= 8'h10 ;
			data[54946] <= 8'h10 ;
			data[54947] <= 8'h10 ;
			data[54948] <= 8'h10 ;
			data[54949] <= 8'h10 ;
			data[54950] <= 8'h10 ;
			data[54951] <= 8'h10 ;
			data[54952] <= 8'h10 ;
			data[54953] <= 8'h10 ;
			data[54954] <= 8'h10 ;
			data[54955] <= 8'h10 ;
			data[54956] <= 8'h10 ;
			data[54957] <= 8'h10 ;
			data[54958] <= 8'h10 ;
			data[54959] <= 8'h10 ;
			data[54960] <= 8'h10 ;
			data[54961] <= 8'h10 ;
			data[54962] <= 8'h10 ;
			data[54963] <= 8'h10 ;
			data[54964] <= 8'h10 ;
			data[54965] <= 8'h10 ;
			data[54966] <= 8'h10 ;
			data[54967] <= 8'h10 ;
			data[54968] <= 8'h10 ;
			data[54969] <= 8'h10 ;
			data[54970] <= 8'h10 ;
			data[54971] <= 8'h10 ;
			data[54972] <= 8'h10 ;
			data[54973] <= 8'h10 ;
			data[54974] <= 8'h10 ;
			data[54975] <= 8'h10 ;
			data[54976] <= 8'h10 ;
			data[54977] <= 8'h10 ;
			data[54978] <= 8'h10 ;
			data[54979] <= 8'h10 ;
			data[54980] <= 8'h10 ;
			data[54981] <= 8'h10 ;
			data[54982] <= 8'h10 ;
			data[54983] <= 8'h10 ;
			data[54984] <= 8'h10 ;
			data[54985] <= 8'h10 ;
			data[54986] <= 8'h10 ;
			data[54987] <= 8'h10 ;
			data[54988] <= 8'h10 ;
			data[54989] <= 8'h10 ;
			data[54990] <= 8'h10 ;
			data[54991] <= 8'h10 ;
			data[54992] <= 8'h10 ;
			data[54993] <= 8'h10 ;
			data[54994] <= 8'h10 ;
			data[54995] <= 8'h10 ;
			data[54996] <= 8'h10 ;
			data[54997] <= 8'h10 ;
			data[54998] <= 8'h10 ;
			data[54999] <= 8'h10 ;
			data[55000] <= 8'h10 ;
			data[55001] <= 8'h10 ;
			data[55002] <= 8'h10 ;
			data[55003] <= 8'h10 ;
			data[55004] <= 8'h10 ;
			data[55005] <= 8'h10 ;
			data[55006] <= 8'h10 ;
			data[55007] <= 8'h10 ;
			data[55008] <= 8'h10 ;
			data[55009] <= 8'h10 ;
			data[55010] <= 8'h10 ;
			data[55011] <= 8'h10 ;
			data[55012] <= 8'h10 ;
			data[55013] <= 8'h10 ;
			data[55014] <= 8'h10 ;
			data[55015] <= 8'h10 ;
			data[55016] <= 8'h10 ;
			data[55017] <= 8'h10 ;
			data[55018] <= 8'h10 ;
			data[55019] <= 8'h10 ;
			data[55020] <= 8'h10 ;
			data[55021] <= 8'h10 ;
			data[55022] <= 8'h10 ;
			data[55023] <= 8'h10 ;
			data[55024] <= 8'h10 ;
			data[55025] <= 8'h10 ;
			data[55026] <= 8'h10 ;
			data[55027] <= 8'h10 ;
			data[55028] <= 8'h10 ;
			data[55029] <= 8'h10 ;
			data[55030] <= 8'h10 ;
			data[55031] <= 8'h10 ;
			data[55032] <= 8'h10 ;
			data[55033] <= 8'h10 ;
			data[55034] <= 8'h10 ;
			data[55035] <= 8'h10 ;
			data[55036] <= 8'h10 ;
			data[55037] <= 8'h10 ;
			data[55038] <= 8'h10 ;
			data[55039] <= 8'h10 ;
			data[55040] <= 8'h10 ;
			data[55041] <= 8'h10 ;
			data[55042] <= 8'h10 ;
			data[55043] <= 8'h10 ;
			data[55044] <= 8'h10 ;
			data[55045] <= 8'h10 ;
			data[55046] <= 8'h10 ;
			data[55047] <= 8'h10 ;
			data[55048] <= 8'h10 ;
			data[55049] <= 8'h10 ;
			data[55050] <= 8'h10 ;
			data[55051] <= 8'h10 ;
			data[55052] <= 8'h10 ;
			data[55053] <= 8'h10 ;
			data[55054] <= 8'h10 ;
			data[55055] <= 8'h10 ;
			data[55056] <= 8'h10 ;
			data[55057] <= 8'h10 ;
			data[55058] <= 8'h10 ;
			data[55059] <= 8'h10 ;
			data[55060] <= 8'h10 ;
			data[55061] <= 8'h10 ;
			data[55062] <= 8'h10 ;
			data[55063] <= 8'h10 ;
			data[55064] <= 8'h10 ;
			data[55065] <= 8'h10 ;
			data[55066] <= 8'h10 ;
			data[55067] <= 8'h10 ;
			data[55068] <= 8'h10 ;
			data[55069] <= 8'h10 ;
			data[55070] <= 8'h10 ;
			data[55071] <= 8'h10 ;
			data[55072] <= 8'h10 ;
			data[55073] <= 8'h10 ;
			data[55074] <= 8'h10 ;
			data[55075] <= 8'h10 ;
			data[55076] <= 8'h10 ;
			data[55077] <= 8'h10 ;
			data[55078] <= 8'h10 ;
			data[55079] <= 8'h10 ;
			data[55080] <= 8'h10 ;
			data[55081] <= 8'h10 ;
			data[55082] <= 8'h10 ;
			data[55083] <= 8'h10 ;
			data[55084] <= 8'h10 ;
			data[55085] <= 8'h10 ;
			data[55086] <= 8'h10 ;
			data[55087] <= 8'h10 ;
			data[55088] <= 8'h10 ;
			data[55089] <= 8'h10 ;
			data[55090] <= 8'h10 ;
			data[55091] <= 8'h10 ;
			data[55092] <= 8'h10 ;
			data[55093] <= 8'h10 ;
			data[55094] <= 8'h10 ;
			data[55095] <= 8'h10 ;
			data[55096] <= 8'h10 ;
			data[55097] <= 8'h10 ;
			data[55098] <= 8'h10 ;
			data[55099] <= 8'h10 ;
			data[55100] <= 8'h10 ;
			data[55101] <= 8'h10 ;
			data[55102] <= 8'h10 ;
			data[55103] <= 8'h10 ;
			data[55104] <= 8'h10 ;
			data[55105] <= 8'h10 ;
			data[55106] <= 8'h10 ;
			data[55107] <= 8'h10 ;
			data[55108] <= 8'h10 ;
			data[55109] <= 8'h10 ;
			data[55110] <= 8'h10 ;
			data[55111] <= 8'h10 ;
			data[55112] <= 8'h10 ;
			data[55113] <= 8'h10 ;
			data[55114] <= 8'h10 ;
			data[55115] <= 8'h10 ;
			data[55116] <= 8'h10 ;
			data[55117] <= 8'h10 ;
			data[55118] <= 8'h10 ;
			data[55119] <= 8'h10 ;
			data[55120] <= 8'h10 ;
			data[55121] <= 8'h10 ;
			data[55122] <= 8'h10 ;
			data[55123] <= 8'h10 ;
			data[55124] <= 8'h10 ;
			data[55125] <= 8'h10 ;
			data[55126] <= 8'h10 ;
			data[55127] <= 8'h10 ;
			data[55128] <= 8'h10 ;
			data[55129] <= 8'h10 ;
			data[55130] <= 8'h10 ;
			data[55131] <= 8'h10 ;
			data[55132] <= 8'h10 ;
			data[55133] <= 8'h10 ;
			data[55134] <= 8'h10 ;
			data[55135] <= 8'h10 ;
			data[55136] <= 8'h10 ;
			data[55137] <= 8'h10 ;
			data[55138] <= 8'h10 ;
			data[55139] <= 8'h10 ;
			data[55140] <= 8'h10 ;
			data[55141] <= 8'h10 ;
			data[55142] <= 8'h10 ;
			data[55143] <= 8'h10 ;
			data[55144] <= 8'h10 ;
			data[55145] <= 8'h10 ;
			data[55146] <= 8'h10 ;
			data[55147] <= 8'h10 ;
			data[55148] <= 8'h10 ;
			data[55149] <= 8'h10 ;
			data[55150] <= 8'h10 ;
			data[55151] <= 8'h10 ;
			data[55152] <= 8'h10 ;
			data[55153] <= 8'h10 ;
			data[55154] <= 8'h10 ;
			data[55155] <= 8'h10 ;
			data[55156] <= 8'h10 ;
			data[55157] <= 8'h10 ;
			data[55158] <= 8'h10 ;
			data[55159] <= 8'h10 ;
			data[55160] <= 8'h10 ;
			data[55161] <= 8'h10 ;
			data[55162] <= 8'h10 ;
			data[55163] <= 8'h10 ;
			data[55164] <= 8'h10 ;
			data[55165] <= 8'h10 ;
			data[55166] <= 8'h10 ;
			data[55167] <= 8'h10 ;
			data[55168] <= 8'h10 ;
			data[55169] <= 8'h10 ;
			data[55170] <= 8'h10 ;
			data[55171] <= 8'h10 ;
			data[55172] <= 8'h10 ;
			data[55173] <= 8'h10 ;
			data[55174] <= 8'h10 ;
			data[55175] <= 8'h10 ;
			data[55176] <= 8'h10 ;
			data[55177] <= 8'h10 ;
			data[55178] <= 8'h10 ;
			data[55179] <= 8'h10 ;
			data[55180] <= 8'h10 ;
			data[55181] <= 8'h10 ;
			data[55182] <= 8'h10 ;
			data[55183] <= 8'h10 ;
			data[55184] <= 8'h10 ;
			data[55185] <= 8'h10 ;
			data[55186] <= 8'h10 ;
			data[55187] <= 8'h10 ;
			data[55188] <= 8'h10 ;
			data[55189] <= 8'h10 ;
			data[55190] <= 8'h10 ;
			data[55191] <= 8'h10 ;
			data[55192] <= 8'h10 ;
			data[55193] <= 8'h10 ;
			data[55194] <= 8'h10 ;
			data[55195] <= 8'h10 ;
			data[55196] <= 8'h10 ;
			data[55197] <= 8'h10 ;
			data[55198] <= 8'h10 ;
			data[55199] <= 8'h10 ;
			data[55200] <= 8'h10 ;
			data[55201] <= 8'h10 ;
			data[55202] <= 8'h10 ;
			data[55203] <= 8'h10 ;
			data[55204] <= 8'h10 ;
			data[55205] <= 8'h10 ;
			data[55206] <= 8'h10 ;
			data[55207] <= 8'h10 ;
			data[55208] <= 8'h10 ;
			data[55209] <= 8'h10 ;
			data[55210] <= 8'h10 ;
			data[55211] <= 8'h10 ;
			data[55212] <= 8'h10 ;
			data[55213] <= 8'h10 ;
			data[55214] <= 8'h10 ;
			data[55215] <= 8'h10 ;
			data[55216] <= 8'h10 ;
			data[55217] <= 8'h10 ;
			data[55218] <= 8'h10 ;
			data[55219] <= 8'h10 ;
			data[55220] <= 8'h10 ;
			data[55221] <= 8'h10 ;
			data[55222] <= 8'h10 ;
			data[55223] <= 8'h10 ;
			data[55224] <= 8'h10 ;
			data[55225] <= 8'h10 ;
			data[55226] <= 8'h10 ;
			data[55227] <= 8'h10 ;
			data[55228] <= 8'h10 ;
			data[55229] <= 8'h10 ;
			data[55230] <= 8'h10 ;
			data[55231] <= 8'h10 ;
			data[55232] <= 8'h10 ;
			data[55233] <= 8'h10 ;
			data[55234] <= 8'h10 ;
			data[55235] <= 8'h10 ;
			data[55236] <= 8'h10 ;
			data[55237] <= 8'h10 ;
			data[55238] <= 8'h10 ;
			data[55239] <= 8'h10 ;
			data[55240] <= 8'h10 ;
			data[55241] <= 8'h10 ;
			data[55242] <= 8'h10 ;
			data[55243] <= 8'h10 ;
			data[55244] <= 8'h10 ;
			data[55245] <= 8'h10 ;
			data[55246] <= 8'h10 ;
			data[55247] <= 8'h10 ;
			data[55248] <= 8'h10 ;
			data[55249] <= 8'h10 ;
			data[55250] <= 8'h10 ;
			data[55251] <= 8'h10 ;
			data[55252] <= 8'h10 ;
			data[55253] <= 8'h10 ;
			data[55254] <= 8'h10 ;
			data[55255] <= 8'h10 ;
			data[55256] <= 8'h10 ;
			data[55257] <= 8'h10 ;
			data[55258] <= 8'h10 ;
			data[55259] <= 8'h10 ;
			data[55260] <= 8'h10 ;
			data[55261] <= 8'h10 ;
			data[55262] <= 8'h10 ;
			data[55263] <= 8'h10 ;
			data[55264] <= 8'h10 ;
			data[55265] <= 8'h10 ;
			data[55266] <= 8'h10 ;
			data[55267] <= 8'h10 ;
			data[55268] <= 8'h10 ;
			data[55269] <= 8'h10 ;
			data[55270] <= 8'h10 ;
			data[55271] <= 8'h10 ;
			data[55272] <= 8'h10 ;
			data[55273] <= 8'h10 ;
			data[55274] <= 8'h10 ;
			data[55275] <= 8'h10 ;
			data[55276] <= 8'h10 ;
			data[55277] <= 8'h10 ;
			data[55278] <= 8'h10 ;
			data[55279] <= 8'h10 ;
			data[55280] <= 8'h10 ;
			data[55281] <= 8'h10 ;
			data[55282] <= 8'h10 ;
			data[55283] <= 8'h10 ;
			data[55284] <= 8'h10 ;
			data[55285] <= 8'h10 ;
			data[55286] <= 8'h10 ;
			data[55287] <= 8'h10 ;
			data[55288] <= 8'h10 ;
			data[55289] <= 8'h10 ;
			data[55290] <= 8'h10 ;
			data[55291] <= 8'h10 ;
			data[55292] <= 8'h10 ;
			data[55293] <= 8'h10 ;
			data[55294] <= 8'h10 ;
			data[55295] <= 8'h10 ;
			data[55296] <= 8'h10 ;
			data[55297] <= 8'h10 ;
			data[55298] <= 8'h10 ;
			data[55299] <= 8'h10 ;
			data[55300] <= 8'h10 ;
			data[55301] <= 8'h10 ;
			data[55302] <= 8'h10 ;
			data[55303] <= 8'h10 ;
			data[55304] <= 8'h10 ;
			data[55305] <= 8'h10 ;
			data[55306] <= 8'h10 ;
			data[55307] <= 8'h10 ;
			data[55308] <= 8'h10 ;
			data[55309] <= 8'h10 ;
			data[55310] <= 8'h10 ;
			data[55311] <= 8'h10 ;
			data[55312] <= 8'h10 ;
			data[55313] <= 8'h10 ;
			data[55314] <= 8'h10 ;
			data[55315] <= 8'h10 ;
			data[55316] <= 8'h10 ;
			data[55317] <= 8'h10 ;
			data[55318] <= 8'h10 ;
			data[55319] <= 8'h10 ;
			data[55320] <= 8'h10 ;
			data[55321] <= 8'h10 ;
			data[55322] <= 8'h10 ;
			data[55323] <= 8'h10 ;
			data[55324] <= 8'h10 ;
			data[55325] <= 8'h10 ;
			data[55326] <= 8'h10 ;
			data[55327] <= 8'h10 ;
			data[55328] <= 8'h10 ;
			data[55329] <= 8'h10 ;
			data[55330] <= 8'h10 ;
			data[55331] <= 8'h10 ;
			data[55332] <= 8'h10 ;
			data[55333] <= 8'h10 ;
			data[55334] <= 8'h10 ;
			data[55335] <= 8'h10 ;
			data[55336] <= 8'h10 ;
			data[55337] <= 8'h10 ;
			data[55338] <= 8'h10 ;
			data[55339] <= 8'h10 ;
			data[55340] <= 8'h10 ;
			data[55341] <= 8'h10 ;
			data[55342] <= 8'h10 ;
			data[55343] <= 8'h10 ;
			data[55344] <= 8'h10 ;
			data[55345] <= 8'h10 ;
			data[55346] <= 8'h10 ;
			data[55347] <= 8'h10 ;
			data[55348] <= 8'h10 ;
			data[55349] <= 8'h10 ;
			data[55350] <= 8'h10 ;
			data[55351] <= 8'h10 ;
			data[55352] <= 8'h10 ;
			data[55353] <= 8'h10 ;
			data[55354] <= 8'h10 ;
			data[55355] <= 8'h10 ;
			data[55356] <= 8'h10 ;
			data[55357] <= 8'h10 ;
			data[55358] <= 8'h10 ;
			data[55359] <= 8'h10 ;
			data[55360] <= 8'h10 ;
			data[55361] <= 8'h10 ;
			data[55362] <= 8'h10 ;
			data[55363] <= 8'h10 ;
			data[55364] <= 8'h10 ;
			data[55365] <= 8'h10 ;
			data[55366] <= 8'h10 ;
			data[55367] <= 8'h10 ;
			data[55368] <= 8'h10 ;
			data[55369] <= 8'h10 ;
			data[55370] <= 8'h10 ;
			data[55371] <= 8'h10 ;
			data[55372] <= 8'h10 ;
			data[55373] <= 8'h10 ;
			data[55374] <= 8'h10 ;
			data[55375] <= 8'h10 ;
			data[55376] <= 8'h10 ;
			data[55377] <= 8'h10 ;
			data[55378] <= 8'h10 ;
			data[55379] <= 8'h10 ;
			data[55380] <= 8'h10 ;
			data[55381] <= 8'h10 ;
			data[55382] <= 8'h10 ;
			data[55383] <= 8'h10 ;
			data[55384] <= 8'h10 ;
			data[55385] <= 8'h10 ;
			data[55386] <= 8'h10 ;
			data[55387] <= 8'h10 ;
			data[55388] <= 8'h10 ;
			data[55389] <= 8'h10 ;
			data[55390] <= 8'h10 ;
			data[55391] <= 8'h10 ;
			data[55392] <= 8'h10 ;
			data[55393] <= 8'h10 ;
			data[55394] <= 8'h10 ;
			data[55395] <= 8'h10 ;
			data[55396] <= 8'h10 ;
			data[55397] <= 8'h10 ;
			data[55398] <= 8'h10 ;
			data[55399] <= 8'h10 ;
			data[55400] <= 8'h10 ;
			data[55401] <= 8'h10 ;
			data[55402] <= 8'h10 ;
			data[55403] <= 8'h10 ;
			data[55404] <= 8'h10 ;
			data[55405] <= 8'h10 ;
			data[55406] <= 8'h10 ;
			data[55407] <= 8'h10 ;
			data[55408] <= 8'h10 ;
			data[55409] <= 8'h10 ;
			data[55410] <= 8'h10 ;
			data[55411] <= 8'h10 ;
			data[55412] <= 8'h10 ;
			data[55413] <= 8'h10 ;
			data[55414] <= 8'h10 ;
			data[55415] <= 8'h10 ;
			data[55416] <= 8'h10 ;
			data[55417] <= 8'h10 ;
			data[55418] <= 8'h10 ;
			data[55419] <= 8'h10 ;
			data[55420] <= 8'h10 ;
			data[55421] <= 8'h10 ;
			data[55422] <= 8'h10 ;
			data[55423] <= 8'h10 ;
			data[55424] <= 8'h10 ;
			data[55425] <= 8'h10 ;
			data[55426] <= 8'h10 ;
			data[55427] <= 8'h10 ;
			data[55428] <= 8'h10 ;
			data[55429] <= 8'h10 ;
			data[55430] <= 8'h10 ;
			data[55431] <= 8'h10 ;
			data[55432] <= 8'h10 ;
			data[55433] <= 8'h10 ;
			data[55434] <= 8'h10 ;
			data[55435] <= 8'h10 ;
			data[55436] <= 8'h10 ;
			data[55437] <= 8'h10 ;
			data[55438] <= 8'h10 ;
			data[55439] <= 8'h10 ;
			data[55440] <= 8'h10 ;
			data[55441] <= 8'h10 ;
			data[55442] <= 8'h10 ;
			data[55443] <= 8'h10 ;
			data[55444] <= 8'h10 ;
			data[55445] <= 8'h10 ;
			data[55446] <= 8'h10 ;
			data[55447] <= 8'h10 ;
			data[55448] <= 8'h10 ;
			data[55449] <= 8'h10 ;
			data[55450] <= 8'h10 ;
			data[55451] <= 8'h10 ;
			data[55452] <= 8'h10 ;
			data[55453] <= 8'h10 ;
			data[55454] <= 8'h10 ;
			data[55455] <= 8'h10 ;
			data[55456] <= 8'h10 ;
			data[55457] <= 8'h10 ;
			data[55458] <= 8'h10 ;
			data[55459] <= 8'h10 ;
			data[55460] <= 8'h10 ;
			data[55461] <= 8'h10 ;
			data[55462] <= 8'h10 ;
			data[55463] <= 8'h10 ;
			data[55464] <= 8'h10 ;
			data[55465] <= 8'h10 ;
			data[55466] <= 8'h10 ;
			data[55467] <= 8'h10 ;
			data[55468] <= 8'h10 ;
			data[55469] <= 8'h10 ;
			data[55470] <= 8'h10 ;
			data[55471] <= 8'h10 ;
			data[55472] <= 8'h10 ;
			data[55473] <= 8'h10 ;
			data[55474] <= 8'h10 ;
			data[55475] <= 8'h10 ;
			data[55476] <= 8'h10 ;
			data[55477] <= 8'h10 ;
			data[55478] <= 8'h10 ;
			data[55479] <= 8'h10 ;
			data[55480] <= 8'h10 ;
			data[55481] <= 8'h10 ;
			data[55482] <= 8'h10 ;
			data[55483] <= 8'h10 ;
			data[55484] <= 8'h10 ;
			data[55485] <= 8'h10 ;
			data[55486] <= 8'h10 ;
			data[55487] <= 8'h10 ;
			data[55488] <= 8'h10 ;
			data[55489] <= 8'h10 ;
			data[55490] <= 8'h10 ;
			data[55491] <= 8'h10 ;
			data[55492] <= 8'h10 ;
			data[55493] <= 8'h10 ;
			data[55494] <= 8'h10 ;
			data[55495] <= 8'h10 ;
			data[55496] <= 8'h10 ;
			data[55497] <= 8'h10 ;
			data[55498] <= 8'h10 ;
			data[55499] <= 8'h10 ;
			data[55500] <= 8'h10 ;
			data[55501] <= 8'h10 ;
			data[55502] <= 8'h10 ;
			data[55503] <= 8'h10 ;
			data[55504] <= 8'h10 ;
			data[55505] <= 8'h10 ;
			data[55506] <= 8'h10 ;
			data[55507] <= 8'h10 ;
			data[55508] <= 8'h10 ;
			data[55509] <= 8'h10 ;
			data[55510] <= 8'h10 ;
			data[55511] <= 8'h10 ;
			data[55512] <= 8'h10 ;
			data[55513] <= 8'h10 ;
			data[55514] <= 8'h10 ;
			data[55515] <= 8'h10 ;
			data[55516] <= 8'h10 ;
			data[55517] <= 8'h10 ;
			data[55518] <= 8'h10 ;
			data[55519] <= 8'h10 ;
			data[55520] <= 8'h10 ;
			data[55521] <= 8'h10 ;
			data[55522] <= 8'h10 ;
			data[55523] <= 8'h10 ;
			data[55524] <= 8'h10 ;
			data[55525] <= 8'h10 ;
			data[55526] <= 8'h10 ;
			data[55527] <= 8'h10 ;
			data[55528] <= 8'h10 ;
			data[55529] <= 8'h10 ;
			data[55530] <= 8'h10 ;
			data[55531] <= 8'h10 ;
			data[55532] <= 8'h10 ;
			data[55533] <= 8'h10 ;
			data[55534] <= 8'h10 ;
			data[55535] <= 8'h10 ;
			data[55536] <= 8'h10 ;
			data[55537] <= 8'h10 ;
			data[55538] <= 8'h10 ;
			data[55539] <= 8'h10 ;
			data[55540] <= 8'h10 ;
			data[55541] <= 8'h10 ;
			data[55542] <= 8'h10 ;
			data[55543] <= 8'h10 ;
			data[55544] <= 8'h10 ;
			data[55545] <= 8'h10 ;
			data[55546] <= 8'h10 ;
			data[55547] <= 8'h10 ;
			data[55548] <= 8'h10 ;
			data[55549] <= 8'h10 ;
			data[55550] <= 8'h10 ;
			data[55551] <= 8'h10 ;
			data[55552] <= 8'h10 ;
			data[55553] <= 8'h10 ;
			data[55554] <= 8'h10 ;
			data[55555] <= 8'h10 ;
			data[55556] <= 8'h10 ;
			data[55557] <= 8'h10 ;
			data[55558] <= 8'h10 ;
			data[55559] <= 8'h10 ;
			data[55560] <= 8'h10 ;
			data[55561] <= 8'h10 ;
			data[55562] <= 8'h10 ;
			data[55563] <= 8'h10 ;
			data[55564] <= 8'h10 ;
			data[55565] <= 8'h10 ;
			data[55566] <= 8'h10 ;
			data[55567] <= 8'h10 ;
			data[55568] <= 8'h10 ;
			data[55569] <= 8'h10 ;
			data[55570] <= 8'h10 ;
			data[55571] <= 8'h10 ;
			data[55572] <= 8'h10 ;
			data[55573] <= 8'h10 ;
			data[55574] <= 8'h10 ;
			data[55575] <= 8'h10 ;
			data[55576] <= 8'h10 ;
			data[55577] <= 8'h10 ;
			data[55578] <= 8'h10 ;
			data[55579] <= 8'h10 ;
			data[55580] <= 8'h10 ;
			data[55581] <= 8'h10 ;
			data[55582] <= 8'h10 ;
			data[55583] <= 8'h10 ;
			data[55584] <= 8'h10 ;
			data[55585] <= 8'h10 ;
			data[55586] <= 8'h10 ;
			data[55587] <= 8'h10 ;
			data[55588] <= 8'h10 ;
			data[55589] <= 8'h10 ;
			data[55590] <= 8'h10 ;
			data[55591] <= 8'h10 ;
			data[55592] <= 8'h10 ;
			data[55593] <= 8'h10 ;
			data[55594] <= 8'h10 ;
			data[55595] <= 8'h10 ;
			data[55596] <= 8'h10 ;
			data[55597] <= 8'h10 ;
			data[55598] <= 8'h10 ;
			data[55599] <= 8'h10 ;
			data[55600] <= 8'h10 ;
			data[55601] <= 8'h10 ;
			data[55602] <= 8'h10 ;
			data[55603] <= 8'h10 ;
			data[55604] <= 8'h10 ;
			data[55605] <= 8'h10 ;
			data[55606] <= 8'h10 ;
			data[55607] <= 8'h10 ;
			data[55608] <= 8'h10 ;
			data[55609] <= 8'h10 ;
			data[55610] <= 8'h10 ;
			data[55611] <= 8'h10 ;
			data[55612] <= 8'h10 ;
			data[55613] <= 8'h10 ;
			data[55614] <= 8'h10 ;
			data[55615] <= 8'h10 ;
			data[55616] <= 8'h10 ;
			data[55617] <= 8'h10 ;
			data[55618] <= 8'h10 ;
			data[55619] <= 8'h10 ;
			data[55620] <= 8'h10 ;
			data[55621] <= 8'h10 ;
			data[55622] <= 8'h10 ;
			data[55623] <= 8'h10 ;
			data[55624] <= 8'h10 ;
			data[55625] <= 8'h10 ;
			data[55626] <= 8'h10 ;
			data[55627] <= 8'h10 ;
			data[55628] <= 8'h10 ;
			data[55629] <= 8'h10 ;
			data[55630] <= 8'h10 ;
			data[55631] <= 8'h10 ;
			data[55632] <= 8'h10 ;
			data[55633] <= 8'h10 ;
			data[55634] <= 8'h10 ;
			data[55635] <= 8'h10 ;
			data[55636] <= 8'h10 ;
			data[55637] <= 8'h10 ;
			data[55638] <= 8'h10 ;
			data[55639] <= 8'h10 ;
			data[55640] <= 8'h10 ;
			data[55641] <= 8'h10 ;
			data[55642] <= 8'h10 ;
			data[55643] <= 8'h10 ;
			data[55644] <= 8'h10 ;
			data[55645] <= 8'h10 ;
			data[55646] <= 8'h10 ;
			data[55647] <= 8'h10 ;
			data[55648] <= 8'h10 ;
			data[55649] <= 8'h10 ;
			data[55650] <= 8'h10 ;
			data[55651] <= 8'h10 ;
			data[55652] <= 8'h10 ;
			data[55653] <= 8'h10 ;
			data[55654] <= 8'h10 ;
			data[55655] <= 8'h10 ;
			data[55656] <= 8'h10 ;
			data[55657] <= 8'h10 ;
			data[55658] <= 8'h10 ;
			data[55659] <= 8'h10 ;
			data[55660] <= 8'h10 ;
			data[55661] <= 8'h10 ;
			data[55662] <= 8'h10 ;
			data[55663] <= 8'h10 ;
			data[55664] <= 8'h10 ;
			data[55665] <= 8'h10 ;
			data[55666] <= 8'h10 ;
			data[55667] <= 8'h10 ;
			data[55668] <= 8'h10 ;
			data[55669] <= 8'h10 ;
			data[55670] <= 8'h10 ;
			data[55671] <= 8'h10 ;
			data[55672] <= 8'h10 ;
			data[55673] <= 8'h10 ;
			data[55674] <= 8'h10 ;
			data[55675] <= 8'h10 ;
			data[55676] <= 8'h10 ;
			data[55677] <= 8'h10 ;
			data[55678] <= 8'h10 ;
			data[55679] <= 8'h10 ;
			data[55680] <= 8'h10 ;
			data[55681] <= 8'h10 ;
			data[55682] <= 8'h10 ;
			data[55683] <= 8'h10 ;
			data[55684] <= 8'h10 ;
			data[55685] <= 8'h10 ;
			data[55686] <= 8'h10 ;
			data[55687] <= 8'h10 ;
			data[55688] <= 8'h10 ;
			data[55689] <= 8'h10 ;
			data[55690] <= 8'h10 ;
			data[55691] <= 8'h10 ;
			data[55692] <= 8'h10 ;
			data[55693] <= 8'h10 ;
			data[55694] <= 8'h10 ;
			data[55695] <= 8'h10 ;
			data[55696] <= 8'h10 ;
			data[55697] <= 8'h10 ;
			data[55698] <= 8'h10 ;
			data[55699] <= 8'h10 ;
			data[55700] <= 8'h10 ;
			data[55701] <= 8'h10 ;
			data[55702] <= 8'h10 ;
			data[55703] <= 8'h10 ;
			data[55704] <= 8'h10 ;
			data[55705] <= 8'h10 ;
			data[55706] <= 8'h10 ;
			data[55707] <= 8'h10 ;
			data[55708] <= 8'h10 ;
			data[55709] <= 8'h10 ;
			data[55710] <= 8'h10 ;
			data[55711] <= 8'h10 ;
			data[55712] <= 8'h10 ;
			data[55713] <= 8'h10 ;
			data[55714] <= 8'h10 ;
			data[55715] <= 8'h10 ;
			data[55716] <= 8'h10 ;
			data[55717] <= 8'h10 ;
			data[55718] <= 8'h10 ;
			data[55719] <= 8'h10 ;
			data[55720] <= 8'h10 ;
			data[55721] <= 8'h10 ;
			data[55722] <= 8'h10 ;
			data[55723] <= 8'h10 ;
			data[55724] <= 8'h10 ;
			data[55725] <= 8'h10 ;
			data[55726] <= 8'h10 ;
			data[55727] <= 8'h10 ;
			data[55728] <= 8'h10 ;
			data[55729] <= 8'h10 ;
			data[55730] <= 8'h10 ;
			data[55731] <= 8'h10 ;
			data[55732] <= 8'h10 ;
			data[55733] <= 8'h10 ;
			data[55734] <= 8'h10 ;
			data[55735] <= 8'h10 ;
			data[55736] <= 8'h10 ;
			data[55737] <= 8'h10 ;
			data[55738] <= 8'h10 ;
			data[55739] <= 8'h10 ;
			data[55740] <= 8'h10 ;
			data[55741] <= 8'h10 ;
			data[55742] <= 8'h10 ;
			data[55743] <= 8'h10 ;
			data[55744] <= 8'h10 ;
			data[55745] <= 8'h10 ;
			data[55746] <= 8'h10 ;
			data[55747] <= 8'h10 ;
			data[55748] <= 8'h10 ;
			data[55749] <= 8'h10 ;
			data[55750] <= 8'h10 ;
			data[55751] <= 8'h10 ;
			data[55752] <= 8'h10 ;
			data[55753] <= 8'h10 ;
			data[55754] <= 8'h10 ;
			data[55755] <= 8'h10 ;
			data[55756] <= 8'h10 ;
			data[55757] <= 8'h10 ;
			data[55758] <= 8'h10 ;
			data[55759] <= 8'h10 ;
			data[55760] <= 8'h10 ;
			data[55761] <= 8'h10 ;
			data[55762] <= 8'h10 ;
			data[55763] <= 8'h10 ;
			data[55764] <= 8'h10 ;
			data[55765] <= 8'h10 ;
			data[55766] <= 8'h10 ;
			data[55767] <= 8'h10 ;
			data[55768] <= 8'h10 ;
			data[55769] <= 8'h10 ;
			data[55770] <= 8'h10 ;
			data[55771] <= 8'h10 ;
			data[55772] <= 8'h10 ;
			data[55773] <= 8'h10 ;
			data[55774] <= 8'h10 ;
			data[55775] <= 8'h10 ;
			data[55776] <= 8'h10 ;
			data[55777] <= 8'h10 ;
			data[55778] <= 8'h10 ;
			data[55779] <= 8'h10 ;
			data[55780] <= 8'h10 ;
			data[55781] <= 8'h10 ;
			data[55782] <= 8'h10 ;
			data[55783] <= 8'h10 ;
			data[55784] <= 8'h10 ;
			data[55785] <= 8'h10 ;
			data[55786] <= 8'h10 ;
			data[55787] <= 8'h10 ;
			data[55788] <= 8'h10 ;
			data[55789] <= 8'h10 ;
			data[55790] <= 8'h10 ;
			data[55791] <= 8'h10 ;
			data[55792] <= 8'h10 ;
			data[55793] <= 8'h10 ;
			data[55794] <= 8'h10 ;
			data[55795] <= 8'h10 ;
			data[55796] <= 8'h10 ;
			data[55797] <= 8'h10 ;
			data[55798] <= 8'h10 ;
			data[55799] <= 8'h10 ;
			data[55800] <= 8'h10 ;
			data[55801] <= 8'h10 ;
			data[55802] <= 8'h10 ;
			data[55803] <= 8'h10 ;
			data[55804] <= 8'h10 ;
			data[55805] <= 8'h10 ;
			data[55806] <= 8'h10 ;
			data[55807] <= 8'h10 ;
			data[55808] <= 8'h10 ;
			data[55809] <= 8'h10 ;
			data[55810] <= 8'h10 ;
			data[55811] <= 8'h10 ;
			data[55812] <= 8'h10 ;
			data[55813] <= 8'h10 ;
			data[55814] <= 8'h10 ;
			data[55815] <= 8'h10 ;
			data[55816] <= 8'h10 ;
			data[55817] <= 8'h10 ;
			data[55818] <= 8'h10 ;
			data[55819] <= 8'h10 ;
			data[55820] <= 8'h10 ;
			data[55821] <= 8'h10 ;
			data[55822] <= 8'h10 ;
			data[55823] <= 8'h10 ;
			data[55824] <= 8'h10 ;
			data[55825] <= 8'h10 ;
			data[55826] <= 8'h10 ;
			data[55827] <= 8'h10 ;
			data[55828] <= 8'h10 ;
			data[55829] <= 8'h10 ;
			data[55830] <= 8'h10 ;
			data[55831] <= 8'h10 ;
			data[55832] <= 8'h10 ;
			data[55833] <= 8'h10 ;
			data[55834] <= 8'h10 ;
			data[55835] <= 8'h10 ;
			data[55836] <= 8'h10 ;
			data[55837] <= 8'h10 ;
			data[55838] <= 8'h10 ;
			data[55839] <= 8'h10 ;
			data[55840] <= 8'h10 ;
			data[55841] <= 8'h10 ;
			data[55842] <= 8'h10 ;
			data[55843] <= 8'h10 ;
			data[55844] <= 8'h10 ;
			data[55845] <= 8'h10 ;
			data[55846] <= 8'h10 ;
			data[55847] <= 8'h10 ;
			data[55848] <= 8'h10 ;
			data[55849] <= 8'h10 ;
			data[55850] <= 8'h10 ;
			data[55851] <= 8'h10 ;
			data[55852] <= 8'h10 ;
			data[55853] <= 8'h10 ;
			data[55854] <= 8'h10 ;
			data[55855] <= 8'h10 ;
			data[55856] <= 8'h10 ;
			data[55857] <= 8'h10 ;
			data[55858] <= 8'h10 ;
			data[55859] <= 8'h10 ;
			data[55860] <= 8'h10 ;
			data[55861] <= 8'h10 ;
			data[55862] <= 8'h10 ;
			data[55863] <= 8'h10 ;
			data[55864] <= 8'h10 ;
			data[55865] <= 8'h10 ;
			data[55866] <= 8'h10 ;
			data[55867] <= 8'h10 ;
			data[55868] <= 8'h10 ;
			data[55869] <= 8'h10 ;
			data[55870] <= 8'h10 ;
			data[55871] <= 8'h10 ;
			data[55872] <= 8'h10 ;
			data[55873] <= 8'h10 ;
			data[55874] <= 8'h10 ;
			data[55875] <= 8'h10 ;
			data[55876] <= 8'h10 ;
			data[55877] <= 8'h10 ;
			data[55878] <= 8'h10 ;
			data[55879] <= 8'h10 ;
			data[55880] <= 8'h10 ;
			data[55881] <= 8'h10 ;
			data[55882] <= 8'h10 ;
			data[55883] <= 8'h10 ;
			data[55884] <= 8'h10 ;
			data[55885] <= 8'h10 ;
			data[55886] <= 8'h10 ;
			data[55887] <= 8'h10 ;
			data[55888] <= 8'h10 ;
			data[55889] <= 8'h10 ;
			data[55890] <= 8'h10 ;
			data[55891] <= 8'h10 ;
			data[55892] <= 8'h10 ;
			data[55893] <= 8'h10 ;
			data[55894] <= 8'h10 ;
			data[55895] <= 8'h10 ;
			data[55896] <= 8'h10 ;
			data[55897] <= 8'h10 ;
			data[55898] <= 8'h10 ;
			data[55899] <= 8'h10 ;
			data[55900] <= 8'h10 ;
			data[55901] <= 8'h10 ;
			data[55902] <= 8'h10 ;
			data[55903] <= 8'h10 ;
			data[55904] <= 8'h10 ;
			data[55905] <= 8'h10 ;
			data[55906] <= 8'h10 ;
			data[55907] <= 8'h10 ;
			data[55908] <= 8'h10 ;
			data[55909] <= 8'h10 ;
			data[55910] <= 8'h10 ;
			data[55911] <= 8'h10 ;
			data[55912] <= 8'h10 ;
			data[55913] <= 8'h10 ;
			data[55914] <= 8'h10 ;
			data[55915] <= 8'h10 ;
			data[55916] <= 8'h10 ;
			data[55917] <= 8'h10 ;
			data[55918] <= 8'h10 ;
			data[55919] <= 8'h10 ;
			data[55920] <= 8'h10 ;
			data[55921] <= 8'h10 ;
			data[55922] <= 8'h10 ;
			data[55923] <= 8'h10 ;
			data[55924] <= 8'h10 ;
			data[55925] <= 8'h10 ;
			data[55926] <= 8'h10 ;
			data[55927] <= 8'h10 ;
			data[55928] <= 8'h10 ;
			data[55929] <= 8'h10 ;
			data[55930] <= 8'h10 ;
			data[55931] <= 8'h10 ;
			data[55932] <= 8'h10 ;
			data[55933] <= 8'h10 ;
			data[55934] <= 8'h10 ;
			data[55935] <= 8'h10 ;
			data[55936] <= 8'h10 ;
			data[55937] <= 8'h10 ;
			data[55938] <= 8'h10 ;
			data[55939] <= 8'h10 ;
			data[55940] <= 8'h10 ;
			data[55941] <= 8'h10 ;
			data[55942] <= 8'h10 ;
			data[55943] <= 8'h10 ;
			data[55944] <= 8'h10 ;
			data[55945] <= 8'h10 ;
			data[55946] <= 8'h10 ;
			data[55947] <= 8'h10 ;
			data[55948] <= 8'h10 ;
			data[55949] <= 8'h10 ;
			data[55950] <= 8'h10 ;
			data[55951] <= 8'h10 ;
			data[55952] <= 8'h10 ;
			data[55953] <= 8'h10 ;
			data[55954] <= 8'h10 ;
			data[55955] <= 8'h10 ;
			data[55956] <= 8'h10 ;
			data[55957] <= 8'h10 ;
			data[55958] <= 8'h10 ;
			data[55959] <= 8'h10 ;
			data[55960] <= 8'h10 ;
			data[55961] <= 8'h10 ;
			data[55962] <= 8'h10 ;
			data[55963] <= 8'h10 ;
			data[55964] <= 8'h10 ;
			data[55965] <= 8'h10 ;
			data[55966] <= 8'h10 ;
			data[55967] <= 8'h10 ;
			data[55968] <= 8'h10 ;
			data[55969] <= 8'h10 ;
			data[55970] <= 8'h10 ;
			data[55971] <= 8'h10 ;
			data[55972] <= 8'h10 ;
			data[55973] <= 8'h10 ;
			data[55974] <= 8'h10 ;
			data[55975] <= 8'h10 ;
			data[55976] <= 8'h10 ;
			data[55977] <= 8'h10 ;
			data[55978] <= 8'h10 ;
			data[55979] <= 8'h10 ;
			data[55980] <= 8'h10 ;
			data[55981] <= 8'h10 ;
			data[55982] <= 8'h10 ;
			data[55983] <= 8'h10 ;
			data[55984] <= 8'h10 ;
			data[55985] <= 8'h10 ;
			data[55986] <= 8'h10 ;
			data[55987] <= 8'h10 ;
			data[55988] <= 8'h10 ;
			data[55989] <= 8'h10 ;
			data[55990] <= 8'h10 ;
			data[55991] <= 8'h10 ;
			data[55992] <= 8'h10 ;
			data[55993] <= 8'h10 ;
			data[55994] <= 8'h10 ;
			data[55995] <= 8'h10 ;
			data[55996] <= 8'h10 ;
			data[55997] <= 8'h10 ;
			data[55998] <= 8'h10 ;
			data[55999] <= 8'h10 ;
			data[56000] <= 8'h10 ;
			data[56001] <= 8'h10 ;
			data[56002] <= 8'h10 ;
			data[56003] <= 8'h10 ;
			data[56004] <= 8'h10 ;
			data[56005] <= 8'h10 ;
			data[56006] <= 8'h10 ;
			data[56007] <= 8'h10 ;
			data[56008] <= 8'h10 ;
			data[56009] <= 8'h10 ;
			data[56010] <= 8'h10 ;
			data[56011] <= 8'h10 ;
			data[56012] <= 8'h10 ;
			data[56013] <= 8'h10 ;
			data[56014] <= 8'h10 ;
			data[56015] <= 8'h10 ;
			data[56016] <= 8'h10 ;
			data[56017] <= 8'h10 ;
			data[56018] <= 8'h10 ;
			data[56019] <= 8'h10 ;
			data[56020] <= 8'h10 ;
			data[56021] <= 8'h10 ;
			data[56022] <= 8'h10 ;
			data[56023] <= 8'h10 ;
			data[56024] <= 8'h10 ;
			data[56025] <= 8'h10 ;
			data[56026] <= 8'h10 ;
			data[56027] <= 8'h10 ;
			data[56028] <= 8'h10 ;
			data[56029] <= 8'h10 ;
			data[56030] <= 8'h10 ;
			data[56031] <= 8'h10 ;
			data[56032] <= 8'h10 ;
			data[56033] <= 8'h10 ;
			data[56034] <= 8'h10 ;
			data[56035] <= 8'h10 ;
			data[56036] <= 8'h10 ;
			data[56037] <= 8'h10 ;
			data[56038] <= 8'h10 ;
			data[56039] <= 8'h10 ;
			data[56040] <= 8'h10 ;
			data[56041] <= 8'h10 ;
			data[56042] <= 8'h10 ;
			data[56043] <= 8'h10 ;
			data[56044] <= 8'h10 ;
			data[56045] <= 8'h10 ;
			data[56046] <= 8'h10 ;
			data[56047] <= 8'h10 ;
			data[56048] <= 8'h10 ;
			data[56049] <= 8'h10 ;
			data[56050] <= 8'h10 ;
			data[56051] <= 8'h10 ;
			data[56052] <= 8'h10 ;
			data[56053] <= 8'h10 ;
			data[56054] <= 8'h10 ;
			data[56055] <= 8'h10 ;
			data[56056] <= 8'h10 ;
			data[56057] <= 8'h10 ;
			data[56058] <= 8'h10 ;
			data[56059] <= 8'h10 ;
			data[56060] <= 8'h10 ;
			data[56061] <= 8'h10 ;
			data[56062] <= 8'h10 ;
			data[56063] <= 8'h10 ;
			data[56064] <= 8'h10 ;
			data[56065] <= 8'h10 ;
			data[56066] <= 8'h10 ;
			data[56067] <= 8'h10 ;
			data[56068] <= 8'h10 ;
			data[56069] <= 8'h10 ;
			data[56070] <= 8'h10 ;
			data[56071] <= 8'h10 ;
			data[56072] <= 8'h10 ;
			data[56073] <= 8'h10 ;
			data[56074] <= 8'h10 ;
			data[56075] <= 8'h10 ;
			data[56076] <= 8'h10 ;
			data[56077] <= 8'h10 ;
			data[56078] <= 8'h10 ;
			data[56079] <= 8'h10 ;
			data[56080] <= 8'h10 ;
			data[56081] <= 8'h10 ;
			data[56082] <= 8'h10 ;
			data[56083] <= 8'h10 ;
			data[56084] <= 8'h10 ;
			data[56085] <= 8'h10 ;
			data[56086] <= 8'h10 ;
			data[56087] <= 8'h10 ;
			data[56088] <= 8'h10 ;
			data[56089] <= 8'h10 ;
			data[56090] <= 8'h10 ;
			data[56091] <= 8'h10 ;
			data[56092] <= 8'h10 ;
			data[56093] <= 8'h10 ;
			data[56094] <= 8'h10 ;
			data[56095] <= 8'h10 ;
			data[56096] <= 8'h10 ;
			data[56097] <= 8'h10 ;
			data[56098] <= 8'h10 ;
			data[56099] <= 8'h10 ;
			data[56100] <= 8'h10 ;
			data[56101] <= 8'h10 ;
			data[56102] <= 8'h10 ;
			data[56103] <= 8'h10 ;
			data[56104] <= 8'h10 ;
			data[56105] <= 8'h10 ;
			data[56106] <= 8'h10 ;
			data[56107] <= 8'h10 ;
			data[56108] <= 8'h10 ;
			data[56109] <= 8'h10 ;
			data[56110] <= 8'h10 ;
			data[56111] <= 8'h10 ;
			data[56112] <= 8'h10 ;
			data[56113] <= 8'h10 ;
			data[56114] <= 8'h10 ;
			data[56115] <= 8'h10 ;
			data[56116] <= 8'h10 ;
			data[56117] <= 8'h10 ;
			data[56118] <= 8'h10 ;
			data[56119] <= 8'h10 ;
			data[56120] <= 8'h10 ;
			data[56121] <= 8'h10 ;
			data[56122] <= 8'h10 ;
			data[56123] <= 8'h10 ;
			data[56124] <= 8'h10 ;
			data[56125] <= 8'h10 ;
			data[56126] <= 8'h10 ;
			data[56127] <= 8'h10 ;
			data[56128] <= 8'h10 ;
			data[56129] <= 8'h10 ;
			data[56130] <= 8'h10 ;
			data[56131] <= 8'h10 ;
			data[56132] <= 8'h10 ;
			data[56133] <= 8'h10 ;
			data[56134] <= 8'h10 ;
			data[56135] <= 8'h10 ;
			data[56136] <= 8'h10 ;
			data[56137] <= 8'h10 ;
			data[56138] <= 8'h10 ;
			data[56139] <= 8'h10 ;
			data[56140] <= 8'h10 ;
			data[56141] <= 8'h10 ;
			data[56142] <= 8'h10 ;
			data[56143] <= 8'h10 ;
			data[56144] <= 8'h10 ;
			data[56145] <= 8'h10 ;
			data[56146] <= 8'h10 ;
			data[56147] <= 8'h10 ;
			data[56148] <= 8'h10 ;
			data[56149] <= 8'h10 ;
			data[56150] <= 8'h10 ;
			data[56151] <= 8'h10 ;
			data[56152] <= 8'h10 ;
			data[56153] <= 8'h10 ;
			data[56154] <= 8'h10 ;
			data[56155] <= 8'h10 ;
			data[56156] <= 8'h10 ;
			data[56157] <= 8'h10 ;
			data[56158] <= 8'h10 ;
			data[56159] <= 8'h10 ;
			data[56160] <= 8'h10 ;
			data[56161] <= 8'h10 ;
			data[56162] <= 8'h10 ;
			data[56163] <= 8'h10 ;
			data[56164] <= 8'h10 ;
			data[56165] <= 8'h10 ;
			data[56166] <= 8'h10 ;
			data[56167] <= 8'h10 ;
			data[56168] <= 8'h10 ;
			data[56169] <= 8'h10 ;
			data[56170] <= 8'h10 ;
			data[56171] <= 8'h10 ;
			data[56172] <= 8'h10 ;
			data[56173] <= 8'h10 ;
			data[56174] <= 8'h10 ;
			data[56175] <= 8'h10 ;
			data[56176] <= 8'h10 ;
			data[56177] <= 8'h10 ;
			data[56178] <= 8'h10 ;
			data[56179] <= 8'h10 ;
			data[56180] <= 8'h10 ;
			data[56181] <= 8'h10 ;
			data[56182] <= 8'h10 ;
			data[56183] <= 8'h10 ;
			data[56184] <= 8'h10 ;
			data[56185] <= 8'h10 ;
			data[56186] <= 8'h10 ;
			data[56187] <= 8'h10 ;
			data[56188] <= 8'h10 ;
			data[56189] <= 8'h10 ;
			data[56190] <= 8'h10 ;
			data[56191] <= 8'h10 ;
			data[56192] <= 8'h10 ;
			data[56193] <= 8'h10 ;
			data[56194] <= 8'h10 ;
			data[56195] <= 8'h10 ;
			data[56196] <= 8'h10 ;
			data[56197] <= 8'h10 ;
			data[56198] <= 8'h10 ;
			data[56199] <= 8'h10 ;
			data[56200] <= 8'h10 ;
			data[56201] <= 8'h10 ;
			data[56202] <= 8'h10 ;
			data[56203] <= 8'h10 ;
			data[56204] <= 8'h10 ;
			data[56205] <= 8'h10 ;
			data[56206] <= 8'h10 ;
			data[56207] <= 8'h10 ;
			data[56208] <= 8'h10 ;
			data[56209] <= 8'h10 ;
			data[56210] <= 8'h10 ;
			data[56211] <= 8'h10 ;
			data[56212] <= 8'h10 ;
			data[56213] <= 8'h10 ;
			data[56214] <= 8'h10 ;
			data[56215] <= 8'h10 ;
			data[56216] <= 8'h10 ;
			data[56217] <= 8'h10 ;
			data[56218] <= 8'h10 ;
			data[56219] <= 8'h10 ;
			data[56220] <= 8'h10 ;
			data[56221] <= 8'h10 ;
			data[56222] <= 8'h10 ;
			data[56223] <= 8'h10 ;
			data[56224] <= 8'h10 ;
			data[56225] <= 8'h10 ;
			data[56226] <= 8'h10 ;
			data[56227] <= 8'h10 ;
			data[56228] <= 8'h10 ;
			data[56229] <= 8'h10 ;
			data[56230] <= 8'h10 ;
			data[56231] <= 8'h10 ;
			data[56232] <= 8'h10 ;
			data[56233] <= 8'h10 ;
			data[56234] <= 8'h10 ;
			data[56235] <= 8'h10 ;
			data[56236] <= 8'h10 ;
			data[56237] <= 8'h10 ;
			data[56238] <= 8'h10 ;
			data[56239] <= 8'h10 ;
			data[56240] <= 8'h10 ;
			data[56241] <= 8'h10 ;
			data[56242] <= 8'h10 ;
			data[56243] <= 8'h10 ;
			data[56244] <= 8'h10 ;
			data[56245] <= 8'h10 ;
			data[56246] <= 8'h10 ;
			data[56247] <= 8'h10 ;
			data[56248] <= 8'h10 ;
			data[56249] <= 8'h10 ;
			data[56250] <= 8'h10 ;
			data[56251] <= 8'h10 ;
			data[56252] <= 8'h10 ;
			data[56253] <= 8'h10 ;
			data[56254] <= 8'h10 ;
			data[56255] <= 8'h10 ;
			data[56256] <= 8'h10 ;
			data[56257] <= 8'h10 ;
			data[56258] <= 8'h10 ;
			data[56259] <= 8'h10 ;
			data[56260] <= 8'h10 ;
			data[56261] <= 8'h10 ;
			data[56262] <= 8'h10 ;
			data[56263] <= 8'h10 ;
			data[56264] <= 8'h10 ;
			data[56265] <= 8'h10 ;
			data[56266] <= 8'h10 ;
			data[56267] <= 8'h10 ;
			data[56268] <= 8'h10 ;
			data[56269] <= 8'h10 ;
			data[56270] <= 8'h10 ;
			data[56271] <= 8'h10 ;
			data[56272] <= 8'h10 ;
			data[56273] <= 8'h10 ;
			data[56274] <= 8'h10 ;
			data[56275] <= 8'h10 ;
			data[56276] <= 8'h10 ;
			data[56277] <= 8'h10 ;
			data[56278] <= 8'h10 ;
			data[56279] <= 8'h10 ;
			data[56280] <= 8'h10 ;
			data[56281] <= 8'h10 ;
			data[56282] <= 8'h10 ;
			data[56283] <= 8'h10 ;
			data[56284] <= 8'h10 ;
			data[56285] <= 8'h10 ;
			data[56286] <= 8'h10 ;
			data[56287] <= 8'h10 ;
			data[56288] <= 8'h10 ;
			data[56289] <= 8'h10 ;
			data[56290] <= 8'h10 ;
			data[56291] <= 8'h10 ;
			data[56292] <= 8'h10 ;
			data[56293] <= 8'h10 ;
			data[56294] <= 8'h10 ;
			data[56295] <= 8'h10 ;
			data[56296] <= 8'h10 ;
			data[56297] <= 8'h10 ;
			data[56298] <= 8'h10 ;
			data[56299] <= 8'h10 ;
			data[56300] <= 8'h10 ;
			data[56301] <= 8'h10 ;
			data[56302] <= 8'h10 ;
			data[56303] <= 8'h10 ;
			data[56304] <= 8'h10 ;
			data[56305] <= 8'h10 ;
			data[56306] <= 8'h10 ;
			data[56307] <= 8'h10 ;
			data[56308] <= 8'h10 ;
			data[56309] <= 8'h10 ;
			data[56310] <= 8'h10 ;
			data[56311] <= 8'h10 ;
			data[56312] <= 8'h10 ;
			data[56313] <= 8'h10 ;
			data[56314] <= 8'h10 ;
			data[56315] <= 8'h10 ;
			data[56316] <= 8'h10 ;
			data[56317] <= 8'h10 ;
			data[56318] <= 8'h10 ;
			data[56319] <= 8'h10 ;
			data[56320] <= 8'h10 ;
			data[56321] <= 8'h10 ;
			data[56322] <= 8'h10 ;
			data[56323] <= 8'h10 ;
			data[56324] <= 8'h10 ;
			data[56325] <= 8'h10 ;
			data[56326] <= 8'h10 ;
			data[56327] <= 8'h10 ;
			data[56328] <= 8'h10 ;
			data[56329] <= 8'h10 ;
			data[56330] <= 8'h10 ;
			data[56331] <= 8'h10 ;
			data[56332] <= 8'h10 ;
			data[56333] <= 8'h10 ;
			data[56334] <= 8'h10 ;
			data[56335] <= 8'h10 ;
			data[56336] <= 8'h10 ;
			data[56337] <= 8'h10 ;
			data[56338] <= 8'h10 ;
			data[56339] <= 8'h10 ;
			data[56340] <= 8'h10 ;
			data[56341] <= 8'h10 ;
			data[56342] <= 8'h10 ;
			data[56343] <= 8'h10 ;
			data[56344] <= 8'h10 ;
			data[56345] <= 8'h10 ;
			data[56346] <= 8'h10 ;
			data[56347] <= 8'h10 ;
			data[56348] <= 8'h10 ;
			data[56349] <= 8'h10 ;
			data[56350] <= 8'h10 ;
			data[56351] <= 8'h10 ;
			data[56352] <= 8'h10 ;
			data[56353] <= 8'h10 ;
			data[56354] <= 8'h10 ;
			data[56355] <= 8'h10 ;
			data[56356] <= 8'h10 ;
			data[56357] <= 8'h10 ;
			data[56358] <= 8'h10 ;
			data[56359] <= 8'h10 ;
			data[56360] <= 8'h10 ;
			data[56361] <= 8'h10 ;
			data[56362] <= 8'h10 ;
			data[56363] <= 8'h10 ;
			data[56364] <= 8'h10 ;
			data[56365] <= 8'h10 ;
			data[56366] <= 8'h10 ;
			data[56367] <= 8'h10 ;
			data[56368] <= 8'h10 ;
			data[56369] <= 8'h10 ;
			data[56370] <= 8'h10 ;
			data[56371] <= 8'h10 ;
			data[56372] <= 8'h10 ;
			data[56373] <= 8'h10 ;
			data[56374] <= 8'h10 ;
			data[56375] <= 8'h10 ;
			data[56376] <= 8'h10 ;
			data[56377] <= 8'h10 ;
			data[56378] <= 8'h10 ;
			data[56379] <= 8'h10 ;
			data[56380] <= 8'h10 ;
			data[56381] <= 8'h10 ;
			data[56382] <= 8'h10 ;
			data[56383] <= 8'h10 ;
			data[56384] <= 8'h10 ;
			data[56385] <= 8'h10 ;
			data[56386] <= 8'h10 ;
			data[56387] <= 8'h10 ;
			data[56388] <= 8'h10 ;
			data[56389] <= 8'h10 ;
			data[56390] <= 8'h10 ;
			data[56391] <= 8'h10 ;
			data[56392] <= 8'h10 ;
			data[56393] <= 8'h10 ;
			data[56394] <= 8'h10 ;
			data[56395] <= 8'h10 ;
			data[56396] <= 8'h10 ;
			data[56397] <= 8'h10 ;
			data[56398] <= 8'h10 ;
			data[56399] <= 8'h10 ;
			data[56400] <= 8'h10 ;
			data[56401] <= 8'h10 ;
			data[56402] <= 8'h10 ;
			data[56403] <= 8'h10 ;
			data[56404] <= 8'h10 ;
			data[56405] <= 8'h10 ;
			data[56406] <= 8'h10 ;
			data[56407] <= 8'h10 ;
			data[56408] <= 8'h10 ;
			data[56409] <= 8'h10 ;
			data[56410] <= 8'h10 ;
			data[56411] <= 8'h10 ;
			data[56412] <= 8'h10 ;
			data[56413] <= 8'h10 ;
			data[56414] <= 8'h10 ;
			data[56415] <= 8'h10 ;
			data[56416] <= 8'h10 ;
			data[56417] <= 8'h10 ;
			data[56418] <= 8'h10 ;
			data[56419] <= 8'h10 ;
			data[56420] <= 8'h10 ;
			data[56421] <= 8'h10 ;
			data[56422] <= 8'h10 ;
			data[56423] <= 8'h10 ;
			data[56424] <= 8'h10 ;
			data[56425] <= 8'h10 ;
			data[56426] <= 8'h10 ;
			data[56427] <= 8'h10 ;
			data[56428] <= 8'h10 ;
			data[56429] <= 8'h10 ;
			data[56430] <= 8'h10 ;
			data[56431] <= 8'h10 ;
			data[56432] <= 8'h10 ;
			data[56433] <= 8'h10 ;
			data[56434] <= 8'h10 ;
			data[56435] <= 8'h10 ;
			data[56436] <= 8'h10 ;
			data[56437] <= 8'h10 ;
			data[56438] <= 8'h10 ;
			data[56439] <= 8'h10 ;
			data[56440] <= 8'h10 ;
			data[56441] <= 8'h10 ;
			data[56442] <= 8'h10 ;
			data[56443] <= 8'h10 ;
			data[56444] <= 8'h10 ;
			data[56445] <= 8'h10 ;
			data[56446] <= 8'h10 ;
			data[56447] <= 8'h10 ;
			data[56448] <= 8'h10 ;
			data[56449] <= 8'h10 ;
			data[56450] <= 8'h10 ;
			data[56451] <= 8'h10 ;
			data[56452] <= 8'h10 ;
			data[56453] <= 8'h10 ;
			data[56454] <= 8'h10 ;
			data[56455] <= 8'h10 ;
			data[56456] <= 8'h10 ;
			data[56457] <= 8'h10 ;
			data[56458] <= 8'h10 ;
			data[56459] <= 8'h10 ;
			data[56460] <= 8'h10 ;
			data[56461] <= 8'h10 ;
			data[56462] <= 8'h10 ;
			data[56463] <= 8'h10 ;
			data[56464] <= 8'h10 ;
			data[56465] <= 8'h10 ;
			data[56466] <= 8'h10 ;
			data[56467] <= 8'h10 ;
			data[56468] <= 8'h10 ;
			data[56469] <= 8'h10 ;
			data[56470] <= 8'h10 ;
			data[56471] <= 8'h10 ;
			data[56472] <= 8'h10 ;
			data[56473] <= 8'h10 ;
			data[56474] <= 8'h10 ;
			data[56475] <= 8'h10 ;
			data[56476] <= 8'h10 ;
			data[56477] <= 8'h10 ;
			data[56478] <= 8'h10 ;
			data[56479] <= 8'h10 ;
			data[56480] <= 8'h10 ;
			data[56481] <= 8'h10 ;
			data[56482] <= 8'h10 ;
			data[56483] <= 8'h10 ;
			data[56484] <= 8'h10 ;
			data[56485] <= 8'h10 ;
			data[56486] <= 8'h10 ;
			data[56487] <= 8'h10 ;
			data[56488] <= 8'h10 ;
			data[56489] <= 8'h10 ;
			data[56490] <= 8'h10 ;
			data[56491] <= 8'h10 ;
			data[56492] <= 8'h10 ;
			data[56493] <= 8'h10 ;
			data[56494] <= 8'h10 ;
			data[56495] <= 8'h10 ;
			data[56496] <= 8'h10 ;
			data[56497] <= 8'h10 ;
			data[56498] <= 8'h10 ;
			data[56499] <= 8'h10 ;
			data[56500] <= 8'h10 ;
			data[56501] <= 8'h10 ;
			data[56502] <= 8'h10 ;
			data[56503] <= 8'h10 ;
			data[56504] <= 8'h10 ;
			data[56505] <= 8'h10 ;
			data[56506] <= 8'h10 ;
			data[56507] <= 8'h10 ;
			data[56508] <= 8'h10 ;
			data[56509] <= 8'h10 ;
			data[56510] <= 8'h10 ;
			data[56511] <= 8'h10 ;
			data[56512] <= 8'h10 ;
			data[56513] <= 8'h10 ;
			data[56514] <= 8'h10 ;
			data[56515] <= 8'h10 ;
			data[56516] <= 8'h10 ;
			data[56517] <= 8'h10 ;
			data[56518] <= 8'h10 ;
			data[56519] <= 8'h10 ;
			data[56520] <= 8'h10 ;
			data[56521] <= 8'h10 ;
			data[56522] <= 8'h10 ;
			data[56523] <= 8'h10 ;
			data[56524] <= 8'h10 ;
			data[56525] <= 8'h10 ;
			data[56526] <= 8'h10 ;
			data[56527] <= 8'h10 ;
			data[56528] <= 8'h10 ;
			data[56529] <= 8'h10 ;
			data[56530] <= 8'h10 ;
			data[56531] <= 8'h10 ;
			data[56532] <= 8'h10 ;
			data[56533] <= 8'h10 ;
			data[56534] <= 8'h10 ;
			data[56535] <= 8'h10 ;
			data[56536] <= 8'h10 ;
			data[56537] <= 8'h10 ;
			data[56538] <= 8'h10 ;
			data[56539] <= 8'h10 ;
			data[56540] <= 8'h10 ;
			data[56541] <= 8'h10 ;
			data[56542] <= 8'h10 ;
			data[56543] <= 8'h10 ;
			data[56544] <= 8'h10 ;
			data[56545] <= 8'h10 ;
			data[56546] <= 8'h10 ;
			data[56547] <= 8'h10 ;
			data[56548] <= 8'h10 ;
			data[56549] <= 8'h10 ;
			data[56550] <= 8'h10 ;
			data[56551] <= 8'h10 ;
			data[56552] <= 8'h10 ;
			data[56553] <= 8'h10 ;
			data[56554] <= 8'h10 ;
			data[56555] <= 8'h10 ;
			data[56556] <= 8'h10 ;
			data[56557] <= 8'h10 ;
			data[56558] <= 8'h10 ;
			data[56559] <= 8'h10 ;
			data[56560] <= 8'h10 ;
			data[56561] <= 8'h10 ;
			data[56562] <= 8'h10 ;
			data[56563] <= 8'h10 ;
			data[56564] <= 8'h10 ;
			data[56565] <= 8'h10 ;
			data[56566] <= 8'h10 ;
			data[56567] <= 8'h10 ;
			data[56568] <= 8'h10 ;
			data[56569] <= 8'h10 ;
			data[56570] <= 8'h10 ;
			data[56571] <= 8'h10 ;
			data[56572] <= 8'h10 ;
			data[56573] <= 8'h10 ;
			data[56574] <= 8'h10 ;
			data[56575] <= 8'h10 ;
			data[56576] <= 8'h10 ;
			data[56577] <= 8'h10 ;
			data[56578] <= 8'h10 ;
			data[56579] <= 8'h10 ;
			data[56580] <= 8'h10 ;
			data[56581] <= 8'h10 ;
			data[56582] <= 8'h10 ;
			data[56583] <= 8'h10 ;
			data[56584] <= 8'h10 ;
			data[56585] <= 8'h10 ;
			data[56586] <= 8'h10 ;
			data[56587] <= 8'h10 ;
			data[56588] <= 8'h10 ;
			data[56589] <= 8'h10 ;
			data[56590] <= 8'h10 ;
			data[56591] <= 8'h10 ;
			data[56592] <= 8'h10 ;
			data[56593] <= 8'h10 ;
			data[56594] <= 8'h10 ;
			data[56595] <= 8'h10 ;
			data[56596] <= 8'h10 ;
			data[56597] <= 8'h10 ;
			data[56598] <= 8'h10 ;
			data[56599] <= 8'h10 ;
			data[56600] <= 8'h10 ;
			data[56601] <= 8'h10 ;
			data[56602] <= 8'h10 ;
			data[56603] <= 8'h10 ;
			data[56604] <= 8'h10 ;
			data[56605] <= 8'h10 ;
			data[56606] <= 8'h10 ;
			data[56607] <= 8'h10 ;
			data[56608] <= 8'h10 ;
			data[56609] <= 8'h10 ;
			data[56610] <= 8'h10 ;
			data[56611] <= 8'h10 ;
			data[56612] <= 8'h10 ;
			data[56613] <= 8'h10 ;
			data[56614] <= 8'h10 ;
			data[56615] <= 8'h10 ;
			data[56616] <= 8'h10 ;
			data[56617] <= 8'h10 ;
			data[56618] <= 8'h10 ;
			data[56619] <= 8'h10 ;
			data[56620] <= 8'h10 ;
			data[56621] <= 8'h10 ;
			data[56622] <= 8'h10 ;
			data[56623] <= 8'h10 ;
			data[56624] <= 8'h10 ;
			data[56625] <= 8'h10 ;
			data[56626] <= 8'h10 ;
			data[56627] <= 8'h10 ;
			data[56628] <= 8'h10 ;
			data[56629] <= 8'h10 ;
			data[56630] <= 8'h10 ;
			data[56631] <= 8'h10 ;
			data[56632] <= 8'h10 ;
			data[56633] <= 8'h10 ;
			data[56634] <= 8'h10 ;
			data[56635] <= 8'h10 ;
			data[56636] <= 8'h10 ;
			data[56637] <= 8'h10 ;
			data[56638] <= 8'h10 ;
			data[56639] <= 8'h10 ;
			data[56640] <= 8'h10 ;
			data[56641] <= 8'h10 ;
			data[56642] <= 8'h10 ;
			data[56643] <= 8'h10 ;
			data[56644] <= 8'h10 ;
			data[56645] <= 8'h10 ;
			data[56646] <= 8'h10 ;
			data[56647] <= 8'h10 ;
			data[56648] <= 8'h10 ;
			data[56649] <= 8'h10 ;
			data[56650] <= 8'h10 ;
			data[56651] <= 8'h10 ;
			data[56652] <= 8'h10 ;
			data[56653] <= 8'h10 ;
			data[56654] <= 8'h10 ;
			data[56655] <= 8'h10 ;
			data[56656] <= 8'h10 ;
			data[56657] <= 8'h10 ;
			data[56658] <= 8'h10 ;
			data[56659] <= 8'h10 ;
			data[56660] <= 8'h10 ;
			data[56661] <= 8'h10 ;
			data[56662] <= 8'h10 ;
			data[56663] <= 8'h10 ;
			data[56664] <= 8'h10 ;
			data[56665] <= 8'h10 ;
			data[56666] <= 8'h10 ;
			data[56667] <= 8'h10 ;
			data[56668] <= 8'h10 ;
			data[56669] <= 8'h10 ;
			data[56670] <= 8'h10 ;
			data[56671] <= 8'h10 ;
			data[56672] <= 8'h10 ;
			data[56673] <= 8'h10 ;
			data[56674] <= 8'h10 ;
			data[56675] <= 8'h10 ;
			data[56676] <= 8'h10 ;
			data[56677] <= 8'h10 ;
			data[56678] <= 8'h10 ;
			data[56679] <= 8'h10 ;
			data[56680] <= 8'h10 ;
			data[56681] <= 8'h10 ;
			data[56682] <= 8'h10 ;
			data[56683] <= 8'h10 ;
			data[56684] <= 8'h10 ;
			data[56685] <= 8'h10 ;
			data[56686] <= 8'h10 ;
			data[56687] <= 8'h10 ;
			data[56688] <= 8'h10 ;
			data[56689] <= 8'h10 ;
			data[56690] <= 8'h10 ;
			data[56691] <= 8'h10 ;
			data[56692] <= 8'h10 ;
			data[56693] <= 8'h10 ;
			data[56694] <= 8'h10 ;
			data[56695] <= 8'h10 ;
			data[56696] <= 8'h10 ;
			data[56697] <= 8'h10 ;
			data[56698] <= 8'h10 ;
			data[56699] <= 8'h10 ;
			data[56700] <= 8'h10 ;
			data[56701] <= 8'h10 ;
			data[56702] <= 8'h10 ;
			data[56703] <= 8'h10 ;
			data[56704] <= 8'h10 ;
			data[56705] <= 8'h10 ;
			data[56706] <= 8'h10 ;
			data[56707] <= 8'h10 ;
			data[56708] <= 8'h10 ;
			data[56709] <= 8'h10 ;
			data[56710] <= 8'h10 ;
			data[56711] <= 8'h10 ;
			data[56712] <= 8'h10 ;
			data[56713] <= 8'h10 ;
			data[56714] <= 8'h10 ;
			data[56715] <= 8'h10 ;
			data[56716] <= 8'h10 ;
			data[56717] <= 8'h10 ;
			data[56718] <= 8'h10 ;
			data[56719] <= 8'h10 ;
			data[56720] <= 8'h10 ;
			data[56721] <= 8'h10 ;
			data[56722] <= 8'h10 ;
			data[56723] <= 8'h10 ;
			data[56724] <= 8'h10 ;
			data[56725] <= 8'h10 ;
			data[56726] <= 8'h10 ;
			data[56727] <= 8'h10 ;
			data[56728] <= 8'h10 ;
			data[56729] <= 8'h10 ;
			data[56730] <= 8'h10 ;
			data[56731] <= 8'h10 ;
			data[56732] <= 8'h10 ;
			data[56733] <= 8'h10 ;
			data[56734] <= 8'h10 ;
			data[56735] <= 8'h10 ;
			data[56736] <= 8'h10 ;
			data[56737] <= 8'h10 ;
			data[56738] <= 8'h10 ;
			data[56739] <= 8'h10 ;
			data[56740] <= 8'h10 ;
			data[56741] <= 8'h10 ;
			data[56742] <= 8'h10 ;
			data[56743] <= 8'h10 ;
			data[56744] <= 8'h10 ;
			data[56745] <= 8'h10 ;
			data[56746] <= 8'h10 ;
			data[56747] <= 8'h10 ;
			data[56748] <= 8'h10 ;
			data[56749] <= 8'h10 ;
			data[56750] <= 8'h10 ;
			data[56751] <= 8'h10 ;
			data[56752] <= 8'h10 ;
			data[56753] <= 8'h10 ;
			data[56754] <= 8'h10 ;
			data[56755] <= 8'h10 ;
			data[56756] <= 8'h10 ;
			data[56757] <= 8'h10 ;
			data[56758] <= 8'h10 ;
			data[56759] <= 8'h10 ;
			data[56760] <= 8'h10 ;
			data[56761] <= 8'h10 ;
			data[56762] <= 8'h10 ;
			data[56763] <= 8'h10 ;
			data[56764] <= 8'h10 ;
			data[56765] <= 8'h10 ;
			data[56766] <= 8'h10 ;
			data[56767] <= 8'h10 ;
			data[56768] <= 8'h10 ;
			data[56769] <= 8'h10 ;
			data[56770] <= 8'h10 ;
			data[56771] <= 8'h10 ;
			data[56772] <= 8'h10 ;
			data[56773] <= 8'h10 ;
			data[56774] <= 8'h10 ;
			data[56775] <= 8'h10 ;
			data[56776] <= 8'h10 ;
			data[56777] <= 8'h10 ;
			data[56778] <= 8'h10 ;
			data[56779] <= 8'h10 ;
			data[56780] <= 8'h10 ;
			data[56781] <= 8'h10 ;
			data[56782] <= 8'h10 ;
			data[56783] <= 8'h10 ;
			data[56784] <= 8'h10 ;
			data[56785] <= 8'h10 ;
			data[56786] <= 8'h10 ;
			data[56787] <= 8'h10 ;
			data[56788] <= 8'h10 ;
			data[56789] <= 8'h10 ;
			data[56790] <= 8'h10 ;
			data[56791] <= 8'h10 ;
			data[56792] <= 8'h10 ;
			data[56793] <= 8'h10 ;
			data[56794] <= 8'h10 ;
			data[56795] <= 8'h10 ;
			data[56796] <= 8'h10 ;
			data[56797] <= 8'h10 ;
			data[56798] <= 8'h10 ;
			data[56799] <= 8'h10 ;
			data[56800] <= 8'h10 ;
			data[56801] <= 8'h10 ;
			data[56802] <= 8'h10 ;
			data[56803] <= 8'h10 ;
			data[56804] <= 8'h10 ;
			data[56805] <= 8'h10 ;
			data[56806] <= 8'h10 ;
			data[56807] <= 8'h10 ;
			data[56808] <= 8'h10 ;
			data[56809] <= 8'h10 ;
			data[56810] <= 8'h10 ;
			data[56811] <= 8'h10 ;
			data[56812] <= 8'h10 ;
			data[56813] <= 8'h10 ;
			data[56814] <= 8'h10 ;
			data[56815] <= 8'h10 ;
			data[56816] <= 8'h10 ;
			data[56817] <= 8'h10 ;
			data[56818] <= 8'h10 ;
			data[56819] <= 8'h10 ;
			data[56820] <= 8'h10 ;
			data[56821] <= 8'h10 ;
			data[56822] <= 8'h10 ;
			data[56823] <= 8'h10 ;
			data[56824] <= 8'h10 ;
			data[56825] <= 8'h10 ;
			data[56826] <= 8'h10 ;
			data[56827] <= 8'h10 ;
			data[56828] <= 8'h10 ;
			data[56829] <= 8'h10 ;
			data[56830] <= 8'h10 ;
			data[56831] <= 8'h10 ;
			data[56832] <= 8'h10 ;
			data[56833] <= 8'h10 ;
			data[56834] <= 8'h10 ;
			data[56835] <= 8'h10 ;
			data[56836] <= 8'h10 ;
			data[56837] <= 8'h10 ;
			data[56838] <= 8'h10 ;
			data[56839] <= 8'h10 ;
			data[56840] <= 8'h10 ;
			data[56841] <= 8'h10 ;
			data[56842] <= 8'h10 ;
			data[56843] <= 8'h10 ;
			data[56844] <= 8'h10 ;
			data[56845] <= 8'h10 ;
			data[56846] <= 8'h10 ;
			data[56847] <= 8'h10 ;
			data[56848] <= 8'h10 ;
			data[56849] <= 8'h10 ;
			data[56850] <= 8'h10 ;
			data[56851] <= 8'h10 ;
			data[56852] <= 8'h10 ;
			data[56853] <= 8'h10 ;
			data[56854] <= 8'h10 ;
			data[56855] <= 8'h10 ;
			data[56856] <= 8'h10 ;
			data[56857] <= 8'h10 ;
			data[56858] <= 8'h10 ;
			data[56859] <= 8'h10 ;
			data[56860] <= 8'h10 ;
			data[56861] <= 8'h10 ;
			data[56862] <= 8'h10 ;
			data[56863] <= 8'h10 ;
			data[56864] <= 8'h10 ;
			data[56865] <= 8'h10 ;
			data[56866] <= 8'h10 ;
			data[56867] <= 8'h10 ;
			data[56868] <= 8'h10 ;
			data[56869] <= 8'h10 ;
			data[56870] <= 8'h10 ;
			data[56871] <= 8'h10 ;
			data[56872] <= 8'h10 ;
			data[56873] <= 8'h10 ;
			data[56874] <= 8'h10 ;
			data[56875] <= 8'h10 ;
			data[56876] <= 8'h10 ;
			data[56877] <= 8'h10 ;
			data[56878] <= 8'h10 ;
			data[56879] <= 8'h10 ;
			data[56880] <= 8'h10 ;
			data[56881] <= 8'h10 ;
			data[56882] <= 8'h10 ;
			data[56883] <= 8'h10 ;
			data[56884] <= 8'h10 ;
			data[56885] <= 8'h10 ;
			data[56886] <= 8'h10 ;
			data[56887] <= 8'h10 ;
			data[56888] <= 8'h10 ;
			data[56889] <= 8'h10 ;
			data[56890] <= 8'h10 ;
			data[56891] <= 8'h10 ;
			data[56892] <= 8'h10 ;
			data[56893] <= 8'h10 ;
			data[56894] <= 8'h10 ;
			data[56895] <= 8'h10 ;
			data[56896] <= 8'h10 ;
			data[56897] <= 8'h10 ;
			data[56898] <= 8'h10 ;
			data[56899] <= 8'h10 ;
			data[56900] <= 8'h10 ;
			data[56901] <= 8'h10 ;
			data[56902] <= 8'h10 ;
			data[56903] <= 8'h10 ;
			data[56904] <= 8'h10 ;
			data[56905] <= 8'h10 ;
			data[56906] <= 8'h10 ;
			data[56907] <= 8'h10 ;
			data[56908] <= 8'h10 ;
			data[56909] <= 8'h10 ;
			data[56910] <= 8'h10 ;
			data[56911] <= 8'h10 ;
			data[56912] <= 8'h10 ;
			data[56913] <= 8'h10 ;
			data[56914] <= 8'h10 ;
			data[56915] <= 8'h10 ;
			data[56916] <= 8'h10 ;
			data[56917] <= 8'h10 ;
			data[56918] <= 8'h10 ;
			data[56919] <= 8'h10 ;
			data[56920] <= 8'h10 ;
			data[56921] <= 8'h10 ;
			data[56922] <= 8'h10 ;
			data[56923] <= 8'h10 ;
			data[56924] <= 8'h10 ;
			data[56925] <= 8'h10 ;
			data[56926] <= 8'h10 ;
			data[56927] <= 8'h10 ;
			data[56928] <= 8'h10 ;
			data[56929] <= 8'h10 ;
			data[56930] <= 8'h10 ;
			data[56931] <= 8'h10 ;
			data[56932] <= 8'h10 ;
			data[56933] <= 8'h10 ;
			data[56934] <= 8'h10 ;
			data[56935] <= 8'h10 ;
			data[56936] <= 8'h10 ;
			data[56937] <= 8'h10 ;
			data[56938] <= 8'h10 ;
			data[56939] <= 8'h10 ;
			data[56940] <= 8'h10 ;
			data[56941] <= 8'h10 ;
			data[56942] <= 8'h10 ;
			data[56943] <= 8'h10 ;
			data[56944] <= 8'h10 ;
			data[56945] <= 8'h10 ;
			data[56946] <= 8'h10 ;
			data[56947] <= 8'h10 ;
			data[56948] <= 8'h10 ;
			data[56949] <= 8'h10 ;
			data[56950] <= 8'h10 ;
			data[56951] <= 8'h10 ;
			data[56952] <= 8'h10 ;
			data[56953] <= 8'h10 ;
			data[56954] <= 8'h10 ;
			data[56955] <= 8'h10 ;
			data[56956] <= 8'h10 ;
			data[56957] <= 8'h10 ;
			data[56958] <= 8'h10 ;
			data[56959] <= 8'h10 ;
			data[56960] <= 8'h10 ;
			data[56961] <= 8'h10 ;
			data[56962] <= 8'h10 ;
			data[56963] <= 8'h10 ;
			data[56964] <= 8'h10 ;
			data[56965] <= 8'h10 ;
			data[56966] <= 8'h10 ;
			data[56967] <= 8'h10 ;
			data[56968] <= 8'h10 ;
			data[56969] <= 8'h10 ;
			data[56970] <= 8'h10 ;
			data[56971] <= 8'h10 ;
			data[56972] <= 8'h10 ;
			data[56973] <= 8'h10 ;
			data[56974] <= 8'h10 ;
			data[56975] <= 8'h10 ;
			data[56976] <= 8'h10 ;
			data[56977] <= 8'h10 ;
			data[56978] <= 8'h10 ;
			data[56979] <= 8'h10 ;
			data[56980] <= 8'h10 ;
			data[56981] <= 8'h10 ;
			data[56982] <= 8'h10 ;
			data[56983] <= 8'h10 ;
			data[56984] <= 8'h10 ;
			data[56985] <= 8'h10 ;
			data[56986] <= 8'h10 ;
			data[56987] <= 8'h10 ;
			data[56988] <= 8'h10 ;
			data[56989] <= 8'h10 ;
			data[56990] <= 8'h10 ;
			data[56991] <= 8'h10 ;
			data[56992] <= 8'h10 ;
			data[56993] <= 8'h10 ;
			data[56994] <= 8'h10 ;
			data[56995] <= 8'h10 ;
			data[56996] <= 8'h10 ;
			data[56997] <= 8'h10 ;
			data[56998] <= 8'h10 ;
			data[56999] <= 8'h10 ;
			data[57000] <= 8'h10 ;
			data[57001] <= 8'h10 ;
			data[57002] <= 8'h10 ;
			data[57003] <= 8'h10 ;
			data[57004] <= 8'h10 ;
			data[57005] <= 8'h10 ;
			data[57006] <= 8'h10 ;
			data[57007] <= 8'h10 ;
			data[57008] <= 8'h10 ;
			data[57009] <= 8'h10 ;
			data[57010] <= 8'h10 ;
			data[57011] <= 8'h10 ;
			data[57012] <= 8'h10 ;
			data[57013] <= 8'h10 ;
			data[57014] <= 8'h10 ;
			data[57015] <= 8'h10 ;
			data[57016] <= 8'h10 ;
			data[57017] <= 8'h10 ;
			data[57018] <= 8'h10 ;
			data[57019] <= 8'h10 ;
			data[57020] <= 8'h10 ;
			data[57021] <= 8'h10 ;
			data[57022] <= 8'h10 ;
			data[57023] <= 8'h10 ;
			data[57024] <= 8'h10 ;
			data[57025] <= 8'h10 ;
			data[57026] <= 8'h10 ;
			data[57027] <= 8'h10 ;
			data[57028] <= 8'h10 ;
			data[57029] <= 8'h10 ;
			data[57030] <= 8'h10 ;
			data[57031] <= 8'h10 ;
			data[57032] <= 8'h10 ;
			data[57033] <= 8'h10 ;
			data[57034] <= 8'h10 ;
			data[57035] <= 8'h10 ;
			data[57036] <= 8'h10 ;
			data[57037] <= 8'h10 ;
			data[57038] <= 8'h10 ;
			data[57039] <= 8'h10 ;
			data[57040] <= 8'h10 ;
			data[57041] <= 8'h10 ;
			data[57042] <= 8'h10 ;
			data[57043] <= 8'h10 ;
			data[57044] <= 8'h10 ;
			data[57045] <= 8'h10 ;
			data[57046] <= 8'h10 ;
			data[57047] <= 8'h10 ;
			data[57048] <= 8'h10 ;
			data[57049] <= 8'h10 ;
			data[57050] <= 8'h10 ;
			data[57051] <= 8'h10 ;
			data[57052] <= 8'h10 ;
			data[57053] <= 8'h10 ;
			data[57054] <= 8'h10 ;
			data[57055] <= 8'h10 ;
			data[57056] <= 8'h10 ;
			data[57057] <= 8'h10 ;
			data[57058] <= 8'h10 ;
			data[57059] <= 8'h10 ;
			data[57060] <= 8'h10 ;
			data[57061] <= 8'h10 ;
			data[57062] <= 8'h10 ;
			data[57063] <= 8'h10 ;
			data[57064] <= 8'h10 ;
			data[57065] <= 8'h10 ;
			data[57066] <= 8'h10 ;
			data[57067] <= 8'h10 ;
			data[57068] <= 8'h10 ;
			data[57069] <= 8'h10 ;
			data[57070] <= 8'h10 ;
			data[57071] <= 8'h10 ;
			data[57072] <= 8'h10 ;
			data[57073] <= 8'h10 ;
			data[57074] <= 8'h10 ;
			data[57075] <= 8'h10 ;
			data[57076] <= 8'h10 ;
			data[57077] <= 8'h10 ;
			data[57078] <= 8'h10 ;
			data[57079] <= 8'h10 ;
			data[57080] <= 8'h10 ;
			data[57081] <= 8'h10 ;
			data[57082] <= 8'h10 ;
			data[57083] <= 8'h10 ;
			data[57084] <= 8'h10 ;
			data[57085] <= 8'h10 ;
			data[57086] <= 8'h10 ;
			data[57087] <= 8'h10 ;
			data[57088] <= 8'h10 ;
			data[57089] <= 8'h10 ;
			data[57090] <= 8'h10 ;
			data[57091] <= 8'h10 ;
			data[57092] <= 8'h10 ;
			data[57093] <= 8'h10 ;
			data[57094] <= 8'h10 ;
			data[57095] <= 8'h10 ;
			data[57096] <= 8'h10 ;
			data[57097] <= 8'h10 ;
			data[57098] <= 8'h10 ;
			data[57099] <= 8'h10 ;
			data[57100] <= 8'h10 ;
			data[57101] <= 8'h10 ;
			data[57102] <= 8'h10 ;
			data[57103] <= 8'h10 ;
			data[57104] <= 8'h10 ;
			data[57105] <= 8'h10 ;
			data[57106] <= 8'h10 ;
			data[57107] <= 8'h10 ;
			data[57108] <= 8'h10 ;
			data[57109] <= 8'h10 ;
			data[57110] <= 8'h10 ;
			data[57111] <= 8'h10 ;
			data[57112] <= 8'h10 ;
			data[57113] <= 8'h10 ;
			data[57114] <= 8'h10 ;
			data[57115] <= 8'h10 ;
			data[57116] <= 8'h10 ;
			data[57117] <= 8'h10 ;
			data[57118] <= 8'h10 ;
			data[57119] <= 8'h10 ;
			data[57120] <= 8'h10 ;
			data[57121] <= 8'h10 ;
			data[57122] <= 8'h10 ;
			data[57123] <= 8'h10 ;
			data[57124] <= 8'h10 ;
			data[57125] <= 8'h10 ;
			data[57126] <= 8'h10 ;
			data[57127] <= 8'h10 ;
			data[57128] <= 8'h10 ;
			data[57129] <= 8'h10 ;
			data[57130] <= 8'h10 ;
			data[57131] <= 8'h10 ;
			data[57132] <= 8'h10 ;
			data[57133] <= 8'h10 ;
			data[57134] <= 8'h10 ;
			data[57135] <= 8'h10 ;
			data[57136] <= 8'h10 ;
			data[57137] <= 8'h10 ;
			data[57138] <= 8'h10 ;
			data[57139] <= 8'h10 ;
			data[57140] <= 8'h10 ;
			data[57141] <= 8'h10 ;
			data[57142] <= 8'h10 ;
			data[57143] <= 8'h10 ;
			data[57144] <= 8'h10 ;
			data[57145] <= 8'h10 ;
			data[57146] <= 8'h10 ;
			data[57147] <= 8'h10 ;
			data[57148] <= 8'h10 ;
			data[57149] <= 8'h10 ;
			data[57150] <= 8'h10 ;
			data[57151] <= 8'h10 ;
			data[57152] <= 8'h10 ;
			data[57153] <= 8'h10 ;
			data[57154] <= 8'h10 ;
			data[57155] <= 8'h10 ;
			data[57156] <= 8'h10 ;
			data[57157] <= 8'h10 ;
			data[57158] <= 8'h10 ;
			data[57159] <= 8'h10 ;
			data[57160] <= 8'h10 ;
			data[57161] <= 8'h10 ;
			data[57162] <= 8'h10 ;
			data[57163] <= 8'h10 ;
			data[57164] <= 8'h10 ;
			data[57165] <= 8'h10 ;
			data[57166] <= 8'h10 ;
			data[57167] <= 8'h10 ;
			data[57168] <= 8'h10 ;
			data[57169] <= 8'h10 ;
			data[57170] <= 8'h10 ;
			data[57171] <= 8'h10 ;
			data[57172] <= 8'h10 ;
			data[57173] <= 8'h10 ;
			data[57174] <= 8'h10 ;
			data[57175] <= 8'h10 ;
			data[57176] <= 8'h10 ;
			data[57177] <= 8'h10 ;
			data[57178] <= 8'h10 ;
			data[57179] <= 8'h10 ;
			data[57180] <= 8'h10 ;
			data[57181] <= 8'h10 ;
			data[57182] <= 8'h10 ;
			data[57183] <= 8'h10 ;
			data[57184] <= 8'h10 ;
			data[57185] <= 8'h10 ;
			data[57186] <= 8'h10 ;
			data[57187] <= 8'h10 ;
			data[57188] <= 8'h10 ;
			data[57189] <= 8'h10 ;
			data[57190] <= 8'h10 ;
			data[57191] <= 8'h10 ;
			data[57192] <= 8'h10 ;
			data[57193] <= 8'h10 ;
			data[57194] <= 8'h10 ;
			data[57195] <= 8'h10 ;
			data[57196] <= 8'h10 ;
			data[57197] <= 8'h10 ;
			data[57198] <= 8'h10 ;
			data[57199] <= 8'h10 ;
			data[57200] <= 8'h10 ;
			data[57201] <= 8'h10 ;
			data[57202] <= 8'h10 ;
			data[57203] <= 8'h10 ;
			data[57204] <= 8'h10 ;
			data[57205] <= 8'h10 ;
			data[57206] <= 8'h10 ;
			data[57207] <= 8'h10 ;
			data[57208] <= 8'h10 ;
			data[57209] <= 8'h10 ;
			data[57210] <= 8'h10 ;
			data[57211] <= 8'h10 ;
			data[57212] <= 8'h10 ;
			data[57213] <= 8'h10 ;
			data[57214] <= 8'h10 ;
			data[57215] <= 8'h10 ;
			data[57216] <= 8'h10 ;
			data[57217] <= 8'h10 ;
			data[57218] <= 8'h10 ;
			data[57219] <= 8'h10 ;
			data[57220] <= 8'h10 ;
			data[57221] <= 8'h10 ;
			data[57222] <= 8'h10 ;
			data[57223] <= 8'h10 ;
			data[57224] <= 8'h10 ;
			data[57225] <= 8'h10 ;
			data[57226] <= 8'h10 ;
			data[57227] <= 8'h10 ;
			data[57228] <= 8'h10 ;
			data[57229] <= 8'h10 ;
			data[57230] <= 8'h10 ;
			data[57231] <= 8'h10 ;
			data[57232] <= 8'h10 ;
			data[57233] <= 8'h10 ;
			data[57234] <= 8'h10 ;
			data[57235] <= 8'h10 ;
			data[57236] <= 8'h10 ;
			data[57237] <= 8'h10 ;
			data[57238] <= 8'h10 ;
			data[57239] <= 8'h10 ;
			data[57240] <= 8'h10 ;
			data[57241] <= 8'h10 ;
			data[57242] <= 8'h10 ;
			data[57243] <= 8'h10 ;
			data[57244] <= 8'h10 ;
			data[57245] <= 8'h10 ;
			data[57246] <= 8'h10 ;
			data[57247] <= 8'h10 ;
			data[57248] <= 8'h10 ;
			data[57249] <= 8'h10 ;
			data[57250] <= 8'h10 ;
			data[57251] <= 8'h10 ;
			data[57252] <= 8'h10 ;
			data[57253] <= 8'h10 ;
			data[57254] <= 8'h10 ;
			data[57255] <= 8'h10 ;
			data[57256] <= 8'h10 ;
			data[57257] <= 8'h10 ;
			data[57258] <= 8'h10 ;
			data[57259] <= 8'h10 ;
			data[57260] <= 8'h10 ;
			data[57261] <= 8'h10 ;
			data[57262] <= 8'h10 ;
			data[57263] <= 8'h10 ;
			data[57264] <= 8'h10 ;
			data[57265] <= 8'h10 ;
			data[57266] <= 8'h10 ;
			data[57267] <= 8'h10 ;
			data[57268] <= 8'h10 ;
			data[57269] <= 8'h10 ;
			data[57270] <= 8'h10 ;
			data[57271] <= 8'h10 ;
			data[57272] <= 8'h10 ;
			data[57273] <= 8'h10 ;
			data[57274] <= 8'h10 ;
			data[57275] <= 8'h10 ;
			data[57276] <= 8'h10 ;
			data[57277] <= 8'h10 ;
			data[57278] <= 8'h10 ;
			data[57279] <= 8'h10 ;
			data[57280] <= 8'h10 ;
			data[57281] <= 8'h10 ;
			data[57282] <= 8'h10 ;
			data[57283] <= 8'h10 ;
			data[57284] <= 8'h10 ;
			data[57285] <= 8'h10 ;
			data[57286] <= 8'h10 ;
			data[57287] <= 8'h10 ;
			data[57288] <= 8'h10 ;
			data[57289] <= 8'h10 ;
			data[57290] <= 8'h10 ;
			data[57291] <= 8'h10 ;
			data[57292] <= 8'h10 ;
			data[57293] <= 8'h10 ;
			data[57294] <= 8'h10 ;
			data[57295] <= 8'h10 ;
			data[57296] <= 8'h10 ;
			data[57297] <= 8'h10 ;
			data[57298] <= 8'h10 ;
			data[57299] <= 8'h10 ;
			data[57300] <= 8'h10 ;
			data[57301] <= 8'h10 ;
			data[57302] <= 8'h10 ;
			data[57303] <= 8'h10 ;
			data[57304] <= 8'h10 ;
			data[57305] <= 8'h10 ;
			data[57306] <= 8'h10 ;
			data[57307] <= 8'h10 ;
			data[57308] <= 8'h10 ;
			data[57309] <= 8'h10 ;
			data[57310] <= 8'h10 ;
			data[57311] <= 8'h10 ;
			data[57312] <= 8'h10 ;
			data[57313] <= 8'h10 ;
			data[57314] <= 8'h10 ;
			data[57315] <= 8'h10 ;
			data[57316] <= 8'h10 ;
			data[57317] <= 8'h10 ;
			data[57318] <= 8'h10 ;
			data[57319] <= 8'h10 ;
			data[57320] <= 8'h10 ;
			data[57321] <= 8'h10 ;
			data[57322] <= 8'h10 ;
			data[57323] <= 8'h10 ;
			data[57324] <= 8'h10 ;
			data[57325] <= 8'h10 ;
			data[57326] <= 8'h10 ;
			data[57327] <= 8'h10 ;
			data[57328] <= 8'h10 ;
			data[57329] <= 8'h10 ;
			data[57330] <= 8'h10 ;
			data[57331] <= 8'h10 ;
			data[57332] <= 8'h10 ;
			data[57333] <= 8'h10 ;
			data[57334] <= 8'h10 ;
			data[57335] <= 8'h10 ;
			data[57336] <= 8'h10 ;
			data[57337] <= 8'h10 ;
			data[57338] <= 8'h10 ;
			data[57339] <= 8'h10 ;
			data[57340] <= 8'h10 ;
			data[57341] <= 8'h10 ;
			data[57342] <= 8'h10 ;
			data[57343] <= 8'h10 ;
			data[57344] <= 8'h10 ;
			data[57345] <= 8'h10 ;
			data[57346] <= 8'h10 ;
			data[57347] <= 8'h10 ;
			data[57348] <= 8'h10 ;
			data[57349] <= 8'h10 ;
			data[57350] <= 8'h10 ;
			data[57351] <= 8'h10 ;
			data[57352] <= 8'h10 ;
			data[57353] <= 8'h10 ;
			data[57354] <= 8'h10 ;
			data[57355] <= 8'h10 ;
			data[57356] <= 8'h10 ;
			data[57357] <= 8'h10 ;
			data[57358] <= 8'h10 ;
			data[57359] <= 8'h10 ;
			data[57360] <= 8'h10 ;
			data[57361] <= 8'h10 ;
			data[57362] <= 8'h10 ;
			data[57363] <= 8'h10 ;
			data[57364] <= 8'h10 ;
			data[57365] <= 8'h10 ;
			data[57366] <= 8'h10 ;
			data[57367] <= 8'h10 ;
			data[57368] <= 8'h10 ;
			data[57369] <= 8'h10 ;
			data[57370] <= 8'h10 ;
			data[57371] <= 8'h10 ;
			data[57372] <= 8'h10 ;
			data[57373] <= 8'h10 ;
			data[57374] <= 8'h10 ;
			data[57375] <= 8'h10 ;
			data[57376] <= 8'h10 ;
			data[57377] <= 8'h10 ;
			data[57378] <= 8'h10 ;
			data[57379] <= 8'h10 ;
			data[57380] <= 8'h10 ;
			data[57381] <= 8'h10 ;
			data[57382] <= 8'h10 ;
			data[57383] <= 8'h10 ;
			data[57384] <= 8'h10 ;
			data[57385] <= 8'h10 ;
			data[57386] <= 8'h10 ;
			data[57387] <= 8'h10 ;
			data[57388] <= 8'h10 ;
			data[57389] <= 8'h10 ;
			data[57390] <= 8'h10 ;
			data[57391] <= 8'h10 ;
			data[57392] <= 8'h10 ;
			data[57393] <= 8'h10 ;
			data[57394] <= 8'h10 ;
			data[57395] <= 8'h10 ;
			data[57396] <= 8'h10 ;
			data[57397] <= 8'h10 ;
			data[57398] <= 8'h10 ;
			data[57399] <= 8'h10 ;
			data[57400] <= 8'h10 ;
			data[57401] <= 8'h10 ;
			data[57402] <= 8'h10 ;
			data[57403] <= 8'h10 ;
			data[57404] <= 8'h10 ;
			data[57405] <= 8'h10 ;
			data[57406] <= 8'h10 ;
			data[57407] <= 8'h10 ;
			data[57408] <= 8'h10 ;
			data[57409] <= 8'h10 ;
			data[57410] <= 8'h10 ;
			data[57411] <= 8'h10 ;
			data[57412] <= 8'h10 ;
			data[57413] <= 8'h10 ;
			data[57414] <= 8'h10 ;
			data[57415] <= 8'h10 ;
			data[57416] <= 8'h10 ;
			data[57417] <= 8'h10 ;
			data[57418] <= 8'h10 ;
			data[57419] <= 8'h10 ;
			data[57420] <= 8'h10 ;
			data[57421] <= 8'h10 ;
			data[57422] <= 8'h10 ;
			data[57423] <= 8'h10 ;
			data[57424] <= 8'h10 ;
			data[57425] <= 8'h10 ;
			data[57426] <= 8'h10 ;
			data[57427] <= 8'h10 ;
			data[57428] <= 8'h10 ;
			data[57429] <= 8'h10 ;
			data[57430] <= 8'h10 ;
			data[57431] <= 8'h10 ;
			data[57432] <= 8'h10 ;
			data[57433] <= 8'h10 ;
			data[57434] <= 8'h10 ;
			data[57435] <= 8'h10 ;
			data[57436] <= 8'h10 ;
			data[57437] <= 8'h10 ;
			data[57438] <= 8'h10 ;
			data[57439] <= 8'h10 ;
			data[57440] <= 8'h10 ;
			data[57441] <= 8'h10 ;
			data[57442] <= 8'h10 ;
			data[57443] <= 8'h10 ;
			data[57444] <= 8'h10 ;
			data[57445] <= 8'h10 ;
			data[57446] <= 8'h10 ;
			data[57447] <= 8'h10 ;
			data[57448] <= 8'h10 ;
			data[57449] <= 8'h10 ;
			data[57450] <= 8'h10 ;
			data[57451] <= 8'h10 ;
			data[57452] <= 8'h10 ;
			data[57453] <= 8'h10 ;
			data[57454] <= 8'h10 ;
			data[57455] <= 8'h10 ;
			data[57456] <= 8'h10 ;
			data[57457] <= 8'h10 ;
			data[57458] <= 8'h10 ;
			data[57459] <= 8'h10 ;
			data[57460] <= 8'h10 ;
			data[57461] <= 8'h10 ;
			data[57462] <= 8'h10 ;
			data[57463] <= 8'h10 ;
			data[57464] <= 8'h10 ;
			data[57465] <= 8'h10 ;
			data[57466] <= 8'h10 ;
			data[57467] <= 8'h10 ;
			data[57468] <= 8'h10 ;
			data[57469] <= 8'h10 ;
			data[57470] <= 8'h10 ;
			data[57471] <= 8'h10 ;
			data[57472] <= 8'h10 ;
			data[57473] <= 8'h10 ;
			data[57474] <= 8'h10 ;
			data[57475] <= 8'h10 ;
			data[57476] <= 8'h10 ;
			data[57477] <= 8'h10 ;
			data[57478] <= 8'h10 ;
			data[57479] <= 8'h10 ;
			data[57480] <= 8'h10 ;
			data[57481] <= 8'h10 ;
			data[57482] <= 8'h10 ;
			data[57483] <= 8'h10 ;
			data[57484] <= 8'h10 ;
			data[57485] <= 8'h10 ;
			data[57486] <= 8'h10 ;
			data[57487] <= 8'h10 ;
			data[57488] <= 8'h10 ;
			data[57489] <= 8'h10 ;
			data[57490] <= 8'h10 ;
			data[57491] <= 8'h10 ;
			data[57492] <= 8'h10 ;
			data[57493] <= 8'h10 ;
			data[57494] <= 8'h10 ;
			data[57495] <= 8'h10 ;
			data[57496] <= 8'h10 ;
			data[57497] <= 8'h10 ;
			data[57498] <= 8'h10 ;
			data[57499] <= 8'h10 ;
			data[57500] <= 8'h10 ;
			data[57501] <= 8'h10 ;
			data[57502] <= 8'h10 ;
			data[57503] <= 8'h10 ;
			data[57504] <= 8'h10 ;
			data[57505] <= 8'h10 ;
			data[57506] <= 8'h10 ;
			data[57507] <= 8'h10 ;
			data[57508] <= 8'h10 ;
			data[57509] <= 8'h10 ;
			data[57510] <= 8'h10 ;
			data[57511] <= 8'h10 ;
			data[57512] <= 8'h10 ;
			data[57513] <= 8'h10 ;
			data[57514] <= 8'h10 ;
			data[57515] <= 8'h10 ;
			data[57516] <= 8'h10 ;
			data[57517] <= 8'h10 ;
			data[57518] <= 8'h10 ;
			data[57519] <= 8'h10 ;
			data[57520] <= 8'h10 ;
			data[57521] <= 8'h10 ;
			data[57522] <= 8'h10 ;
			data[57523] <= 8'h10 ;
			data[57524] <= 8'h10 ;
			data[57525] <= 8'h10 ;
			data[57526] <= 8'h10 ;
			data[57527] <= 8'h10 ;
			data[57528] <= 8'h10 ;
			data[57529] <= 8'h10 ;
			data[57530] <= 8'h10 ;
			data[57531] <= 8'h10 ;
			data[57532] <= 8'h10 ;
			data[57533] <= 8'h10 ;
			data[57534] <= 8'h10 ;
			data[57535] <= 8'h10 ;
			data[57536] <= 8'h10 ;
			data[57537] <= 8'h10 ;
			data[57538] <= 8'h10 ;
			data[57539] <= 8'h10 ;
			data[57540] <= 8'h10 ;
			data[57541] <= 8'h10 ;
			data[57542] <= 8'h10 ;
			data[57543] <= 8'h10 ;
			data[57544] <= 8'h10 ;
			data[57545] <= 8'h10 ;
			data[57546] <= 8'h10 ;
			data[57547] <= 8'h10 ;
			data[57548] <= 8'h10 ;
			data[57549] <= 8'h10 ;
			data[57550] <= 8'h10 ;
			data[57551] <= 8'h10 ;
			data[57552] <= 8'h10 ;
			data[57553] <= 8'h10 ;
			data[57554] <= 8'h10 ;
			data[57555] <= 8'h10 ;
			data[57556] <= 8'h10 ;
			data[57557] <= 8'h10 ;
			data[57558] <= 8'h10 ;
			data[57559] <= 8'h10 ;
			data[57560] <= 8'h10 ;
			data[57561] <= 8'h10 ;
			data[57562] <= 8'h10 ;
			data[57563] <= 8'h10 ;
			data[57564] <= 8'h10 ;
			data[57565] <= 8'h10 ;
			data[57566] <= 8'h10 ;
			data[57567] <= 8'h10 ;
			data[57568] <= 8'h10 ;
			data[57569] <= 8'h10 ;
			data[57570] <= 8'h10 ;
			data[57571] <= 8'h10 ;
			data[57572] <= 8'h10 ;
			data[57573] <= 8'h10 ;
			data[57574] <= 8'h10 ;
			data[57575] <= 8'h10 ;
			data[57576] <= 8'h10 ;
			data[57577] <= 8'h10 ;
			data[57578] <= 8'h10 ;
			data[57579] <= 8'h10 ;
			data[57580] <= 8'h10 ;
			data[57581] <= 8'h10 ;
			data[57582] <= 8'h10 ;
			data[57583] <= 8'h10 ;
			data[57584] <= 8'h10 ;
			data[57585] <= 8'h10 ;
			data[57586] <= 8'h10 ;
			data[57587] <= 8'h10 ;
			data[57588] <= 8'h10 ;
			data[57589] <= 8'h10 ;
			data[57590] <= 8'h10 ;
			data[57591] <= 8'h10 ;
			data[57592] <= 8'h10 ;
			data[57593] <= 8'h10 ;
			data[57594] <= 8'h10 ;
			data[57595] <= 8'h10 ;
			data[57596] <= 8'h10 ;
			data[57597] <= 8'h10 ;
			data[57598] <= 8'h10 ;
			data[57599] <= 8'h10 ;
			data[57600] <= 8'h10 ;
			data[57601] <= 8'h10 ;
			data[57602] <= 8'h10 ;
			data[57603] <= 8'h10 ;
			data[57604] <= 8'h10 ;
			data[57605] <= 8'h10 ;
			data[57606] <= 8'h10 ;
			data[57607] <= 8'h10 ;
			data[57608] <= 8'h10 ;
			data[57609] <= 8'h10 ;
			data[57610] <= 8'h10 ;
			data[57611] <= 8'h10 ;
			data[57612] <= 8'h10 ;
			data[57613] <= 8'h10 ;
			data[57614] <= 8'h10 ;
			data[57615] <= 8'h10 ;
			data[57616] <= 8'h10 ;
			data[57617] <= 8'h10 ;
			data[57618] <= 8'h10 ;
			data[57619] <= 8'h10 ;
			data[57620] <= 8'h10 ;
			data[57621] <= 8'h10 ;
			data[57622] <= 8'h10 ;
			data[57623] <= 8'h10 ;
			data[57624] <= 8'h10 ;
			data[57625] <= 8'h10 ;
			data[57626] <= 8'h10 ;
			data[57627] <= 8'h10 ;
			data[57628] <= 8'h10 ;
			data[57629] <= 8'h10 ;
			data[57630] <= 8'h10 ;
			data[57631] <= 8'h10 ;
			data[57632] <= 8'h10 ;
			data[57633] <= 8'h10 ;
			data[57634] <= 8'h10 ;
			data[57635] <= 8'h10 ;
			data[57636] <= 8'h10 ;
			data[57637] <= 8'h10 ;
			data[57638] <= 8'h10 ;
			data[57639] <= 8'h10 ;
			data[57640] <= 8'h10 ;
			data[57641] <= 8'h10 ;
			data[57642] <= 8'h10 ;
			data[57643] <= 8'h10 ;
			data[57644] <= 8'h10 ;
			data[57645] <= 8'h10 ;
			data[57646] <= 8'h10 ;
			data[57647] <= 8'h10 ;
			data[57648] <= 8'h10 ;
			data[57649] <= 8'h10 ;
			data[57650] <= 8'h10 ;
			data[57651] <= 8'h10 ;
			data[57652] <= 8'h10 ;
			data[57653] <= 8'h10 ;
			data[57654] <= 8'h10 ;
			data[57655] <= 8'h10 ;
			data[57656] <= 8'h10 ;
			data[57657] <= 8'h10 ;
			data[57658] <= 8'h10 ;
			data[57659] <= 8'h10 ;
			data[57660] <= 8'h10 ;
			data[57661] <= 8'h10 ;
			data[57662] <= 8'h10 ;
			data[57663] <= 8'h10 ;
			data[57664] <= 8'h10 ;
			data[57665] <= 8'h10 ;
			data[57666] <= 8'h10 ;
			data[57667] <= 8'h10 ;
			data[57668] <= 8'h10 ;
			data[57669] <= 8'h10 ;
			data[57670] <= 8'h10 ;
			data[57671] <= 8'h10 ;
			data[57672] <= 8'h10 ;
			data[57673] <= 8'h10 ;
			data[57674] <= 8'h10 ;
			data[57675] <= 8'h10 ;
			data[57676] <= 8'h10 ;
			data[57677] <= 8'h10 ;
			data[57678] <= 8'h10 ;
			data[57679] <= 8'h10 ;
			data[57680] <= 8'h10 ;
			data[57681] <= 8'h10 ;
			data[57682] <= 8'h10 ;
			data[57683] <= 8'h10 ;
			data[57684] <= 8'h10 ;
			data[57685] <= 8'h10 ;
			data[57686] <= 8'h10 ;
			data[57687] <= 8'h10 ;
			data[57688] <= 8'h10 ;
			data[57689] <= 8'h10 ;
			data[57690] <= 8'h10 ;
			data[57691] <= 8'h10 ;
			data[57692] <= 8'h10 ;
			data[57693] <= 8'h10 ;
			data[57694] <= 8'h10 ;
			data[57695] <= 8'h10 ;
			data[57696] <= 8'h10 ;
			data[57697] <= 8'h10 ;
			data[57698] <= 8'h10 ;
			data[57699] <= 8'h10 ;
			data[57700] <= 8'h10 ;
			data[57701] <= 8'h10 ;
			data[57702] <= 8'h10 ;
			data[57703] <= 8'h10 ;
			data[57704] <= 8'h10 ;
			data[57705] <= 8'h10 ;
			data[57706] <= 8'h10 ;
			data[57707] <= 8'h10 ;
			data[57708] <= 8'h10 ;
			data[57709] <= 8'h10 ;
			data[57710] <= 8'h10 ;
			data[57711] <= 8'h10 ;
			data[57712] <= 8'h10 ;
			data[57713] <= 8'h10 ;
			data[57714] <= 8'h10 ;
			data[57715] <= 8'h10 ;
			data[57716] <= 8'h10 ;
			data[57717] <= 8'h10 ;
			data[57718] <= 8'h10 ;
			data[57719] <= 8'h10 ;
			data[57720] <= 8'h10 ;
			data[57721] <= 8'h10 ;
			data[57722] <= 8'h10 ;
			data[57723] <= 8'h10 ;
			data[57724] <= 8'h10 ;
			data[57725] <= 8'h10 ;
			data[57726] <= 8'h10 ;
			data[57727] <= 8'h10 ;
			data[57728] <= 8'h10 ;
			data[57729] <= 8'h10 ;
			data[57730] <= 8'h10 ;
			data[57731] <= 8'h10 ;
			data[57732] <= 8'h10 ;
			data[57733] <= 8'h10 ;
			data[57734] <= 8'h10 ;
			data[57735] <= 8'h10 ;
			data[57736] <= 8'h10 ;
			data[57737] <= 8'h10 ;
			data[57738] <= 8'h10 ;
			data[57739] <= 8'h10 ;
			data[57740] <= 8'h10 ;
			data[57741] <= 8'h10 ;
			data[57742] <= 8'h10 ;
			data[57743] <= 8'h10 ;
			data[57744] <= 8'h10 ;
			data[57745] <= 8'h10 ;
			data[57746] <= 8'h10 ;
			data[57747] <= 8'h10 ;
			data[57748] <= 8'h10 ;
			data[57749] <= 8'h10 ;
			data[57750] <= 8'h10 ;
			data[57751] <= 8'h10 ;
			data[57752] <= 8'h10 ;
			data[57753] <= 8'h10 ;
			data[57754] <= 8'h10 ;
			data[57755] <= 8'h10 ;
			data[57756] <= 8'h10 ;
			data[57757] <= 8'h10 ;
			data[57758] <= 8'h10 ;
			data[57759] <= 8'h10 ;
			data[57760] <= 8'h10 ;
			data[57761] <= 8'h10 ;
			data[57762] <= 8'h10 ;
			data[57763] <= 8'h10 ;
			data[57764] <= 8'h10 ;
			data[57765] <= 8'h10 ;
			data[57766] <= 8'h10 ;
			data[57767] <= 8'h10 ;
			data[57768] <= 8'h10 ;
			data[57769] <= 8'h10 ;
			data[57770] <= 8'h10 ;
			data[57771] <= 8'h10 ;
			data[57772] <= 8'h10 ;
			data[57773] <= 8'h10 ;
			data[57774] <= 8'h10 ;
			data[57775] <= 8'h10 ;
			data[57776] <= 8'h10 ;
			data[57777] <= 8'h10 ;
			data[57778] <= 8'h10 ;
			data[57779] <= 8'h10 ;
			data[57780] <= 8'h10 ;
			data[57781] <= 8'h10 ;
			data[57782] <= 8'h10 ;
			data[57783] <= 8'h10 ;
			data[57784] <= 8'h10 ;
			data[57785] <= 8'h10 ;
			data[57786] <= 8'h10 ;
			data[57787] <= 8'h10 ;
			data[57788] <= 8'h10 ;
			data[57789] <= 8'h10 ;
			data[57790] <= 8'h10 ;
			data[57791] <= 8'h10 ;
			data[57792] <= 8'h10 ;
			data[57793] <= 8'h10 ;
			data[57794] <= 8'h10 ;
			data[57795] <= 8'h10 ;
			data[57796] <= 8'h10 ;
			data[57797] <= 8'h10 ;
			data[57798] <= 8'h10 ;
			data[57799] <= 8'h10 ;
			data[57800] <= 8'h10 ;
			data[57801] <= 8'h10 ;
			data[57802] <= 8'h10 ;
			data[57803] <= 8'h10 ;
			data[57804] <= 8'h10 ;
			data[57805] <= 8'h10 ;
			data[57806] <= 8'h10 ;
			data[57807] <= 8'h10 ;
			data[57808] <= 8'h10 ;
			data[57809] <= 8'h10 ;
			data[57810] <= 8'h10 ;
			data[57811] <= 8'h10 ;
			data[57812] <= 8'h10 ;
			data[57813] <= 8'h10 ;
			data[57814] <= 8'h10 ;
			data[57815] <= 8'h10 ;
			data[57816] <= 8'h10 ;
			data[57817] <= 8'h10 ;
			data[57818] <= 8'h10 ;
			data[57819] <= 8'h10 ;
			data[57820] <= 8'h10 ;
			data[57821] <= 8'h10 ;
			data[57822] <= 8'h10 ;
			data[57823] <= 8'h10 ;
			data[57824] <= 8'h10 ;
			data[57825] <= 8'h10 ;
			data[57826] <= 8'h10 ;
			data[57827] <= 8'h10 ;
			data[57828] <= 8'h10 ;
			data[57829] <= 8'h10 ;
			data[57830] <= 8'h10 ;
			data[57831] <= 8'h10 ;
			data[57832] <= 8'h10 ;
			data[57833] <= 8'h10 ;
			data[57834] <= 8'h10 ;
			data[57835] <= 8'h10 ;
			data[57836] <= 8'h10 ;
			data[57837] <= 8'h10 ;
			data[57838] <= 8'h10 ;
			data[57839] <= 8'h10 ;
			data[57840] <= 8'h10 ;
			data[57841] <= 8'h10 ;
			data[57842] <= 8'h10 ;
			data[57843] <= 8'h10 ;
			data[57844] <= 8'h10 ;
			data[57845] <= 8'h10 ;
			data[57846] <= 8'h10 ;
			data[57847] <= 8'h10 ;
			data[57848] <= 8'h10 ;
			data[57849] <= 8'h10 ;
			data[57850] <= 8'h10 ;
			data[57851] <= 8'h10 ;
			data[57852] <= 8'h10 ;
			data[57853] <= 8'h10 ;
			data[57854] <= 8'h10 ;
			data[57855] <= 8'h10 ;
			data[57856] <= 8'h10 ;
			data[57857] <= 8'h10 ;
			data[57858] <= 8'h10 ;
			data[57859] <= 8'h10 ;
			data[57860] <= 8'h10 ;
			data[57861] <= 8'h10 ;
			data[57862] <= 8'h10 ;
			data[57863] <= 8'h10 ;
			data[57864] <= 8'h10 ;
			data[57865] <= 8'h10 ;
			data[57866] <= 8'h10 ;
			data[57867] <= 8'h10 ;
			data[57868] <= 8'h10 ;
			data[57869] <= 8'h10 ;
			data[57870] <= 8'h10 ;
			data[57871] <= 8'h10 ;
			data[57872] <= 8'h10 ;
			data[57873] <= 8'h10 ;
			data[57874] <= 8'h10 ;
			data[57875] <= 8'h10 ;
			data[57876] <= 8'h10 ;
			data[57877] <= 8'h10 ;
			data[57878] <= 8'h10 ;
			data[57879] <= 8'h10 ;
			data[57880] <= 8'h10 ;
			data[57881] <= 8'h10 ;
			data[57882] <= 8'h10 ;
			data[57883] <= 8'h10 ;
			data[57884] <= 8'h10 ;
			data[57885] <= 8'h10 ;
			data[57886] <= 8'h10 ;
			data[57887] <= 8'h10 ;
			data[57888] <= 8'h10 ;
			data[57889] <= 8'h10 ;
			data[57890] <= 8'h10 ;
			data[57891] <= 8'h10 ;
			data[57892] <= 8'h10 ;
			data[57893] <= 8'h10 ;
			data[57894] <= 8'h10 ;
			data[57895] <= 8'h10 ;
			data[57896] <= 8'h10 ;
			data[57897] <= 8'h10 ;
			data[57898] <= 8'h10 ;
			data[57899] <= 8'h10 ;
			data[57900] <= 8'h10 ;
			data[57901] <= 8'h10 ;
			data[57902] <= 8'h10 ;
			data[57903] <= 8'h10 ;
			data[57904] <= 8'h10 ;
			data[57905] <= 8'h10 ;
			data[57906] <= 8'h10 ;
			data[57907] <= 8'h10 ;
			data[57908] <= 8'h10 ;
			data[57909] <= 8'h10 ;
			data[57910] <= 8'h10 ;
			data[57911] <= 8'h10 ;
			data[57912] <= 8'h10 ;
			data[57913] <= 8'h10 ;
			data[57914] <= 8'h10 ;
			data[57915] <= 8'h10 ;
			data[57916] <= 8'h10 ;
			data[57917] <= 8'h10 ;
			data[57918] <= 8'h10 ;
			data[57919] <= 8'h10 ;
			data[57920] <= 8'h10 ;
			data[57921] <= 8'h10 ;
			data[57922] <= 8'h10 ;
			data[57923] <= 8'h10 ;
			data[57924] <= 8'h10 ;
			data[57925] <= 8'h10 ;
			data[57926] <= 8'h10 ;
			data[57927] <= 8'h10 ;
			data[57928] <= 8'h10 ;
			data[57929] <= 8'h10 ;
			data[57930] <= 8'h10 ;
			data[57931] <= 8'h10 ;
			data[57932] <= 8'h10 ;
			data[57933] <= 8'h10 ;
			data[57934] <= 8'h10 ;
			data[57935] <= 8'h10 ;
			data[57936] <= 8'h10 ;
			data[57937] <= 8'h10 ;
			data[57938] <= 8'h10 ;
			data[57939] <= 8'h10 ;
			data[57940] <= 8'h10 ;
			data[57941] <= 8'h10 ;
			data[57942] <= 8'h10 ;
			data[57943] <= 8'h10 ;
			data[57944] <= 8'h10 ;
			data[57945] <= 8'h10 ;
			data[57946] <= 8'h10 ;
			data[57947] <= 8'h10 ;
			data[57948] <= 8'h10 ;
			data[57949] <= 8'h10 ;
			data[57950] <= 8'h10 ;
			data[57951] <= 8'h10 ;
			data[57952] <= 8'h10 ;
			data[57953] <= 8'h10 ;
			data[57954] <= 8'h10 ;
			data[57955] <= 8'h10 ;
			data[57956] <= 8'h10 ;
			data[57957] <= 8'h10 ;
			data[57958] <= 8'h10 ;
			data[57959] <= 8'h10 ;
			data[57960] <= 8'h10 ;
			data[57961] <= 8'h10 ;
			data[57962] <= 8'h10 ;
			data[57963] <= 8'h10 ;
			data[57964] <= 8'h10 ;
			data[57965] <= 8'h10 ;
			data[57966] <= 8'h10 ;
			data[57967] <= 8'h10 ;
			data[57968] <= 8'h10 ;
			data[57969] <= 8'h10 ;
			data[57970] <= 8'h10 ;
			data[57971] <= 8'h10 ;
			data[57972] <= 8'h10 ;
			data[57973] <= 8'h10 ;
			data[57974] <= 8'h10 ;
			data[57975] <= 8'h10 ;
			data[57976] <= 8'h10 ;
			data[57977] <= 8'h10 ;
			data[57978] <= 8'h10 ;
			data[57979] <= 8'h10 ;
			data[57980] <= 8'h10 ;
			data[57981] <= 8'h10 ;
			data[57982] <= 8'h10 ;
			data[57983] <= 8'h10 ;
			data[57984] <= 8'h10 ;
			data[57985] <= 8'h10 ;
			data[57986] <= 8'h10 ;
			data[57987] <= 8'h10 ;
			data[57988] <= 8'h10 ;
			data[57989] <= 8'h10 ;
			data[57990] <= 8'h10 ;
			data[57991] <= 8'h10 ;
			data[57992] <= 8'h10 ;
			data[57993] <= 8'h10 ;
			data[57994] <= 8'h10 ;
			data[57995] <= 8'h10 ;
			data[57996] <= 8'h10 ;
			data[57997] <= 8'h10 ;
			data[57998] <= 8'h10 ;
			data[57999] <= 8'h10 ;
			data[58000] <= 8'h10 ;
			data[58001] <= 8'h10 ;
			data[58002] <= 8'h10 ;
			data[58003] <= 8'h10 ;
			data[58004] <= 8'h10 ;
			data[58005] <= 8'h10 ;
			data[58006] <= 8'h10 ;
			data[58007] <= 8'h10 ;
			data[58008] <= 8'h10 ;
			data[58009] <= 8'h10 ;
			data[58010] <= 8'h10 ;
			data[58011] <= 8'h10 ;
			data[58012] <= 8'h10 ;
			data[58013] <= 8'h10 ;
			data[58014] <= 8'h10 ;
			data[58015] <= 8'h10 ;
			data[58016] <= 8'h10 ;
			data[58017] <= 8'h10 ;
			data[58018] <= 8'h10 ;
			data[58019] <= 8'h10 ;
			data[58020] <= 8'h10 ;
			data[58021] <= 8'h10 ;
			data[58022] <= 8'h10 ;
			data[58023] <= 8'h10 ;
			data[58024] <= 8'h10 ;
			data[58025] <= 8'h10 ;
			data[58026] <= 8'h10 ;
			data[58027] <= 8'h10 ;
			data[58028] <= 8'h10 ;
			data[58029] <= 8'h10 ;
			data[58030] <= 8'h10 ;
			data[58031] <= 8'h10 ;
			data[58032] <= 8'h10 ;
			data[58033] <= 8'h10 ;
			data[58034] <= 8'h10 ;
			data[58035] <= 8'h10 ;
			data[58036] <= 8'h10 ;
			data[58037] <= 8'h10 ;
			data[58038] <= 8'h10 ;
			data[58039] <= 8'h10 ;
			data[58040] <= 8'h10 ;
			data[58041] <= 8'h10 ;
			data[58042] <= 8'h10 ;
			data[58043] <= 8'h10 ;
			data[58044] <= 8'h10 ;
			data[58045] <= 8'h10 ;
			data[58046] <= 8'h10 ;
			data[58047] <= 8'h10 ;
			data[58048] <= 8'h10 ;
			data[58049] <= 8'h10 ;
			data[58050] <= 8'h10 ;
			data[58051] <= 8'h10 ;
			data[58052] <= 8'h10 ;
			data[58053] <= 8'h10 ;
			data[58054] <= 8'h10 ;
			data[58055] <= 8'h10 ;
			data[58056] <= 8'h10 ;
			data[58057] <= 8'h10 ;
			data[58058] <= 8'h10 ;
			data[58059] <= 8'h10 ;
			data[58060] <= 8'h10 ;
			data[58061] <= 8'h10 ;
			data[58062] <= 8'h10 ;
			data[58063] <= 8'h10 ;
			data[58064] <= 8'h10 ;
			data[58065] <= 8'h10 ;
			data[58066] <= 8'h10 ;
			data[58067] <= 8'h10 ;
			data[58068] <= 8'h10 ;
			data[58069] <= 8'h10 ;
			data[58070] <= 8'h10 ;
			data[58071] <= 8'h10 ;
			data[58072] <= 8'h10 ;
			data[58073] <= 8'h10 ;
			data[58074] <= 8'h10 ;
			data[58075] <= 8'h10 ;
			data[58076] <= 8'h10 ;
			data[58077] <= 8'h10 ;
			data[58078] <= 8'h10 ;
			data[58079] <= 8'h10 ;
			data[58080] <= 8'h10 ;
			data[58081] <= 8'h10 ;
			data[58082] <= 8'h10 ;
			data[58083] <= 8'h10 ;
			data[58084] <= 8'h10 ;
			data[58085] <= 8'h10 ;
			data[58086] <= 8'h10 ;
			data[58087] <= 8'h10 ;
			data[58088] <= 8'h10 ;
			data[58089] <= 8'h10 ;
			data[58090] <= 8'h10 ;
			data[58091] <= 8'h10 ;
			data[58092] <= 8'h10 ;
			data[58093] <= 8'h10 ;
			data[58094] <= 8'h10 ;
			data[58095] <= 8'h10 ;
			data[58096] <= 8'h10 ;
			data[58097] <= 8'h10 ;
			data[58098] <= 8'h10 ;
			data[58099] <= 8'h10 ;
			data[58100] <= 8'h10 ;
			data[58101] <= 8'h10 ;
			data[58102] <= 8'h10 ;
			data[58103] <= 8'h10 ;
			data[58104] <= 8'h10 ;
			data[58105] <= 8'h10 ;
			data[58106] <= 8'h10 ;
			data[58107] <= 8'h10 ;
			data[58108] <= 8'h10 ;
			data[58109] <= 8'h10 ;
			data[58110] <= 8'h10 ;
			data[58111] <= 8'h10 ;
			data[58112] <= 8'h10 ;
			data[58113] <= 8'h10 ;
			data[58114] <= 8'h10 ;
			data[58115] <= 8'h10 ;
			data[58116] <= 8'h10 ;
			data[58117] <= 8'h10 ;
			data[58118] <= 8'h10 ;
			data[58119] <= 8'h10 ;
			data[58120] <= 8'h10 ;
			data[58121] <= 8'h10 ;
			data[58122] <= 8'h10 ;
			data[58123] <= 8'h10 ;
			data[58124] <= 8'h10 ;
			data[58125] <= 8'h10 ;
			data[58126] <= 8'h10 ;
			data[58127] <= 8'h10 ;
			data[58128] <= 8'h10 ;
			data[58129] <= 8'h10 ;
			data[58130] <= 8'h10 ;
			data[58131] <= 8'h10 ;
			data[58132] <= 8'h10 ;
			data[58133] <= 8'h10 ;
			data[58134] <= 8'h10 ;
			data[58135] <= 8'h10 ;
			data[58136] <= 8'h10 ;
			data[58137] <= 8'h10 ;
			data[58138] <= 8'h10 ;
			data[58139] <= 8'h10 ;
			data[58140] <= 8'h10 ;
			data[58141] <= 8'h10 ;
			data[58142] <= 8'h10 ;
			data[58143] <= 8'h10 ;
			data[58144] <= 8'h10 ;
			data[58145] <= 8'h10 ;
			data[58146] <= 8'h10 ;
			data[58147] <= 8'h10 ;
			data[58148] <= 8'h10 ;
			data[58149] <= 8'h10 ;
			data[58150] <= 8'h10 ;
			data[58151] <= 8'h10 ;
			data[58152] <= 8'h10 ;
			data[58153] <= 8'h10 ;
			data[58154] <= 8'h10 ;
			data[58155] <= 8'h10 ;
			data[58156] <= 8'h10 ;
			data[58157] <= 8'h10 ;
			data[58158] <= 8'h10 ;
			data[58159] <= 8'h10 ;
			data[58160] <= 8'h10 ;
			data[58161] <= 8'h10 ;
			data[58162] <= 8'h10 ;
			data[58163] <= 8'h10 ;
			data[58164] <= 8'h10 ;
			data[58165] <= 8'h10 ;
			data[58166] <= 8'h10 ;
			data[58167] <= 8'h10 ;
			data[58168] <= 8'h10 ;
			data[58169] <= 8'h10 ;
			data[58170] <= 8'h10 ;
			data[58171] <= 8'h10 ;
			data[58172] <= 8'h10 ;
			data[58173] <= 8'h10 ;
			data[58174] <= 8'h10 ;
			data[58175] <= 8'h10 ;
			data[58176] <= 8'h10 ;
			data[58177] <= 8'h10 ;
			data[58178] <= 8'h10 ;
			data[58179] <= 8'h10 ;
			data[58180] <= 8'h10 ;
			data[58181] <= 8'h10 ;
			data[58182] <= 8'h10 ;
			data[58183] <= 8'h10 ;
			data[58184] <= 8'h10 ;
			data[58185] <= 8'h10 ;
			data[58186] <= 8'h10 ;
			data[58187] <= 8'h10 ;
			data[58188] <= 8'h10 ;
			data[58189] <= 8'h10 ;
			data[58190] <= 8'h10 ;
			data[58191] <= 8'h10 ;
			data[58192] <= 8'h10 ;
			data[58193] <= 8'h10 ;
			data[58194] <= 8'h10 ;
			data[58195] <= 8'h10 ;
			data[58196] <= 8'h10 ;
			data[58197] <= 8'h10 ;
			data[58198] <= 8'h10 ;
			data[58199] <= 8'h10 ;
			data[58200] <= 8'h10 ;
			data[58201] <= 8'h10 ;
			data[58202] <= 8'h10 ;
			data[58203] <= 8'h10 ;
			data[58204] <= 8'h10 ;
			data[58205] <= 8'h10 ;
			data[58206] <= 8'h10 ;
			data[58207] <= 8'h10 ;
			data[58208] <= 8'h10 ;
			data[58209] <= 8'h10 ;
			data[58210] <= 8'h10 ;
			data[58211] <= 8'h10 ;
			data[58212] <= 8'h10 ;
			data[58213] <= 8'h10 ;
			data[58214] <= 8'h10 ;
			data[58215] <= 8'h10 ;
			data[58216] <= 8'h10 ;
			data[58217] <= 8'h10 ;
			data[58218] <= 8'h10 ;
			data[58219] <= 8'h10 ;
			data[58220] <= 8'h10 ;
			data[58221] <= 8'h10 ;
			data[58222] <= 8'h10 ;
			data[58223] <= 8'h10 ;
			data[58224] <= 8'h10 ;
			data[58225] <= 8'h10 ;
			data[58226] <= 8'h10 ;
			data[58227] <= 8'h10 ;
			data[58228] <= 8'h10 ;
			data[58229] <= 8'h10 ;
			data[58230] <= 8'h10 ;
			data[58231] <= 8'h10 ;
			data[58232] <= 8'h10 ;
			data[58233] <= 8'h10 ;
			data[58234] <= 8'h10 ;
			data[58235] <= 8'h10 ;
			data[58236] <= 8'h10 ;
			data[58237] <= 8'h10 ;
			data[58238] <= 8'h10 ;
			data[58239] <= 8'h10 ;
			data[58240] <= 8'h10 ;
			data[58241] <= 8'h10 ;
			data[58242] <= 8'h10 ;
			data[58243] <= 8'h10 ;
			data[58244] <= 8'h10 ;
			data[58245] <= 8'h10 ;
			data[58246] <= 8'h10 ;
			data[58247] <= 8'h10 ;
			data[58248] <= 8'h10 ;
			data[58249] <= 8'h10 ;
			data[58250] <= 8'h10 ;
			data[58251] <= 8'h10 ;
			data[58252] <= 8'h10 ;
			data[58253] <= 8'h10 ;
			data[58254] <= 8'h10 ;
			data[58255] <= 8'h10 ;
			data[58256] <= 8'h10 ;
			data[58257] <= 8'h10 ;
			data[58258] <= 8'h10 ;
			data[58259] <= 8'h10 ;
			data[58260] <= 8'h10 ;
			data[58261] <= 8'h10 ;
			data[58262] <= 8'h10 ;
			data[58263] <= 8'h10 ;
			data[58264] <= 8'h10 ;
			data[58265] <= 8'h10 ;
			data[58266] <= 8'h10 ;
			data[58267] <= 8'h10 ;
			data[58268] <= 8'h10 ;
			data[58269] <= 8'h10 ;
			data[58270] <= 8'h10 ;
			data[58271] <= 8'h10 ;
			data[58272] <= 8'h10 ;
			data[58273] <= 8'h10 ;
			data[58274] <= 8'h10 ;
			data[58275] <= 8'h10 ;
			data[58276] <= 8'h10 ;
			data[58277] <= 8'h10 ;
			data[58278] <= 8'h10 ;
			data[58279] <= 8'h10 ;
			data[58280] <= 8'h10 ;
			data[58281] <= 8'h10 ;
			data[58282] <= 8'h10 ;
			data[58283] <= 8'h10 ;
			data[58284] <= 8'h10 ;
			data[58285] <= 8'h10 ;
			data[58286] <= 8'h10 ;
			data[58287] <= 8'h10 ;
			data[58288] <= 8'h10 ;
			data[58289] <= 8'h10 ;
			data[58290] <= 8'h10 ;
			data[58291] <= 8'h10 ;
			data[58292] <= 8'h10 ;
			data[58293] <= 8'h10 ;
			data[58294] <= 8'h10 ;
			data[58295] <= 8'h10 ;
			data[58296] <= 8'h10 ;
			data[58297] <= 8'h10 ;
			data[58298] <= 8'h10 ;
			data[58299] <= 8'h10 ;
			data[58300] <= 8'h10 ;
			data[58301] <= 8'h10 ;
			data[58302] <= 8'h10 ;
			data[58303] <= 8'h10 ;
			data[58304] <= 8'h10 ;
			data[58305] <= 8'h10 ;
			data[58306] <= 8'h10 ;
			data[58307] <= 8'h10 ;
			data[58308] <= 8'h10 ;
			data[58309] <= 8'h10 ;
			data[58310] <= 8'h10 ;
			data[58311] <= 8'h10 ;
			data[58312] <= 8'h10 ;
			data[58313] <= 8'h10 ;
			data[58314] <= 8'h10 ;
			data[58315] <= 8'h10 ;
			data[58316] <= 8'h10 ;
			data[58317] <= 8'h10 ;
			data[58318] <= 8'h10 ;
			data[58319] <= 8'h10 ;
			data[58320] <= 8'h10 ;
			data[58321] <= 8'h10 ;
			data[58322] <= 8'h10 ;
			data[58323] <= 8'h10 ;
			data[58324] <= 8'h10 ;
			data[58325] <= 8'h10 ;
			data[58326] <= 8'h10 ;
			data[58327] <= 8'h10 ;
			data[58328] <= 8'h10 ;
			data[58329] <= 8'h10 ;
			data[58330] <= 8'h10 ;
			data[58331] <= 8'h10 ;
			data[58332] <= 8'h10 ;
			data[58333] <= 8'h10 ;
			data[58334] <= 8'h10 ;
			data[58335] <= 8'h10 ;
			data[58336] <= 8'h10 ;
			data[58337] <= 8'h10 ;
			data[58338] <= 8'h10 ;
			data[58339] <= 8'h10 ;
			data[58340] <= 8'h10 ;
			data[58341] <= 8'h10 ;
			data[58342] <= 8'h10 ;
			data[58343] <= 8'h10 ;
			data[58344] <= 8'h10 ;
			data[58345] <= 8'h10 ;
			data[58346] <= 8'h10 ;
			data[58347] <= 8'h10 ;
			data[58348] <= 8'h10 ;
			data[58349] <= 8'h10 ;
			data[58350] <= 8'h10 ;
			data[58351] <= 8'h10 ;
			data[58352] <= 8'h10 ;
			data[58353] <= 8'h10 ;
			data[58354] <= 8'h10 ;
			data[58355] <= 8'h10 ;
			data[58356] <= 8'h10 ;
			data[58357] <= 8'h10 ;
			data[58358] <= 8'h10 ;
			data[58359] <= 8'h10 ;
			data[58360] <= 8'h10 ;
			data[58361] <= 8'h10 ;
			data[58362] <= 8'h10 ;
			data[58363] <= 8'h10 ;
			data[58364] <= 8'h10 ;
			data[58365] <= 8'h10 ;
			data[58366] <= 8'h10 ;
			data[58367] <= 8'h10 ;
			data[58368] <= 8'h10 ;
			data[58369] <= 8'h10 ;
			data[58370] <= 8'h10 ;
			data[58371] <= 8'h10 ;
			data[58372] <= 8'h10 ;
			data[58373] <= 8'h10 ;
			data[58374] <= 8'h10 ;
			data[58375] <= 8'h10 ;
			data[58376] <= 8'h10 ;
			data[58377] <= 8'h10 ;
			data[58378] <= 8'h10 ;
			data[58379] <= 8'h10 ;
			data[58380] <= 8'h10 ;
			data[58381] <= 8'h10 ;
			data[58382] <= 8'h10 ;
			data[58383] <= 8'h10 ;
			data[58384] <= 8'h10 ;
			data[58385] <= 8'h10 ;
			data[58386] <= 8'h10 ;
			data[58387] <= 8'h10 ;
			data[58388] <= 8'h10 ;
			data[58389] <= 8'h10 ;
			data[58390] <= 8'h10 ;
			data[58391] <= 8'h10 ;
			data[58392] <= 8'h10 ;
			data[58393] <= 8'h10 ;
			data[58394] <= 8'h10 ;
			data[58395] <= 8'h10 ;
			data[58396] <= 8'h10 ;
			data[58397] <= 8'h10 ;
			data[58398] <= 8'h10 ;
			data[58399] <= 8'h10 ;
			data[58400] <= 8'h10 ;
			data[58401] <= 8'h10 ;
			data[58402] <= 8'h10 ;
			data[58403] <= 8'h10 ;
			data[58404] <= 8'h10 ;
			data[58405] <= 8'h10 ;
			data[58406] <= 8'h10 ;
			data[58407] <= 8'h10 ;
			data[58408] <= 8'h10 ;
			data[58409] <= 8'h10 ;
			data[58410] <= 8'h10 ;
			data[58411] <= 8'h10 ;
			data[58412] <= 8'h10 ;
			data[58413] <= 8'h10 ;
			data[58414] <= 8'h10 ;
			data[58415] <= 8'h10 ;
			data[58416] <= 8'h10 ;
			data[58417] <= 8'h10 ;
			data[58418] <= 8'h10 ;
			data[58419] <= 8'h10 ;
			data[58420] <= 8'h10 ;
			data[58421] <= 8'h10 ;
			data[58422] <= 8'h10 ;
			data[58423] <= 8'h10 ;
			data[58424] <= 8'h10 ;
			data[58425] <= 8'h10 ;
			data[58426] <= 8'h10 ;
			data[58427] <= 8'h10 ;
			data[58428] <= 8'h10 ;
			data[58429] <= 8'h10 ;
			data[58430] <= 8'h10 ;
			data[58431] <= 8'h10 ;
			data[58432] <= 8'h10 ;
			data[58433] <= 8'h10 ;
			data[58434] <= 8'h10 ;
			data[58435] <= 8'h10 ;
			data[58436] <= 8'h10 ;
			data[58437] <= 8'h10 ;
			data[58438] <= 8'h10 ;
			data[58439] <= 8'h10 ;
			data[58440] <= 8'h10 ;
			data[58441] <= 8'h10 ;
			data[58442] <= 8'h10 ;
			data[58443] <= 8'h10 ;
			data[58444] <= 8'h10 ;
			data[58445] <= 8'h10 ;
			data[58446] <= 8'h10 ;
			data[58447] <= 8'h10 ;
			data[58448] <= 8'h10 ;
			data[58449] <= 8'h10 ;
			data[58450] <= 8'h10 ;
			data[58451] <= 8'h10 ;
			data[58452] <= 8'h10 ;
			data[58453] <= 8'h10 ;
			data[58454] <= 8'h10 ;
			data[58455] <= 8'h10 ;
			data[58456] <= 8'h10 ;
			data[58457] <= 8'h10 ;
			data[58458] <= 8'h10 ;
			data[58459] <= 8'h10 ;
			data[58460] <= 8'h10 ;
			data[58461] <= 8'h10 ;
			data[58462] <= 8'h10 ;
			data[58463] <= 8'h10 ;
			data[58464] <= 8'h10 ;
			data[58465] <= 8'h10 ;
			data[58466] <= 8'h10 ;
			data[58467] <= 8'h10 ;
			data[58468] <= 8'h10 ;
			data[58469] <= 8'h10 ;
			data[58470] <= 8'h10 ;
			data[58471] <= 8'h10 ;
			data[58472] <= 8'h10 ;
			data[58473] <= 8'h10 ;
			data[58474] <= 8'h10 ;
			data[58475] <= 8'h10 ;
			data[58476] <= 8'h10 ;
			data[58477] <= 8'h10 ;
			data[58478] <= 8'h10 ;
			data[58479] <= 8'h10 ;
			data[58480] <= 8'h10 ;
			data[58481] <= 8'h10 ;
			data[58482] <= 8'h10 ;
			data[58483] <= 8'h10 ;
			data[58484] <= 8'h10 ;
			data[58485] <= 8'h10 ;
			data[58486] <= 8'h10 ;
			data[58487] <= 8'h10 ;
			data[58488] <= 8'h10 ;
			data[58489] <= 8'h10 ;
			data[58490] <= 8'h10 ;
			data[58491] <= 8'h10 ;
			data[58492] <= 8'h10 ;
			data[58493] <= 8'h10 ;
			data[58494] <= 8'h10 ;
			data[58495] <= 8'h10 ;
			data[58496] <= 8'h10 ;
			data[58497] <= 8'h10 ;
			data[58498] <= 8'h10 ;
			data[58499] <= 8'h10 ;
			data[58500] <= 8'h10 ;
			data[58501] <= 8'h10 ;
			data[58502] <= 8'h10 ;
			data[58503] <= 8'h10 ;
			data[58504] <= 8'h10 ;
			data[58505] <= 8'h10 ;
			data[58506] <= 8'h10 ;
			data[58507] <= 8'h10 ;
			data[58508] <= 8'h10 ;
			data[58509] <= 8'h10 ;
			data[58510] <= 8'h10 ;
			data[58511] <= 8'h10 ;
			data[58512] <= 8'h10 ;
			data[58513] <= 8'h10 ;
			data[58514] <= 8'h10 ;
			data[58515] <= 8'h10 ;
			data[58516] <= 8'h10 ;
			data[58517] <= 8'h10 ;
			data[58518] <= 8'h10 ;
			data[58519] <= 8'h10 ;
			data[58520] <= 8'h10 ;
			data[58521] <= 8'h10 ;
			data[58522] <= 8'h10 ;
			data[58523] <= 8'h10 ;
			data[58524] <= 8'h10 ;
			data[58525] <= 8'h10 ;
			data[58526] <= 8'h10 ;
			data[58527] <= 8'h10 ;
			data[58528] <= 8'h10 ;
			data[58529] <= 8'h10 ;
			data[58530] <= 8'h10 ;
			data[58531] <= 8'h10 ;
			data[58532] <= 8'h10 ;
			data[58533] <= 8'h10 ;
			data[58534] <= 8'h10 ;
			data[58535] <= 8'h10 ;
			data[58536] <= 8'h10 ;
			data[58537] <= 8'h10 ;
			data[58538] <= 8'h10 ;
			data[58539] <= 8'h10 ;
			data[58540] <= 8'h10 ;
			data[58541] <= 8'h10 ;
			data[58542] <= 8'h10 ;
			data[58543] <= 8'h10 ;
			data[58544] <= 8'h10 ;
			data[58545] <= 8'h10 ;
			data[58546] <= 8'h10 ;
			data[58547] <= 8'h10 ;
			data[58548] <= 8'h10 ;
			data[58549] <= 8'h10 ;
			data[58550] <= 8'h10 ;
			data[58551] <= 8'h10 ;
			data[58552] <= 8'h10 ;
			data[58553] <= 8'h10 ;
			data[58554] <= 8'h10 ;
			data[58555] <= 8'h10 ;
			data[58556] <= 8'h10 ;
			data[58557] <= 8'h10 ;
			data[58558] <= 8'h10 ;
			data[58559] <= 8'h10 ;
			data[58560] <= 8'h10 ;
			data[58561] <= 8'h10 ;
			data[58562] <= 8'h10 ;
			data[58563] <= 8'h10 ;
			data[58564] <= 8'h10 ;
			data[58565] <= 8'h10 ;
			data[58566] <= 8'h10 ;
			data[58567] <= 8'h10 ;
			data[58568] <= 8'h10 ;
			data[58569] <= 8'h10 ;
			data[58570] <= 8'h10 ;
			data[58571] <= 8'h10 ;
			data[58572] <= 8'h10 ;
			data[58573] <= 8'h10 ;
			data[58574] <= 8'h10 ;
			data[58575] <= 8'h10 ;
			data[58576] <= 8'h10 ;
			data[58577] <= 8'h10 ;
			data[58578] <= 8'h10 ;
			data[58579] <= 8'h10 ;
			data[58580] <= 8'h10 ;
			data[58581] <= 8'h10 ;
			data[58582] <= 8'h10 ;
			data[58583] <= 8'h10 ;
			data[58584] <= 8'h10 ;
			data[58585] <= 8'h10 ;
			data[58586] <= 8'h10 ;
			data[58587] <= 8'h10 ;
			data[58588] <= 8'h10 ;
			data[58589] <= 8'h10 ;
			data[58590] <= 8'h10 ;
			data[58591] <= 8'h10 ;
			data[58592] <= 8'h10 ;
			data[58593] <= 8'h10 ;
			data[58594] <= 8'h10 ;
			data[58595] <= 8'h10 ;
			data[58596] <= 8'h10 ;
			data[58597] <= 8'h10 ;
			data[58598] <= 8'h10 ;
			data[58599] <= 8'h10 ;
			data[58600] <= 8'h10 ;
			data[58601] <= 8'h10 ;
			data[58602] <= 8'h10 ;
			data[58603] <= 8'h10 ;
			data[58604] <= 8'h10 ;
			data[58605] <= 8'h10 ;
			data[58606] <= 8'h10 ;
			data[58607] <= 8'h10 ;
			data[58608] <= 8'h10 ;
			data[58609] <= 8'h10 ;
			data[58610] <= 8'h10 ;
			data[58611] <= 8'h10 ;
			data[58612] <= 8'h10 ;
			data[58613] <= 8'h10 ;
			data[58614] <= 8'h10 ;
			data[58615] <= 8'h10 ;
			data[58616] <= 8'h10 ;
			data[58617] <= 8'h10 ;
			data[58618] <= 8'h10 ;
			data[58619] <= 8'h10 ;
			data[58620] <= 8'h10 ;
			data[58621] <= 8'h10 ;
			data[58622] <= 8'h10 ;
			data[58623] <= 8'h10 ;
			data[58624] <= 8'h10 ;
			data[58625] <= 8'h10 ;
			data[58626] <= 8'h10 ;
			data[58627] <= 8'h10 ;
			data[58628] <= 8'h10 ;
			data[58629] <= 8'h10 ;
			data[58630] <= 8'h10 ;
			data[58631] <= 8'h10 ;
			data[58632] <= 8'h10 ;
			data[58633] <= 8'h10 ;
			data[58634] <= 8'h10 ;
			data[58635] <= 8'h10 ;
			data[58636] <= 8'h10 ;
			data[58637] <= 8'h10 ;
			data[58638] <= 8'h10 ;
			data[58639] <= 8'h10 ;
			data[58640] <= 8'h10 ;
			data[58641] <= 8'h10 ;
			data[58642] <= 8'h10 ;
			data[58643] <= 8'h10 ;
			data[58644] <= 8'h10 ;
			data[58645] <= 8'h10 ;
			data[58646] <= 8'h10 ;
			data[58647] <= 8'h10 ;
			data[58648] <= 8'h10 ;
			data[58649] <= 8'h10 ;
			data[58650] <= 8'h10 ;
			data[58651] <= 8'h10 ;
			data[58652] <= 8'h10 ;
			data[58653] <= 8'h10 ;
			data[58654] <= 8'h10 ;
			data[58655] <= 8'h10 ;
			data[58656] <= 8'h10 ;
			data[58657] <= 8'h10 ;
			data[58658] <= 8'h10 ;
			data[58659] <= 8'h10 ;
			data[58660] <= 8'h10 ;
			data[58661] <= 8'h10 ;
			data[58662] <= 8'h10 ;
			data[58663] <= 8'h10 ;
			data[58664] <= 8'h10 ;
			data[58665] <= 8'h10 ;
			data[58666] <= 8'h10 ;
			data[58667] <= 8'h10 ;
			data[58668] <= 8'h10 ;
			data[58669] <= 8'h10 ;
			data[58670] <= 8'h10 ;
			data[58671] <= 8'h10 ;
			data[58672] <= 8'h10 ;
			data[58673] <= 8'h10 ;
			data[58674] <= 8'h10 ;
			data[58675] <= 8'h10 ;
			data[58676] <= 8'h10 ;
			data[58677] <= 8'h10 ;
			data[58678] <= 8'h10 ;
			data[58679] <= 8'h10 ;
			data[58680] <= 8'h10 ;
			data[58681] <= 8'h10 ;
			data[58682] <= 8'h10 ;
			data[58683] <= 8'h10 ;
			data[58684] <= 8'h10 ;
			data[58685] <= 8'h10 ;
			data[58686] <= 8'h10 ;
			data[58687] <= 8'h10 ;
			data[58688] <= 8'h10 ;
			data[58689] <= 8'h10 ;
			data[58690] <= 8'h10 ;
			data[58691] <= 8'h10 ;
			data[58692] <= 8'h10 ;
			data[58693] <= 8'h10 ;
			data[58694] <= 8'h10 ;
			data[58695] <= 8'h10 ;
			data[58696] <= 8'h10 ;
			data[58697] <= 8'h10 ;
			data[58698] <= 8'h10 ;
			data[58699] <= 8'h10 ;
			data[58700] <= 8'h10 ;
			data[58701] <= 8'h10 ;
			data[58702] <= 8'h10 ;
			data[58703] <= 8'h10 ;
			data[58704] <= 8'h10 ;
			data[58705] <= 8'h10 ;
			data[58706] <= 8'h10 ;
			data[58707] <= 8'h10 ;
			data[58708] <= 8'h10 ;
			data[58709] <= 8'h10 ;
			data[58710] <= 8'h10 ;
			data[58711] <= 8'h10 ;
			data[58712] <= 8'h10 ;
			data[58713] <= 8'h10 ;
			data[58714] <= 8'h10 ;
			data[58715] <= 8'h10 ;
			data[58716] <= 8'h10 ;
			data[58717] <= 8'h10 ;
			data[58718] <= 8'h10 ;
			data[58719] <= 8'h10 ;
			data[58720] <= 8'h10 ;
			data[58721] <= 8'h10 ;
			data[58722] <= 8'h10 ;
			data[58723] <= 8'h10 ;
			data[58724] <= 8'h10 ;
			data[58725] <= 8'h10 ;
			data[58726] <= 8'h10 ;
			data[58727] <= 8'h10 ;
			data[58728] <= 8'h10 ;
			data[58729] <= 8'h10 ;
			data[58730] <= 8'h10 ;
			data[58731] <= 8'h10 ;
			data[58732] <= 8'h10 ;
			data[58733] <= 8'h10 ;
			data[58734] <= 8'h10 ;
			data[58735] <= 8'h10 ;
			data[58736] <= 8'h10 ;
			data[58737] <= 8'h10 ;
			data[58738] <= 8'h10 ;
			data[58739] <= 8'h10 ;
			data[58740] <= 8'h10 ;
			data[58741] <= 8'h10 ;
			data[58742] <= 8'h10 ;
			data[58743] <= 8'h10 ;
			data[58744] <= 8'h10 ;
			data[58745] <= 8'h10 ;
			data[58746] <= 8'h10 ;
			data[58747] <= 8'h10 ;
			data[58748] <= 8'h10 ;
			data[58749] <= 8'h10 ;
			data[58750] <= 8'h10 ;
			data[58751] <= 8'h10 ;
			data[58752] <= 8'h10 ;
			data[58753] <= 8'h10 ;
			data[58754] <= 8'h10 ;
			data[58755] <= 8'h10 ;
			data[58756] <= 8'h10 ;
			data[58757] <= 8'h10 ;
			data[58758] <= 8'h10 ;
			data[58759] <= 8'h10 ;
			data[58760] <= 8'h10 ;
			data[58761] <= 8'h10 ;
			data[58762] <= 8'h10 ;
			data[58763] <= 8'h10 ;
			data[58764] <= 8'h10 ;
			data[58765] <= 8'h10 ;
			data[58766] <= 8'h10 ;
			data[58767] <= 8'h10 ;
			data[58768] <= 8'h10 ;
			data[58769] <= 8'h10 ;
			data[58770] <= 8'h10 ;
			data[58771] <= 8'h10 ;
			data[58772] <= 8'h10 ;
			data[58773] <= 8'h10 ;
			data[58774] <= 8'h10 ;
			data[58775] <= 8'h10 ;
			data[58776] <= 8'h10 ;
			data[58777] <= 8'h10 ;
			data[58778] <= 8'h10 ;
			data[58779] <= 8'h10 ;
			data[58780] <= 8'h10 ;
			data[58781] <= 8'h10 ;
			data[58782] <= 8'h10 ;
			data[58783] <= 8'h10 ;
			data[58784] <= 8'h10 ;
			data[58785] <= 8'h10 ;
			data[58786] <= 8'h10 ;
			data[58787] <= 8'h10 ;
			data[58788] <= 8'h10 ;
			data[58789] <= 8'h10 ;
			data[58790] <= 8'h10 ;
			data[58791] <= 8'h10 ;
			data[58792] <= 8'h10 ;
			data[58793] <= 8'h10 ;
			data[58794] <= 8'h10 ;
			data[58795] <= 8'h10 ;
			data[58796] <= 8'h10 ;
			data[58797] <= 8'h10 ;
			data[58798] <= 8'h10 ;
			data[58799] <= 8'h10 ;
			data[58800] <= 8'h10 ;
			data[58801] <= 8'h10 ;
			data[58802] <= 8'h10 ;
			data[58803] <= 8'h10 ;
			data[58804] <= 8'h10 ;
			data[58805] <= 8'h10 ;
			data[58806] <= 8'h10 ;
			data[58807] <= 8'h10 ;
			data[58808] <= 8'h10 ;
			data[58809] <= 8'h10 ;
			data[58810] <= 8'h10 ;
			data[58811] <= 8'h10 ;
			data[58812] <= 8'h10 ;
			data[58813] <= 8'h10 ;
			data[58814] <= 8'h10 ;
			data[58815] <= 8'h10 ;
			data[58816] <= 8'h10 ;
			data[58817] <= 8'h10 ;
			data[58818] <= 8'h10 ;
			data[58819] <= 8'h10 ;
			data[58820] <= 8'h10 ;
			data[58821] <= 8'h10 ;
			data[58822] <= 8'h10 ;
			data[58823] <= 8'h10 ;
			data[58824] <= 8'h10 ;
			data[58825] <= 8'h10 ;
			data[58826] <= 8'h10 ;
			data[58827] <= 8'h10 ;
			data[58828] <= 8'h10 ;
			data[58829] <= 8'h10 ;
			data[58830] <= 8'h10 ;
			data[58831] <= 8'h10 ;
			data[58832] <= 8'h10 ;
			data[58833] <= 8'h10 ;
			data[58834] <= 8'h10 ;
			data[58835] <= 8'h10 ;
			data[58836] <= 8'h10 ;
			data[58837] <= 8'h10 ;
			data[58838] <= 8'h10 ;
			data[58839] <= 8'h10 ;
			data[58840] <= 8'h10 ;
			data[58841] <= 8'h10 ;
			data[58842] <= 8'h10 ;
			data[58843] <= 8'h10 ;
			data[58844] <= 8'h10 ;
			data[58845] <= 8'h10 ;
			data[58846] <= 8'h10 ;
			data[58847] <= 8'h10 ;
			data[58848] <= 8'h10 ;
			data[58849] <= 8'h10 ;
			data[58850] <= 8'h10 ;
			data[58851] <= 8'h10 ;
			data[58852] <= 8'h10 ;
			data[58853] <= 8'h10 ;
			data[58854] <= 8'h10 ;
			data[58855] <= 8'h10 ;
			data[58856] <= 8'h10 ;
			data[58857] <= 8'h10 ;
			data[58858] <= 8'h10 ;
			data[58859] <= 8'h10 ;
			data[58860] <= 8'h10 ;
			data[58861] <= 8'h10 ;
			data[58862] <= 8'h10 ;
			data[58863] <= 8'h10 ;
			data[58864] <= 8'h10 ;
			data[58865] <= 8'h10 ;
			data[58866] <= 8'h10 ;
			data[58867] <= 8'h10 ;
			data[58868] <= 8'h10 ;
			data[58869] <= 8'h10 ;
			data[58870] <= 8'h10 ;
			data[58871] <= 8'h10 ;
			data[58872] <= 8'h10 ;
			data[58873] <= 8'h10 ;
			data[58874] <= 8'h10 ;
			data[58875] <= 8'h10 ;
			data[58876] <= 8'h10 ;
			data[58877] <= 8'h10 ;
			data[58878] <= 8'h10 ;
			data[58879] <= 8'h10 ;
			data[58880] <= 8'h10 ;
			data[58881] <= 8'h10 ;
			data[58882] <= 8'h10 ;
			data[58883] <= 8'h10 ;
			data[58884] <= 8'h10 ;
			data[58885] <= 8'h10 ;
			data[58886] <= 8'h10 ;
			data[58887] <= 8'h10 ;
			data[58888] <= 8'h10 ;
			data[58889] <= 8'h10 ;
			data[58890] <= 8'h10 ;
			data[58891] <= 8'h10 ;
			data[58892] <= 8'h10 ;
			data[58893] <= 8'h10 ;
			data[58894] <= 8'h10 ;
			data[58895] <= 8'h10 ;
			data[58896] <= 8'h10 ;
			data[58897] <= 8'h10 ;
			data[58898] <= 8'h10 ;
			data[58899] <= 8'h10 ;
			data[58900] <= 8'h10 ;
			data[58901] <= 8'h10 ;
			data[58902] <= 8'h10 ;
			data[58903] <= 8'h10 ;
			data[58904] <= 8'h10 ;
			data[58905] <= 8'h10 ;
			data[58906] <= 8'h10 ;
			data[58907] <= 8'h10 ;
			data[58908] <= 8'h10 ;
			data[58909] <= 8'h10 ;
			data[58910] <= 8'h10 ;
			data[58911] <= 8'h10 ;
			data[58912] <= 8'h10 ;
			data[58913] <= 8'h10 ;
			data[58914] <= 8'h10 ;
			data[58915] <= 8'h10 ;
			data[58916] <= 8'h10 ;
			data[58917] <= 8'h10 ;
			data[58918] <= 8'h10 ;
			data[58919] <= 8'h10 ;
			data[58920] <= 8'h10 ;
			data[58921] <= 8'h10 ;
			data[58922] <= 8'h10 ;
			data[58923] <= 8'h10 ;
			data[58924] <= 8'h10 ;
			data[58925] <= 8'h10 ;
			data[58926] <= 8'h10 ;
			data[58927] <= 8'h10 ;
			data[58928] <= 8'h10 ;
			data[58929] <= 8'h10 ;
			data[58930] <= 8'h10 ;
			data[58931] <= 8'h10 ;
			data[58932] <= 8'h10 ;
			data[58933] <= 8'h10 ;
			data[58934] <= 8'h10 ;
			data[58935] <= 8'h10 ;
			data[58936] <= 8'h10 ;
			data[58937] <= 8'h10 ;
			data[58938] <= 8'h10 ;
			data[58939] <= 8'h10 ;
			data[58940] <= 8'h10 ;
			data[58941] <= 8'h10 ;
			data[58942] <= 8'h10 ;
			data[58943] <= 8'h10 ;
			data[58944] <= 8'h10 ;
			data[58945] <= 8'h10 ;
			data[58946] <= 8'h10 ;
			data[58947] <= 8'h10 ;
			data[58948] <= 8'h10 ;
			data[58949] <= 8'h10 ;
			data[58950] <= 8'h10 ;
			data[58951] <= 8'h10 ;
			data[58952] <= 8'h10 ;
			data[58953] <= 8'h10 ;
			data[58954] <= 8'h10 ;
			data[58955] <= 8'h10 ;
			data[58956] <= 8'h10 ;
			data[58957] <= 8'h10 ;
			data[58958] <= 8'h10 ;
			data[58959] <= 8'h10 ;
			data[58960] <= 8'h10 ;
			data[58961] <= 8'h10 ;
			data[58962] <= 8'h10 ;
			data[58963] <= 8'h10 ;
			data[58964] <= 8'h10 ;
			data[58965] <= 8'h10 ;
			data[58966] <= 8'h10 ;
			data[58967] <= 8'h10 ;
			data[58968] <= 8'h10 ;
			data[58969] <= 8'h10 ;
			data[58970] <= 8'h10 ;
			data[58971] <= 8'h10 ;
			data[58972] <= 8'h10 ;
			data[58973] <= 8'h10 ;
			data[58974] <= 8'h10 ;
			data[58975] <= 8'h10 ;
			data[58976] <= 8'h10 ;
			data[58977] <= 8'h10 ;
			data[58978] <= 8'h10 ;
			data[58979] <= 8'h10 ;
			data[58980] <= 8'h10 ;
			data[58981] <= 8'h10 ;
			data[58982] <= 8'h10 ;
			data[58983] <= 8'h10 ;
			data[58984] <= 8'h10 ;
			data[58985] <= 8'h10 ;
			data[58986] <= 8'h10 ;
			data[58987] <= 8'h10 ;
			data[58988] <= 8'h10 ;
			data[58989] <= 8'h10 ;
			data[58990] <= 8'h10 ;
			data[58991] <= 8'h10 ;
			data[58992] <= 8'h10 ;
			data[58993] <= 8'h10 ;
			data[58994] <= 8'h10 ;
			data[58995] <= 8'h10 ;
			data[58996] <= 8'h10 ;
			data[58997] <= 8'h10 ;
			data[58998] <= 8'h10 ;
			data[58999] <= 8'h10 ;
			data[59000] <= 8'h10 ;
			data[59001] <= 8'h10 ;
			data[59002] <= 8'h10 ;
			data[59003] <= 8'h10 ;
			data[59004] <= 8'h10 ;
			data[59005] <= 8'h10 ;
			data[59006] <= 8'h10 ;
			data[59007] <= 8'h10 ;
			data[59008] <= 8'h10 ;
			data[59009] <= 8'h10 ;
			data[59010] <= 8'h10 ;
			data[59011] <= 8'h10 ;
			data[59012] <= 8'h10 ;
			data[59013] <= 8'h10 ;
			data[59014] <= 8'h10 ;
			data[59015] <= 8'h10 ;
			data[59016] <= 8'h10 ;
			data[59017] <= 8'h10 ;
			data[59018] <= 8'h10 ;
			data[59019] <= 8'h10 ;
			data[59020] <= 8'h10 ;
			data[59021] <= 8'h10 ;
			data[59022] <= 8'h10 ;
			data[59023] <= 8'h10 ;
			data[59024] <= 8'h10 ;
			data[59025] <= 8'h10 ;
			data[59026] <= 8'h10 ;
			data[59027] <= 8'h10 ;
			data[59028] <= 8'h10 ;
			data[59029] <= 8'h10 ;
			data[59030] <= 8'h10 ;
			data[59031] <= 8'h10 ;
			data[59032] <= 8'h10 ;
			data[59033] <= 8'h10 ;
			data[59034] <= 8'h10 ;
			data[59035] <= 8'h10 ;
			data[59036] <= 8'h10 ;
			data[59037] <= 8'h10 ;
			data[59038] <= 8'h10 ;
			data[59039] <= 8'h10 ;
			data[59040] <= 8'h10 ;
			data[59041] <= 8'h10 ;
			data[59042] <= 8'h10 ;
			data[59043] <= 8'h10 ;
			data[59044] <= 8'h10 ;
			data[59045] <= 8'h10 ;
			data[59046] <= 8'h10 ;
			data[59047] <= 8'h10 ;
			data[59048] <= 8'h10 ;
			data[59049] <= 8'h10 ;
			data[59050] <= 8'h10 ;
			data[59051] <= 8'h10 ;
			data[59052] <= 8'h10 ;
			data[59053] <= 8'h10 ;
			data[59054] <= 8'h10 ;
			data[59055] <= 8'h10 ;
			data[59056] <= 8'h10 ;
			data[59057] <= 8'h10 ;
			data[59058] <= 8'h10 ;
			data[59059] <= 8'h10 ;
			data[59060] <= 8'h10 ;
			data[59061] <= 8'h10 ;
			data[59062] <= 8'h10 ;
			data[59063] <= 8'h10 ;
			data[59064] <= 8'h10 ;
			data[59065] <= 8'h10 ;
			data[59066] <= 8'h10 ;
			data[59067] <= 8'h10 ;
			data[59068] <= 8'h10 ;
			data[59069] <= 8'h10 ;
			data[59070] <= 8'h10 ;
			data[59071] <= 8'h10 ;
			data[59072] <= 8'h10 ;
			data[59073] <= 8'h10 ;
			data[59074] <= 8'h10 ;
			data[59075] <= 8'h10 ;
			data[59076] <= 8'h10 ;
			data[59077] <= 8'h10 ;
			data[59078] <= 8'h10 ;
			data[59079] <= 8'h10 ;
			data[59080] <= 8'h10 ;
			data[59081] <= 8'h10 ;
			data[59082] <= 8'h10 ;
			data[59083] <= 8'h10 ;
			data[59084] <= 8'h10 ;
			data[59085] <= 8'h10 ;
			data[59086] <= 8'h10 ;
			data[59087] <= 8'h10 ;
			data[59088] <= 8'h10 ;
			data[59089] <= 8'h10 ;
			data[59090] <= 8'h10 ;
			data[59091] <= 8'h10 ;
			data[59092] <= 8'h10 ;
			data[59093] <= 8'h10 ;
			data[59094] <= 8'h10 ;
			data[59095] <= 8'h10 ;
			data[59096] <= 8'h10 ;
			data[59097] <= 8'h10 ;
			data[59098] <= 8'h10 ;
			data[59099] <= 8'h10 ;
			data[59100] <= 8'h10 ;
			data[59101] <= 8'h10 ;
			data[59102] <= 8'h10 ;
			data[59103] <= 8'h10 ;
			data[59104] <= 8'h10 ;
			data[59105] <= 8'h10 ;
			data[59106] <= 8'h10 ;
			data[59107] <= 8'h10 ;
			data[59108] <= 8'h10 ;
			data[59109] <= 8'h10 ;
			data[59110] <= 8'h10 ;
			data[59111] <= 8'h10 ;
			data[59112] <= 8'h10 ;
			data[59113] <= 8'h10 ;
			data[59114] <= 8'h10 ;
			data[59115] <= 8'h10 ;
			data[59116] <= 8'h10 ;
			data[59117] <= 8'h10 ;
			data[59118] <= 8'h10 ;
			data[59119] <= 8'h10 ;
			data[59120] <= 8'h10 ;
			data[59121] <= 8'h10 ;
			data[59122] <= 8'h10 ;
			data[59123] <= 8'h10 ;
			data[59124] <= 8'h10 ;
			data[59125] <= 8'h10 ;
			data[59126] <= 8'h10 ;
			data[59127] <= 8'h10 ;
			data[59128] <= 8'h10 ;
			data[59129] <= 8'h10 ;
			data[59130] <= 8'h10 ;
			data[59131] <= 8'h10 ;
			data[59132] <= 8'h10 ;
			data[59133] <= 8'h10 ;
			data[59134] <= 8'h10 ;
			data[59135] <= 8'h10 ;
			data[59136] <= 8'h10 ;
			data[59137] <= 8'h10 ;
			data[59138] <= 8'h10 ;
			data[59139] <= 8'h10 ;
			data[59140] <= 8'h10 ;
			data[59141] <= 8'h10 ;
			data[59142] <= 8'h10 ;
			data[59143] <= 8'h10 ;
			data[59144] <= 8'h10 ;
			data[59145] <= 8'h10 ;
			data[59146] <= 8'h10 ;
			data[59147] <= 8'h10 ;
			data[59148] <= 8'h10 ;
			data[59149] <= 8'h10 ;
			data[59150] <= 8'h10 ;
			data[59151] <= 8'h10 ;
			data[59152] <= 8'h10 ;
			data[59153] <= 8'h10 ;
			data[59154] <= 8'h10 ;
			data[59155] <= 8'h10 ;
			data[59156] <= 8'h10 ;
			data[59157] <= 8'h10 ;
			data[59158] <= 8'h10 ;
			data[59159] <= 8'h10 ;
			data[59160] <= 8'h10 ;
			data[59161] <= 8'h10 ;
			data[59162] <= 8'h10 ;
			data[59163] <= 8'h10 ;
			data[59164] <= 8'h10 ;
			data[59165] <= 8'h10 ;
			data[59166] <= 8'h10 ;
			data[59167] <= 8'h10 ;
			data[59168] <= 8'h10 ;
			data[59169] <= 8'h10 ;
			data[59170] <= 8'h10 ;
			data[59171] <= 8'h10 ;
			data[59172] <= 8'h10 ;
			data[59173] <= 8'h10 ;
			data[59174] <= 8'h10 ;
			data[59175] <= 8'h10 ;
			data[59176] <= 8'h10 ;
			data[59177] <= 8'h10 ;
			data[59178] <= 8'h10 ;
			data[59179] <= 8'h10 ;
			data[59180] <= 8'h10 ;
			data[59181] <= 8'h10 ;
			data[59182] <= 8'h10 ;
			data[59183] <= 8'h10 ;
			data[59184] <= 8'h10 ;
			data[59185] <= 8'h10 ;
			data[59186] <= 8'h10 ;
			data[59187] <= 8'h10 ;
			data[59188] <= 8'h10 ;
			data[59189] <= 8'h10 ;
			data[59190] <= 8'h10 ;
			data[59191] <= 8'h10 ;
			data[59192] <= 8'h10 ;
			data[59193] <= 8'h10 ;
			data[59194] <= 8'h10 ;
			data[59195] <= 8'h10 ;
			data[59196] <= 8'h10 ;
			data[59197] <= 8'h10 ;
			data[59198] <= 8'h10 ;
			data[59199] <= 8'h10 ;
			data[59200] <= 8'h10 ;
			data[59201] <= 8'h10 ;
			data[59202] <= 8'h10 ;
			data[59203] <= 8'h10 ;
			data[59204] <= 8'h10 ;
			data[59205] <= 8'h10 ;
			data[59206] <= 8'h10 ;
			data[59207] <= 8'h10 ;
			data[59208] <= 8'h10 ;
			data[59209] <= 8'h10 ;
			data[59210] <= 8'h10 ;
			data[59211] <= 8'h10 ;
			data[59212] <= 8'h10 ;
			data[59213] <= 8'h10 ;
			data[59214] <= 8'h10 ;
			data[59215] <= 8'h10 ;
			data[59216] <= 8'h10 ;
			data[59217] <= 8'h10 ;
			data[59218] <= 8'h10 ;
			data[59219] <= 8'h10 ;
			data[59220] <= 8'h10 ;
			data[59221] <= 8'h10 ;
			data[59222] <= 8'h10 ;
			data[59223] <= 8'h10 ;
			data[59224] <= 8'h10 ;
			data[59225] <= 8'h10 ;
			data[59226] <= 8'h10 ;
			data[59227] <= 8'h10 ;
			data[59228] <= 8'h10 ;
			data[59229] <= 8'h10 ;
			data[59230] <= 8'h10 ;
			data[59231] <= 8'h10 ;
			data[59232] <= 8'h10 ;
			data[59233] <= 8'h10 ;
			data[59234] <= 8'h10 ;
			data[59235] <= 8'h10 ;
			data[59236] <= 8'h10 ;
			data[59237] <= 8'h10 ;
			data[59238] <= 8'h10 ;
			data[59239] <= 8'h10 ;
			data[59240] <= 8'h10 ;
			data[59241] <= 8'h10 ;
			data[59242] <= 8'h10 ;
			data[59243] <= 8'h10 ;
			data[59244] <= 8'h10 ;
			data[59245] <= 8'h10 ;
			data[59246] <= 8'h10 ;
			data[59247] <= 8'h10 ;
			data[59248] <= 8'h10 ;
			data[59249] <= 8'h10 ;
			data[59250] <= 8'h10 ;
			data[59251] <= 8'h10 ;
			data[59252] <= 8'h10 ;
			data[59253] <= 8'h10 ;
			data[59254] <= 8'h10 ;
			data[59255] <= 8'h10 ;
			data[59256] <= 8'h10 ;
			data[59257] <= 8'h10 ;
			data[59258] <= 8'h10 ;
			data[59259] <= 8'h10 ;
			data[59260] <= 8'h10 ;
			data[59261] <= 8'h10 ;
			data[59262] <= 8'h10 ;
			data[59263] <= 8'h10 ;
			data[59264] <= 8'h10 ;
			data[59265] <= 8'h10 ;
			data[59266] <= 8'h10 ;
			data[59267] <= 8'h10 ;
			data[59268] <= 8'h10 ;
			data[59269] <= 8'h10 ;
			data[59270] <= 8'h10 ;
			data[59271] <= 8'h10 ;
			data[59272] <= 8'h10 ;
			data[59273] <= 8'h10 ;
			data[59274] <= 8'h10 ;
			data[59275] <= 8'h10 ;
			data[59276] <= 8'h10 ;
			data[59277] <= 8'h10 ;
			data[59278] <= 8'h10 ;
			data[59279] <= 8'h10 ;
			data[59280] <= 8'h10 ;
			data[59281] <= 8'h10 ;
			data[59282] <= 8'h10 ;
			data[59283] <= 8'h10 ;
			data[59284] <= 8'h10 ;
			data[59285] <= 8'h10 ;
			data[59286] <= 8'h10 ;
			data[59287] <= 8'h10 ;
			data[59288] <= 8'h10 ;
			data[59289] <= 8'h10 ;
			data[59290] <= 8'h10 ;
			data[59291] <= 8'h10 ;
			data[59292] <= 8'h10 ;
			data[59293] <= 8'h10 ;
			data[59294] <= 8'h10 ;
			data[59295] <= 8'h10 ;
			data[59296] <= 8'h10 ;
			data[59297] <= 8'h10 ;
			data[59298] <= 8'h10 ;
			data[59299] <= 8'h10 ;
			data[59300] <= 8'h10 ;
			data[59301] <= 8'h10 ;
			data[59302] <= 8'h10 ;
			data[59303] <= 8'h10 ;
			data[59304] <= 8'h10 ;
			data[59305] <= 8'h10 ;
			data[59306] <= 8'h10 ;
			data[59307] <= 8'h10 ;
			data[59308] <= 8'h10 ;
			data[59309] <= 8'h10 ;
			data[59310] <= 8'h10 ;
			data[59311] <= 8'h10 ;
			data[59312] <= 8'h10 ;
			data[59313] <= 8'h10 ;
			data[59314] <= 8'h10 ;
			data[59315] <= 8'h10 ;
			data[59316] <= 8'h10 ;
			data[59317] <= 8'h10 ;
			data[59318] <= 8'h10 ;
			data[59319] <= 8'h10 ;
			data[59320] <= 8'h10 ;
			data[59321] <= 8'h10 ;
			data[59322] <= 8'h10 ;
			data[59323] <= 8'h10 ;
			data[59324] <= 8'h10 ;
			data[59325] <= 8'h10 ;
			data[59326] <= 8'h10 ;
			data[59327] <= 8'h10 ;
			data[59328] <= 8'h10 ;
			data[59329] <= 8'h10 ;
			data[59330] <= 8'h10 ;
			data[59331] <= 8'h10 ;
			data[59332] <= 8'h10 ;
			data[59333] <= 8'h10 ;
			data[59334] <= 8'h10 ;
			data[59335] <= 8'h10 ;
			data[59336] <= 8'h10 ;
			data[59337] <= 8'h10 ;
			data[59338] <= 8'h10 ;
			data[59339] <= 8'h10 ;
			data[59340] <= 8'h10 ;
			data[59341] <= 8'h10 ;
			data[59342] <= 8'h10 ;
			data[59343] <= 8'h10 ;
			data[59344] <= 8'h10 ;
			data[59345] <= 8'h10 ;
			data[59346] <= 8'h10 ;
			data[59347] <= 8'h10 ;
			data[59348] <= 8'h10 ;
			data[59349] <= 8'h10 ;
			data[59350] <= 8'h10 ;
			data[59351] <= 8'h10 ;
			data[59352] <= 8'h10 ;
			data[59353] <= 8'h10 ;
			data[59354] <= 8'h10 ;
			data[59355] <= 8'h10 ;
			data[59356] <= 8'h10 ;
			data[59357] <= 8'h10 ;
			data[59358] <= 8'h10 ;
			data[59359] <= 8'h10 ;
			data[59360] <= 8'h10 ;
			data[59361] <= 8'h10 ;
			data[59362] <= 8'h10 ;
			data[59363] <= 8'h10 ;
			data[59364] <= 8'h10 ;
			data[59365] <= 8'h10 ;
			data[59366] <= 8'h10 ;
			data[59367] <= 8'h10 ;
			data[59368] <= 8'h10 ;
			data[59369] <= 8'h10 ;
			data[59370] <= 8'h10 ;
			data[59371] <= 8'h10 ;
			data[59372] <= 8'h10 ;
			data[59373] <= 8'h10 ;
			data[59374] <= 8'h10 ;
			data[59375] <= 8'h10 ;
			data[59376] <= 8'h10 ;
			data[59377] <= 8'h10 ;
			data[59378] <= 8'h10 ;
			data[59379] <= 8'h10 ;
			data[59380] <= 8'h10 ;
			data[59381] <= 8'h10 ;
			data[59382] <= 8'h10 ;
			data[59383] <= 8'h10 ;
			data[59384] <= 8'h10 ;
			data[59385] <= 8'h10 ;
			data[59386] <= 8'h10 ;
			data[59387] <= 8'h10 ;
			data[59388] <= 8'h10 ;
			data[59389] <= 8'h10 ;
			data[59390] <= 8'h10 ;
			data[59391] <= 8'h10 ;
			data[59392] <= 8'h10 ;
			data[59393] <= 8'h10 ;
			data[59394] <= 8'h10 ;
			data[59395] <= 8'h10 ;
			data[59396] <= 8'h10 ;
			data[59397] <= 8'h10 ;
			data[59398] <= 8'h10 ;
			data[59399] <= 8'h10 ;
			data[59400] <= 8'h10 ;
			data[59401] <= 8'h10 ;
			data[59402] <= 8'h10 ;
			data[59403] <= 8'h10 ;
			data[59404] <= 8'h10 ;
			data[59405] <= 8'h10 ;
			data[59406] <= 8'h10 ;
			data[59407] <= 8'h10 ;
			data[59408] <= 8'h10 ;
			data[59409] <= 8'h10 ;
			data[59410] <= 8'h10 ;
			data[59411] <= 8'h10 ;
			data[59412] <= 8'h10 ;
			data[59413] <= 8'h10 ;
			data[59414] <= 8'h10 ;
			data[59415] <= 8'h10 ;
			data[59416] <= 8'h10 ;
			data[59417] <= 8'h10 ;
			data[59418] <= 8'h10 ;
			data[59419] <= 8'h10 ;
			data[59420] <= 8'h10 ;
			data[59421] <= 8'h10 ;
			data[59422] <= 8'h10 ;
			data[59423] <= 8'h10 ;
			data[59424] <= 8'h10 ;
			data[59425] <= 8'h10 ;
			data[59426] <= 8'h10 ;
			data[59427] <= 8'h10 ;
			data[59428] <= 8'h10 ;
			data[59429] <= 8'h10 ;
			data[59430] <= 8'h10 ;
			data[59431] <= 8'h10 ;
			data[59432] <= 8'h10 ;
			data[59433] <= 8'h10 ;
			data[59434] <= 8'h10 ;
			data[59435] <= 8'h10 ;
			data[59436] <= 8'h10 ;
			data[59437] <= 8'h10 ;
			data[59438] <= 8'h10 ;
			data[59439] <= 8'h10 ;
			data[59440] <= 8'h10 ;
			data[59441] <= 8'h10 ;
			data[59442] <= 8'h10 ;
			data[59443] <= 8'h10 ;
			data[59444] <= 8'h10 ;
			data[59445] <= 8'h10 ;
			data[59446] <= 8'h10 ;
			data[59447] <= 8'h10 ;
			data[59448] <= 8'h10 ;
			data[59449] <= 8'h10 ;
			data[59450] <= 8'h10 ;
			data[59451] <= 8'h10 ;
			data[59452] <= 8'h10 ;
			data[59453] <= 8'h10 ;
			data[59454] <= 8'h10 ;
			data[59455] <= 8'h10 ;
			data[59456] <= 8'h10 ;
			data[59457] <= 8'h10 ;
			data[59458] <= 8'h10 ;
			data[59459] <= 8'h10 ;
			data[59460] <= 8'h10 ;
			data[59461] <= 8'h10 ;
			data[59462] <= 8'h10 ;
			data[59463] <= 8'h10 ;
			data[59464] <= 8'h10 ;
			data[59465] <= 8'h10 ;
			data[59466] <= 8'h10 ;
			data[59467] <= 8'h10 ;
			data[59468] <= 8'h10 ;
			data[59469] <= 8'h10 ;
			data[59470] <= 8'h10 ;
			data[59471] <= 8'h10 ;
			data[59472] <= 8'h10 ;
			data[59473] <= 8'h10 ;
			data[59474] <= 8'h10 ;
			data[59475] <= 8'h10 ;
			data[59476] <= 8'h10 ;
			data[59477] <= 8'h10 ;
			data[59478] <= 8'h10 ;
			data[59479] <= 8'h10 ;
			data[59480] <= 8'h10 ;
			data[59481] <= 8'h10 ;
			data[59482] <= 8'h10 ;
			data[59483] <= 8'h10 ;
			data[59484] <= 8'h10 ;
			data[59485] <= 8'h10 ;
			data[59486] <= 8'h10 ;
			data[59487] <= 8'h10 ;
			data[59488] <= 8'h10 ;
			data[59489] <= 8'h10 ;
			data[59490] <= 8'h10 ;
			data[59491] <= 8'h10 ;
			data[59492] <= 8'h10 ;
			data[59493] <= 8'h10 ;
			data[59494] <= 8'h10 ;
			data[59495] <= 8'h10 ;
			data[59496] <= 8'h10 ;
			data[59497] <= 8'h10 ;
			data[59498] <= 8'h10 ;
			data[59499] <= 8'h10 ;
			data[59500] <= 8'h10 ;
			data[59501] <= 8'h10 ;
			data[59502] <= 8'h10 ;
			data[59503] <= 8'h10 ;
			data[59504] <= 8'h10 ;
			data[59505] <= 8'h10 ;
			data[59506] <= 8'h10 ;
			data[59507] <= 8'h10 ;
			data[59508] <= 8'h10 ;
			data[59509] <= 8'h10 ;
			data[59510] <= 8'h10 ;
			data[59511] <= 8'h10 ;
			data[59512] <= 8'h10 ;
			data[59513] <= 8'h10 ;
			data[59514] <= 8'h10 ;
			data[59515] <= 8'h10 ;
			data[59516] <= 8'h10 ;
			data[59517] <= 8'h10 ;
			data[59518] <= 8'h10 ;
			data[59519] <= 8'h10 ;
			data[59520] <= 8'h10 ;
			data[59521] <= 8'h10 ;
			data[59522] <= 8'h10 ;
			data[59523] <= 8'h10 ;
			data[59524] <= 8'h10 ;
			data[59525] <= 8'h10 ;
			data[59526] <= 8'h10 ;
			data[59527] <= 8'h10 ;
			data[59528] <= 8'h10 ;
			data[59529] <= 8'h10 ;
			data[59530] <= 8'h10 ;
			data[59531] <= 8'h10 ;
			data[59532] <= 8'h10 ;
			data[59533] <= 8'h10 ;
			data[59534] <= 8'h10 ;
			data[59535] <= 8'h10 ;
			data[59536] <= 8'h10 ;
			data[59537] <= 8'h10 ;
			data[59538] <= 8'h10 ;
			data[59539] <= 8'h10 ;
			data[59540] <= 8'h10 ;
			data[59541] <= 8'h10 ;
			data[59542] <= 8'h10 ;
			data[59543] <= 8'h10 ;
			data[59544] <= 8'h10 ;
			data[59545] <= 8'h10 ;
			data[59546] <= 8'h10 ;
			data[59547] <= 8'h10 ;
			data[59548] <= 8'h10 ;
			data[59549] <= 8'h10 ;
			data[59550] <= 8'h10 ;
			data[59551] <= 8'h10 ;
			data[59552] <= 8'h10 ;
			data[59553] <= 8'h10 ;
			data[59554] <= 8'h10 ;
			data[59555] <= 8'h10 ;
			data[59556] <= 8'h10 ;
			data[59557] <= 8'h10 ;
			data[59558] <= 8'h10 ;
			data[59559] <= 8'h10 ;
			data[59560] <= 8'h10 ;
			data[59561] <= 8'h10 ;
			data[59562] <= 8'h10 ;
			data[59563] <= 8'h10 ;
			data[59564] <= 8'h10 ;
			data[59565] <= 8'h10 ;
			data[59566] <= 8'h10 ;
			data[59567] <= 8'h10 ;
			data[59568] <= 8'h10 ;
			data[59569] <= 8'h10 ;
			data[59570] <= 8'h10 ;
			data[59571] <= 8'h10 ;
			data[59572] <= 8'h10 ;
			data[59573] <= 8'h10 ;
			data[59574] <= 8'h10 ;
			data[59575] <= 8'h10 ;
			data[59576] <= 8'h10 ;
			data[59577] <= 8'h10 ;
			data[59578] <= 8'h10 ;
			data[59579] <= 8'h10 ;
			data[59580] <= 8'h10 ;
			data[59581] <= 8'h10 ;
			data[59582] <= 8'h10 ;
			data[59583] <= 8'h10 ;
			data[59584] <= 8'h10 ;
			data[59585] <= 8'h10 ;
			data[59586] <= 8'h10 ;
			data[59587] <= 8'h10 ;
			data[59588] <= 8'h10 ;
			data[59589] <= 8'h10 ;
			data[59590] <= 8'h10 ;
			data[59591] <= 8'h10 ;
			data[59592] <= 8'h10 ;
			data[59593] <= 8'h10 ;
			data[59594] <= 8'h10 ;
			data[59595] <= 8'h10 ;
			data[59596] <= 8'h10 ;
			data[59597] <= 8'h10 ;
			data[59598] <= 8'h10 ;
			data[59599] <= 8'h10 ;
			data[59600] <= 8'h10 ;
			data[59601] <= 8'h10 ;
			data[59602] <= 8'h10 ;
			data[59603] <= 8'h10 ;
			data[59604] <= 8'h10 ;
			data[59605] <= 8'h10 ;
			data[59606] <= 8'h10 ;
			data[59607] <= 8'h10 ;
			data[59608] <= 8'h10 ;
			data[59609] <= 8'h10 ;
			data[59610] <= 8'h10 ;
			data[59611] <= 8'h10 ;
			data[59612] <= 8'h10 ;
			data[59613] <= 8'h10 ;
			data[59614] <= 8'h10 ;
			data[59615] <= 8'h10 ;
			data[59616] <= 8'h10 ;
			data[59617] <= 8'h10 ;
			data[59618] <= 8'h10 ;
			data[59619] <= 8'h10 ;
			data[59620] <= 8'h10 ;
			data[59621] <= 8'h10 ;
			data[59622] <= 8'h10 ;
			data[59623] <= 8'h10 ;
			data[59624] <= 8'h10 ;
			data[59625] <= 8'h10 ;
			data[59626] <= 8'h10 ;
			data[59627] <= 8'h10 ;
			data[59628] <= 8'h10 ;
			data[59629] <= 8'h10 ;
			data[59630] <= 8'h10 ;
			data[59631] <= 8'h10 ;
			data[59632] <= 8'h10 ;
			data[59633] <= 8'h10 ;
			data[59634] <= 8'h10 ;
			data[59635] <= 8'h10 ;
			data[59636] <= 8'h10 ;
			data[59637] <= 8'h10 ;
			data[59638] <= 8'h10 ;
			data[59639] <= 8'h10 ;
			data[59640] <= 8'h10 ;
			data[59641] <= 8'h10 ;
			data[59642] <= 8'h10 ;
			data[59643] <= 8'h10 ;
			data[59644] <= 8'h10 ;
			data[59645] <= 8'h10 ;
			data[59646] <= 8'h10 ;
			data[59647] <= 8'h10 ;
			data[59648] <= 8'h10 ;
			data[59649] <= 8'h10 ;
			data[59650] <= 8'h10 ;
			data[59651] <= 8'h10 ;
			data[59652] <= 8'h10 ;
			data[59653] <= 8'h10 ;
			data[59654] <= 8'h10 ;
			data[59655] <= 8'h10 ;
			data[59656] <= 8'h10 ;
			data[59657] <= 8'h10 ;
			data[59658] <= 8'h10 ;
			data[59659] <= 8'h10 ;
			data[59660] <= 8'h10 ;
			data[59661] <= 8'h10 ;
			data[59662] <= 8'h10 ;
			data[59663] <= 8'h10 ;
			data[59664] <= 8'h10 ;
			data[59665] <= 8'h10 ;
			data[59666] <= 8'h10 ;
			data[59667] <= 8'h10 ;
			data[59668] <= 8'h10 ;
			data[59669] <= 8'h10 ;
			data[59670] <= 8'h10 ;
			data[59671] <= 8'h10 ;
			data[59672] <= 8'h10 ;
			data[59673] <= 8'h10 ;
			data[59674] <= 8'h10 ;
			data[59675] <= 8'h10 ;
			data[59676] <= 8'h10 ;
			data[59677] <= 8'h10 ;
			data[59678] <= 8'h10 ;
			data[59679] <= 8'h10 ;
			data[59680] <= 8'h10 ;
			data[59681] <= 8'h10 ;
			data[59682] <= 8'h10 ;
			data[59683] <= 8'h10 ;
			data[59684] <= 8'h10 ;
			data[59685] <= 8'h10 ;
			data[59686] <= 8'h10 ;
			data[59687] <= 8'h10 ;
			data[59688] <= 8'h10 ;
			data[59689] <= 8'h10 ;
			data[59690] <= 8'h10 ;
			data[59691] <= 8'h10 ;
			data[59692] <= 8'h10 ;
			data[59693] <= 8'h10 ;
			data[59694] <= 8'h10 ;
			data[59695] <= 8'h10 ;
			data[59696] <= 8'h10 ;
			data[59697] <= 8'h10 ;
			data[59698] <= 8'h10 ;
			data[59699] <= 8'h10 ;
			data[59700] <= 8'h10 ;
			data[59701] <= 8'h10 ;
			data[59702] <= 8'h10 ;
			data[59703] <= 8'h10 ;
			data[59704] <= 8'h10 ;
			data[59705] <= 8'h10 ;
			data[59706] <= 8'h10 ;
			data[59707] <= 8'h10 ;
			data[59708] <= 8'h10 ;
			data[59709] <= 8'h10 ;
			data[59710] <= 8'h10 ;
			data[59711] <= 8'h10 ;
			data[59712] <= 8'h10 ;
			data[59713] <= 8'h10 ;
			data[59714] <= 8'h10 ;
			data[59715] <= 8'h10 ;
			data[59716] <= 8'h10 ;
			data[59717] <= 8'h10 ;
			data[59718] <= 8'h10 ;
			data[59719] <= 8'h10 ;
			data[59720] <= 8'h10 ;
			data[59721] <= 8'h10 ;
			data[59722] <= 8'h10 ;
			data[59723] <= 8'h10 ;
			data[59724] <= 8'h10 ;
			data[59725] <= 8'h10 ;
			data[59726] <= 8'h10 ;
			data[59727] <= 8'h10 ;
			data[59728] <= 8'h10 ;
			data[59729] <= 8'h10 ;
			data[59730] <= 8'h10 ;
			data[59731] <= 8'h10 ;
			data[59732] <= 8'h10 ;
			data[59733] <= 8'h10 ;
			data[59734] <= 8'h10 ;
			data[59735] <= 8'h10 ;
			data[59736] <= 8'h10 ;
			data[59737] <= 8'h10 ;
			data[59738] <= 8'h10 ;
			data[59739] <= 8'h10 ;
			data[59740] <= 8'h10 ;
			data[59741] <= 8'h10 ;
			data[59742] <= 8'h10 ;
			data[59743] <= 8'h10 ;
			data[59744] <= 8'h10 ;
			data[59745] <= 8'h10 ;
			data[59746] <= 8'h10 ;
			data[59747] <= 8'h10 ;
			data[59748] <= 8'h10 ;
			data[59749] <= 8'h10 ;
			data[59750] <= 8'h10 ;
			data[59751] <= 8'h10 ;
			data[59752] <= 8'h10 ;
			data[59753] <= 8'h10 ;
			data[59754] <= 8'h10 ;
			data[59755] <= 8'h10 ;
			data[59756] <= 8'h10 ;
			data[59757] <= 8'h10 ;
			data[59758] <= 8'h10 ;
			data[59759] <= 8'h10 ;
			data[59760] <= 8'h10 ;
			data[59761] <= 8'h10 ;
			data[59762] <= 8'h10 ;
			data[59763] <= 8'h10 ;
			data[59764] <= 8'h10 ;
			data[59765] <= 8'h10 ;
			data[59766] <= 8'h10 ;
			data[59767] <= 8'h10 ;
			data[59768] <= 8'h10 ;
			data[59769] <= 8'h10 ;
			data[59770] <= 8'h10 ;
			data[59771] <= 8'h10 ;
			data[59772] <= 8'h10 ;
			data[59773] <= 8'h10 ;
			data[59774] <= 8'h10 ;
			data[59775] <= 8'h10 ;
			data[59776] <= 8'h10 ;
			data[59777] <= 8'h10 ;
			data[59778] <= 8'h10 ;
			data[59779] <= 8'h10 ;
			data[59780] <= 8'h10 ;
			data[59781] <= 8'h10 ;
			data[59782] <= 8'h10 ;
			data[59783] <= 8'h10 ;
			data[59784] <= 8'h10 ;
			data[59785] <= 8'h10 ;
			data[59786] <= 8'h10 ;
			data[59787] <= 8'h10 ;
			data[59788] <= 8'h10 ;
			data[59789] <= 8'h10 ;
			data[59790] <= 8'h10 ;
			data[59791] <= 8'h10 ;
			data[59792] <= 8'h10 ;
			data[59793] <= 8'h10 ;
			data[59794] <= 8'h10 ;
			data[59795] <= 8'h10 ;
			data[59796] <= 8'h10 ;
			data[59797] <= 8'h10 ;
			data[59798] <= 8'h10 ;
			data[59799] <= 8'h10 ;
			data[59800] <= 8'h10 ;
			data[59801] <= 8'h10 ;
			data[59802] <= 8'h10 ;
			data[59803] <= 8'h10 ;
			data[59804] <= 8'h10 ;
			data[59805] <= 8'h10 ;
			data[59806] <= 8'h10 ;
			data[59807] <= 8'h10 ;
			data[59808] <= 8'h10 ;
			data[59809] <= 8'h10 ;
			data[59810] <= 8'h10 ;
			data[59811] <= 8'h10 ;
			data[59812] <= 8'h10 ;
			data[59813] <= 8'h10 ;
			data[59814] <= 8'h10 ;
			data[59815] <= 8'h10 ;
			data[59816] <= 8'h10 ;
			data[59817] <= 8'h10 ;
			data[59818] <= 8'h10 ;
			data[59819] <= 8'h10 ;
			data[59820] <= 8'h10 ;
			data[59821] <= 8'h10 ;
			data[59822] <= 8'h10 ;
			data[59823] <= 8'h10 ;
			data[59824] <= 8'h10 ;
			data[59825] <= 8'h10 ;
			data[59826] <= 8'h10 ;
			data[59827] <= 8'h10 ;
			data[59828] <= 8'h10 ;
			data[59829] <= 8'h10 ;
			data[59830] <= 8'h10 ;
			data[59831] <= 8'h10 ;
			data[59832] <= 8'h10 ;
			data[59833] <= 8'h10 ;
			data[59834] <= 8'h10 ;
			data[59835] <= 8'h10 ;
			data[59836] <= 8'h10 ;
			data[59837] <= 8'h10 ;
			data[59838] <= 8'h10 ;
			data[59839] <= 8'h10 ;
			data[59840] <= 8'h10 ;
			data[59841] <= 8'h10 ;
			data[59842] <= 8'h10 ;
			data[59843] <= 8'h10 ;
			data[59844] <= 8'h10 ;
			data[59845] <= 8'h10 ;
			data[59846] <= 8'h10 ;
			data[59847] <= 8'h10 ;
			data[59848] <= 8'h10 ;
			data[59849] <= 8'h10 ;
			data[59850] <= 8'h10 ;
			data[59851] <= 8'h10 ;
			data[59852] <= 8'h10 ;
			data[59853] <= 8'h10 ;
			data[59854] <= 8'h10 ;
			data[59855] <= 8'h10 ;
			data[59856] <= 8'h10 ;
			data[59857] <= 8'h10 ;
			data[59858] <= 8'h10 ;
			data[59859] <= 8'h10 ;
			data[59860] <= 8'h10 ;
			data[59861] <= 8'h10 ;
			data[59862] <= 8'h10 ;
			data[59863] <= 8'h10 ;
			data[59864] <= 8'h10 ;
			data[59865] <= 8'h10 ;
			data[59866] <= 8'h10 ;
			data[59867] <= 8'h10 ;
			data[59868] <= 8'h10 ;
			data[59869] <= 8'h10 ;
			data[59870] <= 8'h10 ;
			data[59871] <= 8'h10 ;
			data[59872] <= 8'h10 ;
			data[59873] <= 8'h10 ;
			data[59874] <= 8'h10 ;
			data[59875] <= 8'h10 ;
			data[59876] <= 8'h10 ;
			data[59877] <= 8'h10 ;
			data[59878] <= 8'h10 ;
			data[59879] <= 8'h10 ;
			data[59880] <= 8'h10 ;
			data[59881] <= 8'h10 ;
			data[59882] <= 8'h10 ;
			data[59883] <= 8'h10 ;
			data[59884] <= 8'h10 ;
			data[59885] <= 8'h10 ;
			data[59886] <= 8'h10 ;
			data[59887] <= 8'h10 ;
			data[59888] <= 8'h10 ;
			data[59889] <= 8'h10 ;
			data[59890] <= 8'h10 ;
			data[59891] <= 8'h10 ;
			data[59892] <= 8'h10 ;
			data[59893] <= 8'h10 ;
			data[59894] <= 8'h10 ;
			data[59895] <= 8'h10 ;
			data[59896] <= 8'h10 ;
			data[59897] <= 8'h10 ;
			data[59898] <= 8'h10 ;
			data[59899] <= 8'h10 ;
			data[59900] <= 8'h10 ;
			data[59901] <= 8'h10 ;
			data[59902] <= 8'h10 ;
			data[59903] <= 8'h10 ;
			data[59904] <= 8'h10 ;
			data[59905] <= 8'h10 ;
			data[59906] <= 8'h10 ;
			data[59907] <= 8'h10 ;
			data[59908] <= 8'h10 ;
			data[59909] <= 8'h10 ;
			data[59910] <= 8'h10 ;
			data[59911] <= 8'h10 ;
			data[59912] <= 8'h10 ;
			data[59913] <= 8'h10 ;
			data[59914] <= 8'h10 ;
			data[59915] <= 8'h10 ;
			data[59916] <= 8'h10 ;
			data[59917] <= 8'h10 ;
			data[59918] <= 8'h10 ;
			data[59919] <= 8'h10 ;
			data[59920] <= 8'h10 ;
			data[59921] <= 8'h10 ;
			data[59922] <= 8'h10 ;
			data[59923] <= 8'h10 ;
			data[59924] <= 8'h10 ;
			data[59925] <= 8'h10 ;
			data[59926] <= 8'h10 ;
			data[59927] <= 8'h10 ;
			data[59928] <= 8'h10 ;
			data[59929] <= 8'h10 ;
			data[59930] <= 8'h10 ;
			data[59931] <= 8'h10 ;
			data[59932] <= 8'h10 ;
			data[59933] <= 8'h10 ;
			data[59934] <= 8'h10 ;
			data[59935] <= 8'h10 ;
			data[59936] <= 8'h10 ;
			data[59937] <= 8'h10 ;
			data[59938] <= 8'h10 ;
			data[59939] <= 8'h10 ;
			data[59940] <= 8'h10 ;
			data[59941] <= 8'h10 ;
			data[59942] <= 8'h10 ;
			data[59943] <= 8'h10 ;
			data[59944] <= 8'h10 ;
			data[59945] <= 8'h10 ;
			data[59946] <= 8'h10 ;
			data[59947] <= 8'h10 ;
			data[59948] <= 8'h10 ;
			data[59949] <= 8'h10 ;
			data[59950] <= 8'h10 ;
			data[59951] <= 8'h10 ;
			data[59952] <= 8'h10 ;
			data[59953] <= 8'h10 ;
			data[59954] <= 8'h10 ;
			data[59955] <= 8'h10 ;
			data[59956] <= 8'h10 ;
			data[59957] <= 8'h10 ;
			data[59958] <= 8'h10 ;
			data[59959] <= 8'h10 ;
			data[59960] <= 8'h10 ;
			data[59961] <= 8'h10 ;
			data[59962] <= 8'h10 ;
			data[59963] <= 8'h10 ;
			data[59964] <= 8'h10 ;
			data[59965] <= 8'h10 ;
			data[59966] <= 8'h10 ;
			data[59967] <= 8'h10 ;
			data[59968] <= 8'h10 ;
			data[59969] <= 8'h10 ;
			data[59970] <= 8'h10 ;
			data[59971] <= 8'h10 ;
			data[59972] <= 8'h10 ;
			data[59973] <= 8'h10 ;
			data[59974] <= 8'h10 ;
			data[59975] <= 8'h10 ;
			data[59976] <= 8'h10 ;
			data[59977] <= 8'h10 ;
			data[59978] <= 8'h10 ;
			data[59979] <= 8'h10 ;
			data[59980] <= 8'h10 ;
			data[59981] <= 8'h10 ;
			data[59982] <= 8'h10 ;
			data[59983] <= 8'h10 ;
			data[59984] <= 8'h10 ;
			data[59985] <= 8'h10 ;
			data[59986] <= 8'h10 ;
			data[59987] <= 8'h10 ;
			data[59988] <= 8'h10 ;
			data[59989] <= 8'h10 ;
			data[59990] <= 8'h10 ;
			data[59991] <= 8'h10 ;
			data[59992] <= 8'h10 ;
			data[59993] <= 8'h10 ;
			data[59994] <= 8'h10 ;
			data[59995] <= 8'h10 ;
			data[59996] <= 8'h10 ;
			data[59997] <= 8'h10 ;
			data[59998] <= 8'h10 ;
			data[59999] <= 8'h10 ;
			data[60000] <= 8'h10 ;
			data[60001] <= 8'h10 ;
			data[60002] <= 8'h10 ;
			data[60003] <= 8'h10 ;
			data[60004] <= 8'h10 ;
			data[60005] <= 8'h10 ;
			data[60006] <= 8'h10 ;
			data[60007] <= 8'h10 ;
			data[60008] <= 8'h10 ;
			data[60009] <= 8'h10 ;
			data[60010] <= 8'h10 ;
			data[60011] <= 8'h10 ;
			data[60012] <= 8'h10 ;
			data[60013] <= 8'h10 ;
			data[60014] <= 8'h10 ;
			data[60015] <= 8'h10 ;
			data[60016] <= 8'h10 ;
			data[60017] <= 8'h10 ;
			data[60018] <= 8'h10 ;
			data[60019] <= 8'h10 ;
			data[60020] <= 8'h10 ;
			data[60021] <= 8'h10 ;
			data[60022] <= 8'h10 ;
			data[60023] <= 8'h10 ;
			data[60024] <= 8'h10 ;
			data[60025] <= 8'h10 ;
			data[60026] <= 8'h10 ;
			data[60027] <= 8'h10 ;
			data[60028] <= 8'h10 ;
			data[60029] <= 8'h10 ;
			data[60030] <= 8'h10 ;
			data[60031] <= 8'h10 ;
			data[60032] <= 8'h10 ;
			data[60033] <= 8'h10 ;
			data[60034] <= 8'h10 ;
			data[60035] <= 8'h10 ;
			data[60036] <= 8'h10 ;
			data[60037] <= 8'h10 ;
			data[60038] <= 8'h10 ;
			data[60039] <= 8'h10 ;
			data[60040] <= 8'h10 ;
			data[60041] <= 8'h10 ;
			data[60042] <= 8'h10 ;
			data[60043] <= 8'h10 ;
			data[60044] <= 8'h10 ;
			data[60045] <= 8'h10 ;
			data[60046] <= 8'h10 ;
			data[60047] <= 8'h10 ;
			data[60048] <= 8'h10 ;
			data[60049] <= 8'h10 ;
			data[60050] <= 8'h10 ;
			data[60051] <= 8'h10 ;
			data[60052] <= 8'h10 ;
			data[60053] <= 8'h10 ;
			data[60054] <= 8'h10 ;
			data[60055] <= 8'h10 ;
			data[60056] <= 8'h10 ;
			data[60057] <= 8'h10 ;
			data[60058] <= 8'h10 ;
			data[60059] <= 8'h10 ;
			data[60060] <= 8'h10 ;
			data[60061] <= 8'h10 ;
			data[60062] <= 8'h10 ;
			data[60063] <= 8'h10 ;
			data[60064] <= 8'h10 ;
			data[60065] <= 8'h10 ;
			data[60066] <= 8'h10 ;
			data[60067] <= 8'h10 ;
			data[60068] <= 8'h10 ;
			data[60069] <= 8'h10 ;
			data[60070] <= 8'h10 ;
			data[60071] <= 8'h10 ;
			data[60072] <= 8'h10 ;
			data[60073] <= 8'h10 ;
			data[60074] <= 8'h10 ;
			data[60075] <= 8'h10 ;
			data[60076] <= 8'h10 ;
			data[60077] <= 8'h10 ;
			data[60078] <= 8'h10 ;
			data[60079] <= 8'h10 ;
			data[60080] <= 8'h10 ;
			data[60081] <= 8'h10 ;
			data[60082] <= 8'h10 ;
			data[60083] <= 8'h10 ;
			data[60084] <= 8'h10 ;
			data[60085] <= 8'h10 ;
			data[60086] <= 8'h10 ;
			data[60087] <= 8'h10 ;
			data[60088] <= 8'h10 ;
			data[60089] <= 8'h10 ;
			data[60090] <= 8'h10 ;
			data[60091] <= 8'h10 ;
			data[60092] <= 8'h10 ;
			data[60093] <= 8'h10 ;
			data[60094] <= 8'h10 ;
			data[60095] <= 8'h10 ;
			data[60096] <= 8'h10 ;
			data[60097] <= 8'h10 ;
			data[60098] <= 8'h10 ;
			data[60099] <= 8'h10 ;
			data[60100] <= 8'h10 ;
			data[60101] <= 8'h10 ;
			data[60102] <= 8'h10 ;
			data[60103] <= 8'h10 ;
			data[60104] <= 8'h10 ;
			data[60105] <= 8'h10 ;
			data[60106] <= 8'h10 ;
			data[60107] <= 8'h10 ;
			data[60108] <= 8'h10 ;
			data[60109] <= 8'h10 ;
			data[60110] <= 8'h10 ;
			data[60111] <= 8'h10 ;
			data[60112] <= 8'h10 ;
			data[60113] <= 8'h10 ;
			data[60114] <= 8'h10 ;
			data[60115] <= 8'h10 ;
			data[60116] <= 8'h10 ;
			data[60117] <= 8'h10 ;
			data[60118] <= 8'h10 ;
			data[60119] <= 8'h10 ;
			data[60120] <= 8'h10 ;
			data[60121] <= 8'h10 ;
			data[60122] <= 8'h10 ;
			data[60123] <= 8'h10 ;
			data[60124] <= 8'h10 ;
			data[60125] <= 8'h10 ;
			data[60126] <= 8'h10 ;
			data[60127] <= 8'h10 ;
			data[60128] <= 8'h10 ;
			data[60129] <= 8'h10 ;
			data[60130] <= 8'h10 ;
			data[60131] <= 8'h10 ;
			data[60132] <= 8'h10 ;
			data[60133] <= 8'h10 ;
			data[60134] <= 8'h10 ;
			data[60135] <= 8'h10 ;
			data[60136] <= 8'h10 ;
			data[60137] <= 8'h10 ;
			data[60138] <= 8'h10 ;
			data[60139] <= 8'h10 ;
			data[60140] <= 8'h10 ;
			data[60141] <= 8'h10 ;
			data[60142] <= 8'h10 ;
			data[60143] <= 8'h10 ;
			data[60144] <= 8'h10 ;
			data[60145] <= 8'h10 ;
			data[60146] <= 8'h10 ;
			data[60147] <= 8'h10 ;
			data[60148] <= 8'h10 ;
			data[60149] <= 8'h10 ;
			data[60150] <= 8'h10 ;
			data[60151] <= 8'h10 ;
			data[60152] <= 8'h10 ;
			data[60153] <= 8'h10 ;
			data[60154] <= 8'h10 ;
			data[60155] <= 8'h10 ;
			data[60156] <= 8'h10 ;
			data[60157] <= 8'h10 ;
			data[60158] <= 8'h10 ;
			data[60159] <= 8'h10 ;
			data[60160] <= 8'h10 ;
			data[60161] <= 8'h10 ;
			data[60162] <= 8'h10 ;
			data[60163] <= 8'h10 ;
			data[60164] <= 8'h10 ;
			data[60165] <= 8'h10 ;
			data[60166] <= 8'h10 ;
			data[60167] <= 8'h10 ;
			data[60168] <= 8'h10 ;
			data[60169] <= 8'h10 ;
			data[60170] <= 8'h10 ;
			data[60171] <= 8'h10 ;
			data[60172] <= 8'h10 ;
			data[60173] <= 8'h10 ;
			data[60174] <= 8'h10 ;
			data[60175] <= 8'h10 ;
			data[60176] <= 8'h10 ;
			data[60177] <= 8'h10 ;
			data[60178] <= 8'h10 ;
			data[60179] <= 8'h10 ;
			data[60180] <= 8'h10 ;
			data[60181] <= 8'h10 ;
			data[60182] <= 8'h10 ;
			data[60183] <= 8'h10 ;
			data[60184] <= 8'h10 ;
			data[60185] <= 8'h10 ;
			data[60186] <= 8'h10 ;
			data[60187] <= 8'h10 ;
			data[60188] <= 8'h10 ;
			data[60189] <= 8'h10 ;
			data[60190] <= 8'h10 ;
			data[60191] <= 8'h10 ;
			data[60192] <= 8'h10 ;
			data[60193] <= 8'h10 ;
			data[60194] <= 8'h10 ;
			data[60195] <= 8'h10 ;
			data[60196] <= 8'h10 ;
			data[60197] <= 8'h10 ;
			data[60198] <= 8'h10 ;
			data[60199] <= 8'h10 ;
			data[60200] <= 8'h10 ;
			data[60201] <= 8'h10 ;
			data[60202] <= 8'h10 ;
			data[60203] <= 8'h10 ;
			data[60204] <= 8'h10 ;
			data[60205] <= 8'h10 ;
			data[60206] <= 8'h10 ;
			data[60207] <= 8'h10 ;
			data[60208] <= 8'h10 ;
			data[60209] <= 8'h10 ;
			data[60210] <= 8'h10 ;
			data[60211] <= 8'h10 ;
			data[60212] <= 8'h10 ;
			data[60213] <= 8'h10 ;
			data[60214] <= 8'h10 ;
			data[60215] <= 8'h10 ;
			data[60216] <= 8'h10 ;
			data[60217] <= 8'h10 ;
			data[60218] <= 8'h10 ;
			data[60219] <= 8'h10 ;
			data[60220] <= 8'h10 ;
			data[60221] <= 8'h10 ;
			data[60222] <= 8'h10 ;
			data[60223] <= 8'h10 ;
			data[60224] <= 8'h10 ;
			data[60225] <= 8'h10 ;
			data[60226] <= 8'h10 ;
			data[60227] <= 8'h10 ;
			data[60228] <= 8'h10 ;
			data[60229] <= 8'h10 ;
			data[60230] <= 8'h10 ;
			data[60231] <= 8'h10 ;
			data[60232] <= 8'h10 ;
			data[60233] <= 8'h10 ;
			data[60234] <= 8'h10 ;
			data[60235] <= 8'h10 ;
			data[60236] <= 8'h10 ;
			data[60237] <= 8'h10 ;
			data[60238] <= 8'h10 ;
			data[60239] <= 8'h10 ;
			data[60240] <= 8'h10 ;
			data[60241] <= 8'h10 ;
			data[60242] <= 8'h10 ;
			data[60243] <= 8'h10 ;
			data[60244] <= 8'h10 ;
			data[60245] <= 8'h10 ;
			data[60246] <= 8'h10 ;
			data[60247] <= 8'h10 ;
			data[60248] <= 8'h10 ;
			data[60249] <= 8'h10 ;
			data[60250] <= 8'h10 ;
			data[60251] <= 8'h10 ;
			data[60252] <= 8'h10 ;
			data[60253] <= 8'h10 ;
			data[60254] <= 8'h10 ;
			data[60255] <= 8'h10 ;
			data[60256] <= 8'h10 ;
			data[60257] <= 8'h10 ;
			data[60258] <= 8'h10 ;
			data[60259] <= 8'h10 ;
			data[60260] <= 8'h10 ;
			data[60261] <= 8'h10 ;
			data[60262] <= 8'h10 ;
			data[60263] <= 8'h10 ;
			data[60264] <= 8'h10 ;
			data[60265] <= 8'h10 ;
			data[60266] <= 8'h10 ;
			data[60267] <= 8'h10 ;
			data[60268] <= 8'h10 ;
			data[60269] <= 8'h10 ;
			data[60270] <= 8'h10 ;
			data[60271] <= 8'h10 ;
			data[60272] <= 8'h10 ;
			data[60273] <= 8'h10 ;
			data[60274] <= 8'h10 ;
			data[60275] <= 8'h10 ;
			data[60276] <= 8'h10 ;
			data[60277] <= 8'h10 ;
			data[60278] <= 8'h10 ;
			data[60279] <= 8'h10 ;
			data[60280] <= 8'h10 ;
			data[60281] <= 8'h10 ;
			data[60282] <= 8'h10 ;
			data[60283] <= 8'h10 ;
			data[60284] <= 8'h10 ;
			data[60285] <= 8'h10 ;
			data[60286] <= 8'h10 ;
			data[60287] <= 8'h10 ;
			data[60288] <= 8'h10 ;
			data[60289] <= 8'h10 ;
			data[60290] <= 8'h10 ;
			data[60291] <= 8'h10 ;
			data[60292] <= 8'h10 ;
			data[60293] <= 8'h10 ;
			data[60294] <= 8'h10 ;
			data[60295] <= 8'h10 ;
			data[60296] <= 8'h10 ;
			data[60297] <= 8'h10 ;
			data[60298] <= 8'h10 ;
			data[60299] <= 8'h10 ;
			data[60300] <= 8'h10 ;
			data[60301] <= 8'h10 ;
			data[60302] <= 8'h10 ;
			data[60303] <= 8'h10 ;
			data[60304] <= 8'h10 ;
			data[60305] <= 8'h10 ;
			data[60306] <= 8'h10 ;
			data[60307] <= 8'h10 ;
			data[60308] <= 8'h10 ;
			data[60309] <= 8'h10 ;
			data[60310] <= 8'h10 ;
			data[60311] <= 8'h10 ;
			data[60312] <= 8'h10 ;
			data[60313] <= 8'h10 ;
			data[60314] <= 8'h10 ;
			data[60315] <= 8'h10 ;
			data[60316] <= 8'h10 ;
			data[60317] <= 8'h10 ;
			data[60318] <= 8'h10 ;
			data[60319] <= 8'h10 ;
			data[60320] <= 8'h10 ;
			data[60321] <= 8'h10 ;
			data[60322] <= 8'h10 ;
			data[60323] <= 8'h10 ;
			data[60324] <= 8'h10 ;
			data[60325] <= 8'h10 ;
			data[60326] <= 8'h10 ;
			data[60327] <= 8'h10 ;
			data[60328] <= 8'h10 ;
			data[60329] <= 8'h10 ;
			data[60330] <= 8'h10 ;
			data[60331] <= 8'h10 ;
			data[60332] <= 8'h10 ;
			data[60333] <= 8'h10 ;
			data[60334] <= 8'h10 ;
			data[60335] <= 8'h10 ;
			data[60336] <= 8'h10 ;
			data[60337] <= 8'h10 ;
			data[60338] <= 8'h10 ;
			data[60339] <= 8'h10 ;
			data[60340] <= 8'h10 ;
			data[60341] <= 8'h10 ;
			data[60342] <= 8'h10 ;
			data[60343] <= 8'h10 ;
			data[60344] <= 8'h10 ;
			data[60345] <= 8'h10 ;
			data[60346] <= 8'h10 ;
			data[60347] <= 8'h10 ;
			data[60348] <= 8'h10 ;
			data[60349] <= 8'h10 ;
			data[60350] <= 8'h10 ;
			data[60351] <= 8'h10 ;
			data[60352] <= 8'h10 ;
			data[60353] <= 8'h10 ;
			data[60354] <= 8'h10 ;
			data[60355] <= 8'h10 ;
			data[60356] <= 8'h10 ;
			data[60357] <= 8'h10 ;
			data[60358] <= 8'h10 ;
			data[60359] <= 8'h10 ;
			data[60360] <= 8'h10 ;
			data[60361] <= 8'h10 ;
			data[60362] <= 8'h10 ;
			data[60363] <= 8'h10 ;
			data[60364] <= 8'h10 ;
			data[60365] <= 8'h10 ;
			data[60366] <= 8'h10 ;
			data[60367] <= 8'h10 ;
			data[60368] <= 8'h10 ;
			data[60369] <= 8'h10 ;
			data[60370] <= 8'h10 ;
			data[60371] <= 8'h10 ;
			data[60372] <= 8'h10 ;
			data[60373] <= 8'h10 ;
			data[60374] <= 8'h10 ;
			data[60375] <= 8'h10 ;
			data[60376] <= 8'h10 ;
			data[60377] <= 8'h10 ;
			data[60378] <= 8'h10 ;
			data[60379] <= 8'h10 ;
			data[60380] <= 8'h10 ;
			data[60381] <= 8'h10 ;
			data[60382] <= 8'h10 ;
			data[60383] <= 8'h10 ;
			data[60384] <= 8'h10 ;
			data[60385] <= 8'h10 ;
			data[60386] <= 8'h10 ;
			data[60387] <= 8'h10 ;
			data[60388] <= 8'h10 ;
			data[60389] <= 8'h10 ;
			data[60390] <= 8'h10 ;
			data[60391] <= 8'h10 ;
			data[60392] <= 8'h10 ;
			data[60393] <= 8'h10 ;
			data[60394] <= 8'h10 ;
			data[60395] <= 8'h10 ;
			data[60396] <= 8'h10 ;
			data[60397] <= 8'h10 ;
			data[60398] <= 8'h10 ;
			data[60399] <= 8'h10 ;
			data[60400] <= 8'h10 ;
			data[60401] <= 8'h10 ;
			data[60402] <= 8'h10 ;
			data[60403] <= 8'h10 ;
			data[60404] <= 8'h10 ;
			data[60405] <= 8'h10 ;
			data[60406] <= 8'h10 ;
			data[60407] <= 8'h10 ;
			data[60408] <= 8'h10 ;
			data[60409] <= 8'h10 ;
			data[60410] <= 8'h10 ;
			data[60411] <= 8'h10 ;
			data[60412] <= 8'h10 ;
			data[60413] <= 8'h10 ;
			data[60414] <= 8'h10 ;
			data[60415] <= 8'h10 ;
			data[60416] <= 8'h10 ;
			data[60417] <= 8'h10 ;
			data[60418] <= 8'h10 ;
			data[60419] <= 8'h10 ;
			data[60420] <= 8'h10 ;
			data[60421] <= 8'h10 ;
			data[60422] <= 8'h10 ;
			data[60423] <= 8'h10 ;
			data[60424] <= 8'h10 ;
			data[60425] <= 8'h10 ;
			data[60426] <= 8'h10 ;
			data[60427] <= 8'h10 ;
			data[60428] <= 8'h10 ;
			data[60429] <= 8'h10 ;
			data[60430] <= 8'h10 ;
			data[60431] <= 8'h10 ;
			data[60432] <= 8'h10 ;
			data[60433] <= 8'h10 ;
			data[60434] <= 8'h10 ;
			data[60435] <= 8'h10 ;
			data[60436] <= 8'h10 ;
			data[60437] <= 8'h10 ;
			data[60438] <= 8'h10 ;
			data[60439] <= 8'h10 ;
			data[60440] <= 8'h10 ;
			data[60441] <= 8'h10 ;
			data[60442] <= 8'h10 ;
			data[60443] <= 8'h10 ;
			data[60444] <= 8'h10 ;
			data[60445] <= 8'h10 ;
			data[60446] <= 8'h10 ;
			data[60447] <= 8'h10 ;
			data[60448] <= 8'h10 ;
			data[60449] <= 8'h10 ;
			data[60450] <= 8'h10 ;
			data[60451] <= 8'h10 ;
			data[60452] <= 8'h10 ;
			data[60453] <= 8'h10 ;
			data[60454] <= 8'h10 ;
			data[60455] <= 8'h10 ;
			data[60456] <= 8'h10 ;
			data[60457] <= 8'h10 ;
			data[60458] <= 8'h10 ;
			data[60459] <= 8'h10 ;
			data[60460] <= 8'h10 ;
			data[60461] <= 8'h10 ;
			data[60462] <= 8'h10 ;
			data[60463] <= 8'h10 ;
			data[60464] <= 8'h10 ;
			data[60465] <= 8'h10 ;
			data[60466] <= 8'h10 ;
			data[60467] <= 8'h10 ;
			data[60468] <= 8'h10 ;
			data[60469] <= 8'h10 ;
			data[60470] <= 8'h10 ;
			data[60471] <= 8'h10 ;
			data[60472] <= 8'h10 ;
			data[60473] <= 8'h10 ;
			data[60474] <= 8'h10 ;
			data[60475] <= 8'h10 ;
			data[60476] <= 8'h10 ;
			data[60477] <= 8'h10 ;
			data[60478] <= 8'h10 ;
			data[60479] <= 8'h10 ;
			data[60480] <= 8'h10 ;
			data[60481] <= 8'h10 ;
			data[60482] <= 8'h10 ;
			data[60483] <= 8'h10 ;
			data[60484] <= 8'h10 ;
			data[60485] <= 8'h10 ;
			data[60486] <= 8'h10 ;
			data[60487] <= 8'h10 ;
			data[60488] <= 8'h10 ;
			data[60489] <= 8'h10 ;
			data[60490] <= 8'h10 ;
			data[60491] <= 8'h10 ;
			data[60492] <= 8'h10 ;
			data[60493] <= 8'h10 ;
			data[60494] <= 8'h10 ;
			data[60495] <= 8'h10 ;
			data[60496] <= 8'h10 ;
			data[60497] <= 8'h10 ;
			data[60498] <= 8'h10 ;
			data[60499] <= 8'h10 ;
			data[60500] <= 8'h10 ;
			data[60501] <= 8'h10 ;
			data[60502] <= 8'h10 ;
			data[60503] <= 8'h10 ;
			data[60504] <= 8'h10 ;
			data[60505] <= 8'h10 ;
			data[60506] <= 8'h10 ;
			data[60507] <= 8'h10 ;
			data[60508] <= 8'h10 ;
			data[60509] <= 8'h10 ;
			data[60510] <= 8'h10 ;
			data[60511] <= 8'h10 ;
			data[60512] <= 8'h10 ;
			data[60513] <= 8'h10 ;
			data[60514] <= 8'h10 ;
			data[60515] <= 8'h10 ;
			data[60516] <= 8'h10 ;
			data[60517] <= 8'h10 ;
			data[60518] <= 8'h10 ;
			data[60519] <= 8'h10 ;
			data[60520] <= 8'h10 ;
			data[60521] <= 8'h10 ;
			data[60522] <= 8'h10 ;
			data[60523] <= 8'h10 ;
			data[60524] <= 8'h10 ;
			data[60525] <= 8'h10 ;
			data[60526] <= 8'h10 ;
			data[60527] <= 8'h10 ;
			data[60528] <= 8'h10 ;
			data[60529] <= 8'h10 ;
			data[60530] <= 8'h10 ;
			data[60531] <= 8'h10 ;
			data[60532] <= 8'h10 ;
			data[60533] <= 8'h10 ;
			data[60534] <= 8'h10 ;
			data[60535] <= 8'h10 ;
			data[60536] <= 8'h10 ;
			data[60537] <= 8'h10 ;
			data[60538] <= 8'h10 ;
			data[60539] <= 8'h10 ;
			data[60540] <= 8'h10 ;
			data[60541] <= 8'h10 ;
			data[60542] <= 8'h10 ;
			data[60543] <= 8'h10 ;
			data[60544] <= 8'h10 ;
			data[60545] <= 8'h10 ;
			data[60546] <= 8'h10 ;
			data[60547] <= 8'h10 ;
			data[60548] <= 8'h10 ;
			data[60549] <= 8'h10 ;
			data[60550] <= 8'h10 ;
			data[60551] <= 8'h10 ;
			data[60552] <= 8'h10 ;
			data[60553] <= 8'h10 ;
			data[60554] <= 8'h10 ;
			data[60555] <= 8'h10 ;
			data[60556] <= 8'h10 ;
			data[60557] <= 8'h10 ;
			data[60558] <= 8'h10 ;
			data[60559] <= 8'h10 ;
			data[60560] <= 8'h10 ;
			data[60561] <= 8'h10 ;
			data[60562] <= 8'h10 ;
			data[60563] <= 8'h10 ;
			data[60564] <= 8'h10 ;
			data[60565] <= 8'h10 ;
			data[60566] <= 8'h10 ;
			data[60567] <= 8'h10 ;
			data[60568] <= 8'h10 ;
			data[60569] <= 8'h10 ;
			data[60570] <= 8'h10 ;
			data[60571] <= 8'h10 ;
			data[60572] <= 8'h10 ;
			data[60573] <= 8'h10 ;
			data[60574] <= 8'h10 ;
			data[60575] <= 8'h10 ;
			data[60576] <= 8'h10 ;
			data[60577] <= 8'h10 ;
			data[60578] <= 8'h10 ;
			data[60579] <= 8'h10 ;
			data[60580] <= 8'h10 ;
			data[60581] <= 8'h10 ;
			data[60582] <= 8'h10 ;
			data[60583] <= 8'h10 ;
			data[60584] <= 8'h10 ;
			data[60585] <= 8'h10 ;
			data[60586] <= 8'h10 ;
			data[60587] <= 8'h10 ;
			data[60588] <= 8'h10 ;
			data[60589] <= 8'h10 ;
			data[60590] <= 8'h10 ;
			data[60591] <= 8'h10 ;
			data[60592] <= 8'h10 ;
			data[60593] <= 8'h10 ;
			data[60594] <= 8'h10 ;
			data[60595] <= 8'h10 ;
			data[60596] <= 8'h10 ;
			data[60597] <= 8'h10 ;
			data[60598] <= 8'h10 ;
			data[60599] <= 8'h10 ;
			data[60600] <= 8'h10 ;
			data[60601] <= 8'h10 ;
			data[60602] <= 8'h10 ;
			data[60603] <= 8'h10 ;
			data[60604] <= 8'h10 ;
			data[60605] <= 8'h10 ;
			data[60606] <= 8'h10 ;
			data[60607] <= 8'h10 ;
			data[60608] <= 8'h10 ;
			data[60609] <= 8'h10 ;
			data[60610] <= 8'h10 ;
			data[60611] <= 8'h10 ;
			data[60612] <= 8'h10 ;
			data[60613] <= 8'h10 ;
			data[60614] <= 8'h10 ;
			data[60615] <= 8'h10 ;
			data[60616] <= 8'h10 ;
			data[60617] <= 8'h10 ;
			data[60618] <= 8'h10 ;
			data[60619] <= 8'h10 ;
			data[60620] <= 8'h10 ;
			data[60621] <= 8'h10 ;
			data[60622] <= 8'h10 ;
			data[60623] <= 8'h10 ;
			data[60624] <= 8'h10 ;
			data[60625] <= 8'h10 ;
			data[60626] <= 8'h10 ;
			data[60627] <= 8'h10 ;
			data[60628] <= 8'h10 ;
			data[60629] <= 8'h10 ;
			data[60630] <= 8'h10 ;
			data[60631] <= 8'h10 ;
			data[60632] <= 8'h10 ;
			data[60633] <= 8'h10 ;
			data[60634] <= 8'h10 ;
			data[60635] <= 8'h10 ;
			data[60636] <= 8'h10 ;
			data[60637] <= 8'h10 ;
			data[60638] <= 8'h10 ;
			data[60639] <= 8'h10 ;
			data[60640] <= 8'h10 ;
			data[60641] <= 8'h10 ;
			data[60642] <= 8'h10 ;
			data[60643] <= 8'h10 ;
			data[60644] <= 8'h10 ;
			data[60645] <= 8'h10 ;
			data[60646] <= 8'h10 ;
			data[60647] <= 8'h10 ;
			data[60648] <= 8'h10 ;
			data[60649] <= 8'h10 ;
			data[60650] <= 8'h10 ;
			data[60651] <= 8'h10 ;
			data[60652] <= 8'h10 ;
			data[60653] <= 8'h10 ;
			data[60654] <= 8'h10 ;
			data[60655] <= 8'h10 ;
			data[60656] <= 8'h10 ;
			data[60657] <= 8'h10 ;
			data[60658] <= 8'h10 ;
			data[60659] <= 8'h10 ;
			data[60660] <= 8'h10 ;
			data[60661] <= 8'h10 ;
			data[60662] <= 8'h10 ;
			data[60663] <= 8'h10 ;
			data[60664] <= 8'h10 ;
			data[60665] <= 8'h10 ;
			data[60666] <= 8'h10 ;
			data[60667] <= 8'h10 ;
			data[60668] <= 8'h10 ;
			data[60669] <= 8'h10 ;
			data[60670] <= 8'h10 ;
			data[60671] <= 8'h10 ;
			data[60672] <= 8'h10 ;
			data[60673] <= 8'h10 ;
			data[60674] <= 8'h10 ;
			data[60675] <= 8'h10 ;
			data[60676] <= 8'h10 ;
			data[60677] <= 8'h10 ;
			data[60678] <= 8'h10 ;
			data[60679] <= 8'h10 ;
			data[60680] <= 8'h10 ;
			data[60681] <= 8'h10 ;
			data[60682] <= 8'h10 ;
			data[60683] <= 8'h10 ;
			data[60684] <= 8'h10 ;
			data[60685] <= 8'h10 ;
			data[60686] <= 8'h10 ;
			data[60687] <= 8'h10 ;
			data[60688] <= 8'h10 ;
			data[60689] <= 8'h10 ;
			data[60690] <= 8'h10 ;
			data[60691] <= 8'h10 ;
			data[60692] <= 8'h10 ;
			data[60693] <= 8'h10 ;
			data[60694] <= 8'h10 ;
			data[60695] <= 8'h10 ;
			data[60696] <= 8'h10 ;
			data[60697] <= 8'h10 ;
			data[60698] <= 8'h10 ;
			data[60699] <= 8'h10 ;
			data[60700] <= 8'h10 ;
			data[60701] <= 8'h10 ;
			data[60702] <= 8'h10 ;
			data[60703] <= 8'h10 ;
			data[60704] <= 8'h10 ;
			data[60705] <= 8'h10 ;
			data[60706] <= 8'h10 ;
			data[60707] <= 8'h10 ;
			data[60708] <= 8'h10 ;
			data[60709] <= 8'h10 ;
			data[60710] <= 8'h10 ;
			data[60711] <= 8'h10 ;
			data[60712] <= 8'h10 ;
			data[60713] <= 8'h10 ;
			data[60714] <= 8'h10 ;
			data[60715] <= 8'h10 ;
			data[60716] <= 8'h10 ;
			data[60717] <= 8'h10 ;
			data[60718] <= 8'h10 ;
			data[60719] <= 8'h10 ;
			data[60720] <= 8'h10 ;
			data[60721] <= 8'h10 ;
			data[60722] <= 8'h10 ;
			data[60723] <= 8'h10 ;
			data[60724] <= 8'h10 ;
			data[60725] <= 8'h10 ;
			data[60726] <= 8'h10 ;
			data[60727] <= 8'h10 ;
			data[60728] <= 8'h10 ;
			data[60729] <= 8'h10 ;
			data[60730] <= 8'h10 ;
			data[60731] <= 8'h10 ;
			data[60732] <= 8'h10 ;
			data[60733] <= 8'h10 ;
			data[60734] <= 8'h10 ;
			data[60735] <= 8'h10 ;
			data[60736] <= 8'h10 ;
			data[60737] <= 8'h10 ;
			data[60738] <= 8'h10 ;
			data[60739] <= 8'h10 ;
			data[60740] <= 8'h10 ;
			data[60741] <= 8'h10 ;
			data[60742] <= 8'h10 ;
			data[60743] <= 8'h10 ;
			data[60744] <= 8'h10 ;
			data[60745] <= 8'h10 ;
			data[60746] <= 8'h10 ;
			data[60747] <= 8'h10 ;
			data[60748] <= 8'h10 ;
			data[60749] <= 8'h10 ;
			data[60750] <= 8'h10 ;
			data[60751] <= 8'h10 ;
			data[60752] <= 8'h10 ;
			data[60753] <= 8'h10 ;
			data[60754] <= 8'h10 ;
			data[60755] <= 8'h10 ;
			data[60756] <= 8'h10 ;
			data[60757] <= 8'h10 ;
			data[60758] <= 8'h10 ;
			data[60759] <= 8'h10 ;
			data[60760] <= 8'h10 ;
			data[60761] <= 8'h10 ;
			data[60762] <= 8'h10 ;
			data[60763] <= 8'h10 ;
			data[60764] <= 8'h10 ;
			data[60765] <= 8'h10 ;
			data[60766] <= 8'h10 ;
			data[60767] <= 8'h10 ;
			data[60768] <= 8'h10 ;
			data[60769] <= 8'h10 ;
			data[60770] <= 8'h10 ;
			data[60771] <= 8'h10 ;
			data[60772] <= 8'h10 ;
			data[60773] <= 8'h10 ;
			data[60774] <= 8'h10 ;
			data[60775] <= 8'h10 ;
			data[60776] <= 8'h10 ;
			data[60777] <= 8'h10 ;
			data[60778] <= 8'h10 ;
			data[60779] <= 8'h10 ;
			data[60780] <= 8'h10 ;
			data[60781] <= 8'h10 ;
			data[60782] <= 8'h10 ;
			data[60783] <= 8'h10 ;
			data[60784] <= 8'h10 ;
			data[60785] <= 8'h10 ;
			data[60786] <= 8'h10 ;
			data[60787] <= 8'h10 ;
			data[60788] <= 8'h10 ;
			data[60789] <= 8'h10 ;
			data[60790] <= 8'h10 ;
			data[60791] <= 8'h10 ;
			data[60792] <= 8'h10 ;
			data[60793] <= 8'h10 ;
			data[60794] <= 8'h10 ;
			data[60795] <= 8'h10 ;
			data[60796] <= 8'h10 ;
			data[60797] <= 8'h10 ;
			data[60798] <= 8'h10 ;
			data[60799] <= 8'h10 ;
			data[60800] <= 8'h10 ;
			data[60801] <= 8'h10 ;
			data[60802] <= 8'h10 ;
			data[60803] <= 8'h10 ;
			data[60804] <= 8'h10 ;
			data[60805] <= 8'h10 ;
			data[60806] <= 8'h10 ;
			data[60807] <= 8'h10 ;
			data[60808] <= 8'h10 ;
			data[60809] <= 8'h10 ;
			data[60810] <= 8'h10 ;
			data[60811] <= 8'h10 ;
			data[60812] <= 8'h10 ;
			data[60813] <= 8'h10 ;
			data[60814] <= 8'h10 ;
			data[60815] <= 8'h10 ;
			data[60816] <= 8'h10 ;
			data[60817] <= 8'h10 ;
			data[60818] <= 8'h10 ;
			data[60819] <= 8'h10 ;
			data[60820] <= 8'h10 ;
			data[60821] <= 8'h10 ;
			data[60822] <= 8'h10 ;
			data[60823] <= 8'h10 ;
			data[60824] <= 8'h10 ;
			data[60825] <= 8'h10 ;
			data[60826] <= 8'h10 ;
			data[60827] <= 8'h10 ;
			data[60828] <= 8'h10 ;
			data[60829] <= 8'h10 ;
			data[60830] <= 8'h10 ;
			data[60831] <= 8'h10 ;
			data[60832] <= 8'h10 ;
			data[60833] <= 8'h10 ;
			data[60834] <= 8'h10 ;
			data[60835] <= 8'h10 ;
			data[60836] <= 8'h10 ;
			data[60837] <= 8'h10 ;
			data[60838] <= 8'h10 ;
			data[60839] <= 8'h10 ;
			data[60840] <= 8'h10 ;
			data[60841] <= 8'h10 ;
			data[60842] <= 8'h10 ;
			data[60843] <= 8'h10 ;
			data[60844] <= 8'h10 ;
			data[60845] <= 8'h10 ;
			data[60846] <= 8'h10 ;
			data[60847] <= 8'h10 ;
			data[60848] <= 8'h10 ;
			data[60849] <= 8'h10 ;
			data[60850] <= 8'h10 ;
			data[60851] <= 8'h10 ;
			data[60852] <= 8'h10 ;
			data[60853] <= 8'h10 ;
			data[60854] <= 8'h10 ;
			data[60855] <= 8'h10 ;
			data[60856] <= 8'h10 ;
			data[60857] <= 8'h10 ;
			data[60858] <= 8'h10 ;
			data[60859] <= 8'h10 ;
			data[60860] <= 8'h10 ;
			data[60861] <= 8'h10 ;
			data[60862] <= 8'h10 ;
			data[60863] <= 8'h10 ;
			data[60864] <= 8'h10 ;
			data[60865] <= 8'h10 ;
			data[60866] <= 8'h10 ;
			data[60867] <= 8'h10 ;
			data[60868] <= 8'h10 ;
			data[60869] <= 8'h10 ;
			data[60870] <= 8'h10 ;
			data[60871] <= 8'h10 ;
			data[60872] <= 8'h10 ;
			data[60873] <= 8'h10 ;
			data[60874] <= 8'h10 ;
			data[60875] <= 8'h10 ;
			data[60876] <= 8'h10 ;
			data[60877] <= 8'h10 ;
			data[60878] <= 8'h10 ;
			data[60879] <= 8'h10 ;
			data[60880] <= 8'h10 ;
			data[60881] <= 8'h10 ;
			data[60882] <= 8'h10 ;
			data[60883] <= 8'h10 ;
			data[60884] <= 8'h10 ;
			data[60885] <= 8'h10 ;
			data[60886] <= 8'h10 ;
			data[60887] <= 8'h10 ;
			data[60888] <= 8'h10 ;
			data[60889] <= 8'h10 ;
			data[60890] <= 8'h10 ;
			data[60891] <= 8'h10 ;
			data[60892] <= 8'h10 ;
			data[60893] <= 8'h10 ;
			data[60894] <= 8'h10 ;
			data[60895] <= 8'h10 ;
			data[60896] <= 8'h10 ;
			data[60897] <= 8'h10 ;
			data[60898] <= 8'h10 ;
			data[60899] <= 8'h10 ;
			data[60900] <= 8'h10 ;
			data[60901] <= 8'h10 ;
			data[60902] <= 8'h10 ;
			data[60903] <= 8'h10 ;
			data[60904] <= 8'h10 ;
			data[60905] <= 8'h10 ;
			data[60906] <= 8'h10 ;
			data[60907] <= 8'h10 ;
			data[60908] <= 8'h10 ;
			data[60909] <= 8'h10 ;
			data[60910] <= 8'h10 ;
			data[60911] <= 8'h10 ;
			data[60912] <= 8'h10 ;
			data[60913] <= 8'h10 ;
			data[60914] <= 8'h10 ;
			data[60915] <= 8'h10 ;
			data[60916] <= 8'h10 ;
			data[60917] <= 8'h10 ;
			data[60918] <= 8'h10 ;
			data[60919] <= 8'h10 ;
			data[60920] <= 8'h10 ;
			data[60921] <= 8'h10 ;
			data[60922] <= 8'h10 ;
			data[60923] <= 8'h10 ;
			data[60924] <= 8'h10 ;
			data[60925] <= 8'h10 ;
			data[60926] <= 8'h10 ;
			data[60927] <= 8'h10 ;
			data[60928] <= 8'h10 ;
			data[60929] <= 8'h10 ;
			data[60930] <= 8'h10 ;
			data[60931] <= 8'h10 ;
			data[60932] <= 8'h10 ;
			data[60933] <= 8'h10 ;
			data[60934] <= 8'h10 ;
			data[60935] <= 8'h10 ;
			data[60936] <= 8'h10 ;
			data[60937] <= 8'h10 ;
			data[60938] <= 8'h10 ;
			data[60939] <= 8'h10 ;
			data[60940] <= 8'h10 ;
			data[60941] <= 8'h10 ;
			data[60942] <= 8'h10 ;
			data[60943] <= 8'h10 ;
			data[60944] <= 8'h10 ;
			data[60945] <= 8'h10 ;
			data[60946] <= 8'h10 ;
			data[60947] <= 8'h10 ;
			data[60948] <= 8'h10 ;
			data[60949] <= 8'h10 ;
			data[60950] <= 8'h10 ;
			data[60951] <= 8'h10 ;
			data[60952] <= 8'h10 ;
			data[60953] <= 8'h10 ;
			data[60954] <= 8'h10 ;
			data[60955] <= 8'h10 ;
			data[60956] <= 8'h10 ;
			data[60957] <= 8'h10 ;
			data[60958] <= 8'h10 ;
			data[60959] <= 8'h10 ;
			data[60960] <= 8'h10 ;
			data[60961] <= 8'h10 ;
			data[60962] <= 8'h10 ;
			data[60963] <= 8'h10 ;
			data[60964] <= 8'h10 ;
			data[60965] <= 8'h10 ;
			data[60966] <= 8'h10 ;
			data[60967] <= 8'h10 ;
			data[60968] <= 8'h10 ;
			data[60969] <= 8'h10 ;
			data[60970] <= 8'h10 ;
			data[60971] <= 8'h10 ;
			data[60972] <= 8'h10 ;
			data[60973] <= 8'h10 ;
			data[60974] <= 8'h10 ;
			data[60975] <= 8'h10 ;
			data[60976] <= 8'h10 ;
			data[60977] <= 8'h10 ;
			data[60978] <= 8'h10 ;
			data[60979] <= 8'h10 ;
			data[60980] <= 8'h10 ;
			data[60981] <= 8'h10 ;
			data[60982] <= 8'h10 ;
			data[60983] <= 8'h10 ;
			data[60984] <= 8'h10 ;
			data[60985] <= 8'h10 ;
			data[60986] <= 8'h10 ;
			data[60987] <= 8'h10 ;
			data[60988] <= 8'h10 ;
			data[60989] <= 8'h10 ;
			data[60990] <= 8'h10 ;
			data[60991] <= 8'h10 ;
			data[60992] <= 8'h10 ;
			data[60993] <= 8'h10 ;
			data[60994] <= 8'h10 ;
			data[60995] <= 8'h10 ;
			data[60996] <= 8'h10 ;
			data[60997] <= 8'h10 ;
			data[60998] <= 8'h10 ;
			data[60999] <= 8'h10 ;
			data[61000] <= 8'h10 ;
			data[61001] <= 8'h10 ;
			data[61002] <= 8'h10 ;
			data[61003] <= 8'h10 ;
			data[61004] <= 8'h10 ;
			data[61005] <= 8'h10 ;
			data[61006] <= 8'h10 ;
			data[61007] <= 8'h10 ;
			data[61008] <= 8'h10 ;
			data[61009] <= 8'h10 ;
			data[61010] <= 8'h10 ;
			data[61011] <= 8'h10 ;
			data[61012] <= 8'h10 ;
			data[61013] <= 8'h10 ;
			data[61014] <= 8'h10 ;
			data[61015] <= 8'h10 ;
			data[61016] <= 8'h10 ;
			data[61017] <= 8'h10 ;
			data[61018] <= 8'h10 ;
			data[61019] <= 8'h10 ;
			data[61020] <= 8'h10 ;
			data[61021] <= 8'h10 ;
			data[61022] <= 8'h10 ;
			data[61023] <= 8'h10 ;
			data[61024] <= 8'h10 ;
			data[61025] <= 8'h10 ;
			data[61026] <= 8'h10 ;
			data[61027] <= 8'h10 ;
			data[61028] <= 8'h10 ;
			data[61029] <= 8'h10 ;
			data[61030] <= 8'h10 ;
			data[61031] <= 8'h10 ;
			data[61032] <= 8'h10 ;
			data[61033] <= 8'h10 ;
			data[61034] <= 8'h10 ;
			data[61035] <= 8'h10 ;
			data[61036] <= 8'h10 ;
			data[61037] <= 8'h10 ;
			data[61038] <= 8'h10 ;
			data[61039] <= 8'h10 ;
			data[61040] <= 8'h10 ;
			data[61041] <= 8'h10 ;
			data[61042] <= 8'h10 ;
			data[61043] <= 8'h10 ;
			data[61044] <= 8'h10 ;
			data[61045] <= 8'h10 ;
			data[61046] <= 8'h10 ;
			data[61047] <= 8'h10 ;
			data[61048] <= 8'h10 ;
			data[61049] <= 8'h10 ;
			data[61050] <= 8'h10 ;
			data[61051] <= 8'h10 ;
			data[61052] <= 8'h10 ;
			data[61053] <= 8'h10 ;
			data[61054] <= 8'h10 ;
			data[61055] <= 8'h10 ;
			data[61056] <= 8'h10 ;
			data[61057] <= 8'h10 ;
			data[61058] <= 8'h10 ;
			data[61059] <= 8'h10 ;
			data[61060] <= 8'h10 ;
			data[61061] <= 8'h10 ;
			data[61062] <= 8'h10 ;
			data[61063] <= 8'h10 ;
			data[61064] <= 8'h10 ;
			data[61065] <= 8'h10 ;
			data[61066] <= 8'h10 ;
			data[61067] <= 8'h10 ;
			data[61068] <= 8'h10 ;
			data[61069] <= 8'h10 ;
			data[61070] <= 8'h10 ;
			data[61071] <= 8'h10 ;
			data[61072] <= 8'h10 ;
			data[61073] <= 8'h10 ;
			data[61074] <= 8'h10 ;
			data[61075] <= 8'h10 ;
			data[61076] <= 8'h10 ;
			data[61077] <= 8'h10 ;
			data[61078] <= 8'h10 ;
			data[61079] <= 8'h10 ;
			data[61080] <= 8'h10 ;
			data[61081] <= 8'h10 ;
			data[61082] <= 8'h10 ;
			data[61083] <= 8'h10 ;
			data[61084] <= 8'h10 ;
			data[61085] <= 8'h10 ;
			data[61086] <= 8'h10 ;
			data[61087] <= 8'h10 ;
			data[61088] <= 8'h10 ;
			data[61089] <= 8'h10 ;
			data[61090] <= 8'h10 ;
			data[61091] <= 8'h10 ;
			data[61092] <= 8'h10 ;
			data[61093] <= 8'h10 ;
			data[61094] <= 8'h10 ;
			data[61095] <= 8'h10 ;
			data[61096] <= 8'h10 ;
			data[61097] <= 8'h10 ;
			data[61098] <= 8'h10 ;
			data[61099] <= 8'h10 ;
			data[61100] <= 8'h10 ;
			data[61101] <= 8'h10 ;
			data[61102] <= 8'h10 ;
			data[61103] <= 8'h10 ;
			data[61104] <= 8'h10 ;
			data[61105] <= 8'h10 ;
			data[61106] <= 8'h10 ;
			data[61107] <= 8'h10 ;
			data[61108] <= 8'h10 ;
			data[61109] <= 8'h10 ;
			data[61110] <= 8'h10 ;
			data[61111] <= 8'h10 ;
			data[61112] <= 8'h10 ;
			data[61113] <= 8'h10 ;
			data[61114] <= 8'h10 ;
			data[61115] <= 8'h10 ;
			data[61116] <= 8'h10 ;
			data[61117] <= 8'h10 ;
			data[61118] <= 8'h10 ;
			data[61119] <= 8'h10 ;
			data[61120] <= 8'h10 ;
			data[61121] <= 8'h10 ;
			data[61122] <= 8'h10 ;
			data[61123] <= 8'h10 ;
			data[61124] <= 8'h10 ;
			data[61125] <= 8'h10 ;
			data[61126] <= 8'h10 ;
			data[61127] <= 8'h10 ;
			data[61128] <= 8'h10 ;
			data[61129] <= 8'h10 ;
			data[61130] <= 8'h10 ;
			data[61131] <= 8'h10 ;
			data[61132] <= 8'h10 ;
			data[61133] <= 8'h10 ;
			data[61134] <= 8'h10 ;
			data[61135] <= 8'h10 ;
			data[61136] <= 8'h10 ;
			data[61137] <= 8'h10 ;
			data[61138] <= 8'h10 ;
			data[61139] <= 8'h10 ;
			data[61140] <= 8'h10 ;
			data[61141] <= 8'h10 ;
			data[61142] <= 8'h10 ;
			data[61143] <= 8'h10 ;
			data[61144] <= 8'h10 ;
			data[61145] <= 8'h10 ;
			data[61146] <= 8'h10 ;
			data[61147] <= 8'h10 ;
			data[61148] <= 8'h10 ;
			data[61149] <= 8'h10 ;
			data[61150] <= 8'h10 ;
			data[61151] <= 8'h10 ;
			data[61152] <= 8'h10 ;
			data[61153] <= 8'h10 ;
			data[61154] <= 8'h10 ;
			data[61155] <= 8'h10 ;
			data[61156] <= 8'h10 ;
			data[61157] <= 8'h10 ;
			data[61158] <= 8'h10 ;
			data[61159] <= 8'h10 ;
			data[61160] <= 8'h10 ;
			data[61161] <= 8'h10 ;
			data[61162] <= 8'h10 ;
			data[61163] <= 8'h10 ;
			data[61164] <= 8'h10 ;
			data[61165] <= 8'h10 ;
			data[61166] <= 8'h10 ;
			data[61167] <= 8'h10 ;
			data[61168] <= 8'h10 ;
			data[61169] <= 8'h10 ;
			data[61170] <= 8'h10 ;
			data[61171] <= 8'h10 ;
			data[61172] <= 8'h10 ;
			data[61173] <= 8'h10 ;
			data[61174] <= 8'h10 ;
			data[61175] <= 8'h10 ;
			data[61176] <= 8'h10 ;
			data[61177] <= 8'h10 ;
			data[61178] <= 8'h10 ;
			data[61179] <= 8'h10 ;
			data[61180] <= 8'h10 ;
			data[61181] <= 8'h10 ;
			data[61182] <= 8'h10 ;
			data[61183] <= 8'h10 ;
			data[61184] <= 8'h10 ;
			data[61185] <= 8'h10 ;
			data[61186] <= 8'h10 ;
			data[61187] <= 8'h10 ;
			data[61188] <= 8'h10 ;
			data[61189] <= 8'h10 ;
			data[61190] <= 8'h10 ;
			data[61191] <= 8'h10 ;
			data[61192] <= 8'h10 ;
			data[61193] <= 8'h10 ;
			data[61194] <= 8'h10 ;
			data[61195] <= 8'h10 ;
			data[61196] <= 8'h10 ;
			data[61197] <= 8'h10 ;
			data[61198] <= 8'h10 ;
			data[61199] <= 8'h10 ;
			data[61200] <= 8'h10 ;
			data[61201] <= 8'h10 ;
			data[61202] <= 8'h10 ;
			data[61203] <= 8'h10 ;
			data[61204] <= 8'h10 ;
			data[61205] <= 8'h10 ;
			data[61206] <= 8'h10 ;
			data[61207] <= 8'h10 ;
			data[61208] <= 8'h10 ;
			data[61209] <= 8'h10 ;
			data[61210] <= 8'h10 ;
			data[61211] <= 8'h10 ;
			data[61212] <= 8'h10 ;
			data[61213] <= 8'h10 ;
			data[61214] <= 8'h10 ;
			data[61215] <= 8'h10 ;
			data[61216] <= 8'h10 ;
			data[61217] <= 8'h10 ;
			data[61218] <= 8'h10 ;
			data[61219] <= 8'h10 ;
			data[61220] <= 8'h10 ;
			data[61221] <= 8'h10 ;
			data[61222] <= 8'h10 ;
			data[61223] <= 8'h10 ;
			data[61224] <= 8'h10 ;
			data[61225] <= 8'h10 ;
			data[61226] <= 8'h10 ;
			data[61227] <= 8'h10 ;
			data[61228] <= 8'h10 ;
			data[61229] <= 8'h10 ;
			data[61230] <= 8'h10 ;
			data[61231] <= 8'h10 ;
			data[61232] <= 8'h10 ;
			data[61233] <= 8'h10 ;
			data[61234] <= 8'h10 ;
			data[61235] <= 8'h10 ;
			data[61236] <= 8'h10 ;
			data[61237] <= 8'h10 ;
			data[61238] <= 8'h10 ;
			data[61239] <= 8'h10 ;
			data[61240] <= 8'h10 ;
			data[61241] <= 8'h10 ;
			data[61242] <= 8'h10 ;
			data[61243] <= 8'h10 ;
			data[61244] <= 8'h10 ;
			data[61245] <= 8'h10 ;
			data[61246] <= 8'h10 ;
			data[61247] <= 8'h10 ;
			data[61248] <= 8'h10 ;
			data[61249] <= 8'h10 ;
			data[61250] <= 8'h10 ;
			data[61251] <= 8'h10 ;
			data[61252] <= 8'h10 ;
			data[61253] <= 8'h10 ;
			data[61254] <= 8'h10 ;
			data[61255] <= 8'h10 ;
			data[61256] <= 8'h10 ;
			data[61257] <= 8'h10 ;
			data[61258] <= 8'h10 ;
			data[61259] <= 8'h10 ;
			data[61260] <= 8'h10 ;
			data[61261] <= 8'h10 ;
			data[61262] <= 8'h10 ;
			data[61263] <= 8'h10 ;
			data[61264] <= 8'h10 ;
			data[61265] <= 8'h10 ;
			data[61266] <= 8'h10 ;
			data[61267] <= 8'h10 ;
			data[61268] <= 8'h10 ;
			data[61269] <= 8'h10 ;
			data[61270] <= 8'h10 ;
			data[61271] <= 8'h10 ;
			data[61272] <= 8'h10 ;
			data[61273] <= 8'h10 ;
			data[61274] <= 8'h10 ;
			data[61275] <= 8'h10 ;
			data[61276] <= 8'h10 ;
			data[61277] <= 8'h10 ;
			data[61278] <= 8'h10 ;
			data[61279] <= 8'h10 ;
			data[61280] <= 8'h10 ;
			data[61281] <= 8'h10 ;
			data[61282] <= 8'h10 ;
			data[61283] <= 8'h10 ;
			data[61284] <= 8'h10 ;
			data[61285] <= 8'h10 ;
			data[61286] <= 8'h10 ;
			data[61287] <= 8'h10 ;
			data[61288] <= 8'h10 ;
			data[61289] <= 8'h10 ;
			data[61290] <= 8'h10 ;
			data[61291] <= 8'h10 ;
			data[61292] <= 8'h10 ;
			data[61293] <= 8'h10 ;
			data[61294] <= 8'h10 ;
			data[61295] <= 8'h10 ;
			data[61296] <= 8'h10 ;
			data[61297] <= 8'h10 ;
			data[61298] <= 8'h10 ;
			data[61299] <= 8'h10 ;
			data[61300] <= 8'h10 ;
			data[61301] <= 8'h10 ;
			data[61302] <= 8'h10 ;
			data[61303] <= 8'h10 ;
			data[61304] <= 8'h10 ;
			data[61305] <= 8'h10 ;
			data[61306] <= 8'h10 ;
			data[61307] <= 8'h10 ;
			data[61308] <= 8'h10 ;
			data[61309] <= 8'h10 ;
			data[61310] <= 8'h10 ;
			data[61311] <= 8'h10 ;
			data[61312] <= 8'h10 ;
			data[61313] <= 8'h10 ;
			data[61314] <= 8'h10 ;
			data[61315] <= 8'h10 ;
			data[61316] <= 8'h10 ;
			data[61317] <= 8'h10 ;
			data[61318] <= 8'h10 ;
			data[61319] <= 8'h10 ;
			data[61320] <= 8'h10 ;
			data[61321] <= 8'h10 ;
			data[61322] <= 8'h10 ;
			data[61323] <= 8'h10 ;
			data[61324] <= 8'h10 ;
			data[61325] <= 8'h10 ;
			data[61326] <= 8'h10 ;
			data[61327] <= 8'h10 ;
			data[61328] <= 8'h10 ;
			data[61329] <= 8'h10 ;
			data[61330] <= 8'h10 ;
			data[61331] <= 8'h10 ;
			data[61332] <= 8'h10 ;
			data[61333] <= 8'h10 ;
			data[61334] <= 8'h10 ;
			data[61335] <= 8'h10 ;
			data[61336] <= 8'h10 ;
			data[61337] <= 8'h10 ;
			data[61338] <= 8'h10 ;
			data[61339] <= 8'h10 ;
			data[61340] <= 8'h10 ;
			data[61341] <= 8'h10 ;
			data[61342] <= 8'h10 ;
			data[61343] <= 8'h10 ;
			data[61344] <= 8'h10 ;
			data[61345] <= 8'h10 ;
			data[61346] <= 8'h10 ;
			data[61347] <= 8'h10 ;
			data[61348] <= 8'h10 ;
			data[61349] <= 8'h10 ;
			data[61350] <= 8'h10 ;
			data[61351] <= 8'h10 ;
			data[61352] <= 8'h10 ;
			data[61353] <= 8'h10 ;
			data[61354] <= 8'h10 ;
			data[61355] <= 8'h10 ;
			data[61356] <= 8'h10 ;
			data[61357] <= 8'h10 ;
			data[61358] <= 8'h10 ;
			data[61359] <= 8'h10 ;
			data[61360] <= 8'h10 ;
			data[61361] <= 8'h10 ;
			data[61362] <= 8'h10 ;
			data[61363] <= 8'h10 ;
			data[61364] <= 8'h10 ;
			data[61365] <= 8'h10 ;
			data[61366] <= 8'h10 ;
			data[61367] <= 8'h10 ;
			data[61368] <= 8'h10 ;
			data[61369] <= 8'h10 ;
			data[61370] <= 8'h10 ;
			data[61371] <= 8'h10 ;
			data[61372] <= 8'h10 ;
			data[61373] <= 8'h10 ;
			data[61374] <= 8'h10 ;
			data[61375] <= 8'h10 ;
			data[61376] <= 8'h10 ;
			data[61377] <= 8'h10 ;
			data[61378] <= 8'h10 ;
			data[61379] <= 8'h10 ;
			data[61380] <= 8'h10 ;
			data[61381] <= 8'h10 ;
			data[61382] <= 8'h10 ;
			data[61383] <= 8'h10 ;
			data[61384] <= 8'h10 ;
			data[61385] <= 8'h10 ;
			data[61386] <= 8'h10 ;
			data[61387] <= 8'h10 ;
			data[61388] <= 8'h10 ;
			data[61389] <= 8'h10 ;
			data[61390] <= 8'h10 ;
			data[61391] <= 8'h10 ;
			data[61392] <= 8'h10 ;
			data[61393] <= 8'h10 ;
			data[61394] <= 8'h10 ;
			data[61395] <= 8'h10 ;
			data[61396] <= 8'h10 ;
			data[61397] <= 8'h10 ;
			data[61398] <= 8'h10 ;
			data[61399] <= 8'h10 ;
			data[61400] <= 8'h10 ;
			data[61401] <= 8'h10 ;
			data[61402] <= 8'h10 ;
			data[61403] <= 8'h10 ;
			data[61404] <= 8'h10 ;
			data[61405] <= 8'h10 ;
			data[61406] <= 8'h10 ;
			data[61407] <= 8'h10 ;
			data[61408] <= 8'h10 ;
			data[61409] <= 8'h10 ;
			data[61410] <= 8'h10 ;
			data[61411] <= 8'h10 ;
			data[61412] <= 8'h10 ;
			data[61413] <= 8'h10 ;
			data[61414] <= 8'h10 ;
			data[61415] <= 8'h10 ;
			data[61416] <= 8'h10 ;
			data[61417] <= 8'h10 ;
			data[61418] <= 8'h10 ;
			data[61419] <= 8'h10 ;
			data[61420] <= 8'h10 ;
			data[61421] <= 8'h10 ;
			data[61422] <= 8'h10 ;
			data[61423] <= 8'h10 ;
			data[61424] <= 8'h10 ;
			data[61425] <= 8'h10 ;
			data[61426] <= 8'h10 ;
			data[61427] <= 8'h10 ;
			data[61428] <= 8'h10 ;
			data[61429] <= 8'h10 ;
			data[61430] <= 8'h10 ;
			data[61431] <= 8'h10 ;
			data[61432] <= 8'h10 ;
			data[61433] <= 8'h10 ;
			data[61434] <= 8'h10 ;
			data[61435] <= 8'h10 ;
			data[61436] <= 8'h10 ;
			data[61437] <= 8'h10 ;
			data[61438] <= 8'h10 ;
			data[61439] <= 8'h10 ;
			data[61440] <= 8'h10 ;
			data[61441] <= 8'h10 ;
			data[61442] <= 8'h10 ;
			data[61443] <= 8'h10 ;
			data[61444] <= 8'h10 ;
			data[61445] <= 8'h10 ;
			data[61446] <= 8'h10 ;
			data[61447] <= 8'h10 ;
			data[61448] <= 8'h10 ;
			data[61449] <= 8'h10 ;
			data[61450] <= 8'h10 ;
			data[61451] <= 8'h10 ;
			data[61452] <= 8'h10 ;
			data[61453] <= 8'h10 ;
			data[61454] <= 8'h10 ;
			data[61455] <= 8'h10 ;
			data[61456] <= 8'h10 ;
			data[61457] <= 8'h10 ;
			data[61458] <= 8'h10 ;
			data[61459] <= 8'h10 ;
			data[61460] <= 8'h10 ;
			data[61461] <= 8'h10 ;
			data[61462] <= 8'h10 ;
			data[61463] <= 8'h10 ;
			data[61464] <= 8'h10 ;
			data[61465] <= 8'h10 ;
			data[61466] <= 8'h10 ;
			data[61467] <= 8'h10 ;
			data[61468] <= 8'h10 ;
			data[61469] <= 8'h10 ;
			data[61470] <= 8'h10 ;
			data[61471] <= 8'h10 ;
			data[61472] <= 8'h10 ;
			data[61473] <= 8'h10 ;
			data[61474] <= 8'h10 ;
			data[61475] <= 8'h10 ;
			data[61476] <= 8'h10 ;
			data[61477] <= 8'h10 ;
			data[61478] <= 8'h10 ;
			data[61479] <= 8'h10 ;
			data[61480] <= 8'h10 ;
			data[61481] <= 8'h10 ;
			data[61482] <= 8'h10 ;
			data[61483] <= 8'h10 ;
			data[61484] <= 8'h10 ;
			data[61485] <= 8'h10 ;
			data[61486] <= 8'h10 ;
			data[61487] <= 8'h10 ;
			data[61488] <= 8'h10 ;
			data[61489] <= 8'h10 ;
			data[61490] <= 8'h10 ;
			data[61491] <= 8'h10 ;
			data[61492] <= 8'h10 ;
			data[61493] <= 8'h10 ;
			data[61494] <= 8'h10 ;
			data[61495] <= 8'h10 ;
			data[61496] <= 8'h10 ;
			data[61497] <= 8'h10 ;
			data[61498] <= 8'h10 ;
			data[61499] <= 8'h10 ;
			data[61500] <= 8'h10 ;
			data[61501] <= 8'h10 ;
			data[61502] <= 8'h10 ;
			data[61503] <= 8'h10 ;
			data[61504] <= 8'h10 ;
			data[61505] <= 8'h10 ;
			data[61506] <= 8'h10 ;
			data[61507] <= 8'h10 ;
			data[61508] <= 8'h10 ;
			data[61509] <= 8'h10 ;
			data[61510] <= 8'h10 ;
			data[61511] <= 8'h10 ;
			data[61512] <= 8'h10 ;
			data[61513] <= 8'h10 ;
			data[61514] <= 8'h10 ;
			data[61515] <= 8'h10 ;
			data[61516] <= 8'h10 ;
			data[61517] <= 8'h10 ;
			data[61518] <= 8'h10 ;
			data[61519] <= 8'h10 ;
			data[61520] <= 8'h10 ;
			data[61521] <= 8'h10 ;
			data[61522] <= 8'h10 ;
			data[61523] <= 8'h10 ;
			data[61524] <= 8'h10 ;
			data[61525] <= 8'h10 ;
			data[61526] <= 8'h10 ;
			data[61527] <= 8'h10 ;
			data[61528] <= 8'h10 ;
			data[61529] <= 8'h10 ;
			data[61530] <= 8'h10 ;
			data[61531] <= 8'h10 ;
			data[61532] <= 8'h10 ;
			data[61533] <= 8'h10 ;
			data[61534] <= 8'h10 ;
			data[61535] <= 8'h10 ;
			data[61536] <= 8'h10 ;
			data[61537] <= 8'h10 ;
			data[61538] <= 8'h10 ;
			data[61539] <= 8'h10 ;
			data[61540] <= 8'h10 ;
			data[61541] <= 8'h10 ;
			data[61542] <= 8'h10 ;
			data[61543] <= 8'h10 ;
			data[61544] <= 8'h10 ;
			data[61545] <= 8'h10 ;
			data[61546] <= 8'h10 ;
			data[61547] <= 8'h10 ;
			data[61548] <= 8'h10 ;
			data[61549] <= 8'h10 ;
			data[61550] <= 8'h10 ;
			data[61551] <= 8'h10 ;
			data[61552] <= 8'h10 ;
			data[61553] <= 8'h10 ;
			data[61554] <= 8'h10 ;
			data[61555] <= 8'h10 ;
			data[61556] <= 8'h10 ;
			data[61557] <= 8'h10 ;
			data[61558] <= 8'h10 ;
			data[61559] <= 8'h10 ;
			data[61560] <= 8'h10 ;
			data[61561] <= 8'h10 ;
			data[61562] <= 8'h10 ;
			data[61563] <= 8'h10 ;
			data[61564] <= 8'h10 ;
			data[61565] <= 8'h10 ;
			data[61566] <= 8'h10 ;
			data[61567] <= 8'h10 ;
			data[61568] <= 8'h10 ;
			data[61569] <= 8'h10 ;
			data[61570] <= 8'h10 ;
			data[61571] <= 8'h10 ;
			data[61572] <= 8'h10 ;
			data[61573] <= 8'h10 ;
			data[61574] <= 8'h10 ;
			data[61575] <= 8'h10 ;
			data[61576] <= 8'h10 ;
			data[61577] <= 8'h10 ;
			data[61578] <= 8'h10 ;
			data[61579] <= 8'h10 ;
			data[61580] <= 8'h10 ;
			data[61581] <= 8'h10 ;
			data[61582] <= 8'h10 ;
			data[61583] <= 8'h10 ;
			data[61584] <= 8'h10 ;
			data[61585] <= 8'h10 ;
			data[61586] <= 8'h10 ;
			data[61587] <= 8'h10 ;
			data[61588] <= 8'h10 ;
			data[61589] <= 8'h10 ;
			data[61590] <= 8'h10 ;
			data[61591] <= 8'h10 ;
			data[61592] <= 8'h10 ;
			data[61593] <= 8'h10 ;
			data[61594] <= 8'h10 ;
			data[61595] <= 8'h10 ;
			data[61596] <= 8'h10 ;
			data[61597] <= 8'h10 ;
			data[61598] <= 8'h10 ;
			data[61599] <= 8'h10 ;
			data[61600] <= 8'h10 ;
			data[61601] <= 8'h10 ;
			data[61602] <= 8'h10 ;
			data[61603] <= 8'h10 ;
			data[61604] <= 8'h10 ;
			data[61605] <= 8'h10 ;
			data[61606] <= 8'h10 ;
			data[61607] <= 8'h10 ;
			data[61608] <= 8'h10 ;
			data[61609] <= 8'h10 ;
			data[61610] <= 8'h10 ;
			data[61611] <= 8'h10 ;
			data[61612] <= 8'h10 ;
			data[61613] <= 8'h10 ;
			data[61614] <= 8'h10 ;
			data[61615] <= 8'h10 ;
			data[61616] <= 8'h10 ;
			data[61617] <= 8'h10 ;
			data[61618] <= 8'h10 ;
			data[61619] <= 8'h10 ;
			data[61620] <= 8'h10 ;
			data[61621] <= 8'h10 ;
			data[61622] <= 8'h10 ;
			data[61623] <= 8'h10 ;
			data[61624] <= 8'h10 ;
			data[61625] <= 8'h10 ;
			data[61626] <= 8'h10 ;
			data[61627] <= 8'h10 ;
			data[61628] <= 8'h10 ;
			data[61629] <= 8'h10 ;
			data[61630] <= 8'h10 ;
			data[61631] <= 8'h10 ;
			data[61632] <= 8'h10 ;
			data[61633] <= 8'h10 ;
			data[61634] <= 8'h10 ;
			data[61635] <= 8'h10 ;
			data[61636] <= 8'h10 ;
			data[61637] <= 8'h10 ;
			data[61638] <= 8'h10 ;
			data[61639] <= 8'h10 ;
			data[61640] <= 8'h10 ;
			data[61641] <= 8'h10 ;
			data[61642] <= 8'h10 ;
			data[61643] <= 8'h10 ;
			data[61644] <= 8'h10 ;
			data[61645] <= 8'h10 ;
			data[61646] <= 8'h10 ;
			data[61647] <= 8'h10 ;
			data[61648] <= 8'h10 ;
			data[61649] <= 8'h10 ;
			data[61650] <= 8'h10 ;
			data[61651] <= 8'h10 ;
			data[61652] <= 8'h10 ;
			data[61653] <= 8'h10 ;
			data[61654] <= 8'h10 ;
			data[61655] <= 8'h10 ;
			data[61656] <= 8'h10 ;
			data[61657] <= 8'h10 ;
			data[61658] <= 8'h10 ;
			data[61659] <= 8'h10 ;
			data[61660] <= 8'h10 ;
			data[61661] <= 8'h10 ;
			data[61662] <= 8'h10 ;
			data[61663] <= 8'h10 ;
			data[61664] <= 8'h10 ;
			data[61665] <= 8'h10 ;
			data[61666] <= 8'h10 ;
			data[61667] <= 8'h10 ;
			data[61668] <= 8'h10 ;
			data[61669] <= 8'h10 ;
			data[61670] <= 8'h10 ;
			data[61671] <= 8'h10 ;
			data[61672] <= 8'h10 ;
			data[61673] <= 8'h10 ;
			data[61674] <= 8'h10 ;
			data[61675] <= 8'h10 ;
			data[61676] <= 8'h10 ;
			data[61677] <= 8'h10 ;
			data[61678] <= 8'h10 ;
			data[61679] <= 8'h10 ;
			data[61680] <= 8'h10 ;
			data[61681] <= 8'h10 ;
			data[61682] <= 8'h10 ;
			data[61683] <= 8'h10 ;
			data[61684] <= 8'h10 ;
			data[61685] <= 8'h10 ;
			data[61686] <= 8'h10 ;
			data[61687] <= 8'h10 ;
			data[61688] <= 8'h10 ;
			data[61689] <= 8'h10 ;
			data[61690] <= 8'h10 ;
			data[61691] <= 8'h10 ;
			data[61692] <= 8'h10 ;
			data[61693] <= 8'h10 ;
			data[61694] <= 8'h10 ;
			data[61695] <= 8'h10 ;
			data[61696] <= 8'h10 ;
			data[61697] <= 8'h10 ;
			data[61698] <= 8'h10 ;
			data[61699] <= 8'h10 ;
			data[61700] <= 8'h10 ;
			data[61701] <= 8'h10 ;
			data[61702] <= 8'h10 ;
			data[61703] <= 8'h10 ;
			data[61704] <= 8'h10 ;
			data[61705] <= 8'h10 ;
			data[61706] <= 8'h10 ;
			data[61707] <= 8'h10 ;
			data[61708] <= 8'h10 ;
			data[61709] <= 8'h10 ;
			data[61710] <= 8'h10 ;
			data[61711] <= 8'h10 ;
			data[61712] <= 8'h10 ;
			data[61713] <= 8'h10 ;
			data[61714] <= 8'h10 ;
			data[61715] <= 8'h10 ;
			data[61716] <= 8'h10 ;
			data[61717] <= 8'h10 ;
			data[61718] <= 8'h10 ;
			data[61719] <= 8'h10 ;
			data[61720] <= 8'h10 ;
			data[61721] <= 8'h10 ;
			data[61722] <= 8'h10 ;
			data[61723] <= 8'h10 ;
			data[61724] <= 8'h10 ;
			data[61725] <= 8'h10 ;
			data[61726] <= 8'h10 ;
			data[61727] <= 8'h10 ;
			data[61728] <= 8'h10 ;
			data[61729] <= 8'h10 ;
			data[61730] <= 8'h10 ;
			data[61731] <= 8'h10 ;
			data[61732] <= 8'h10 ;
			data[61733] <= 8'h10 ;
			data[61734] <= 8'h10 ;
			data[61735] <= 8'h10 ;
			data[61736] <= 8'h10 ;
			data[61737] <= 8'h10 ;
			data[61738] <= 8'h10 ;
			data[61739] <= 8'h10 ;
			data[61740] <= 8'h10 ;
			data[61741] <= 8'h10 ;
			data[61742] <= 8'h10 ;
			data[61743] <= 8'h10 ;
			data[61744] <= 8'h10 ;
			data[61745] <= 8'h10 ;
			data[61746] <= 8'h10 ;
			data[61747] <= 8'h10 ;
			data[61748] <= 8'h10 ;
			data[61749] <= 8'h10 ;
			data[61750] <= 8'h10 ;
			data[61751] <= 8'h10 ;
			data[61752] <= 8'h10 ;
			data[61753] <= 8'h10 ;
			data[61754] <= 8'h10 ;
			data[61755] <= 8'h10 ;
			data[61756] <= 8'h10 ;
			data[61757] <= 8'h10 ;
			data[61758] <= 8'h10 ;
			data[61759] <= 8'h10 ;
			data[61760] <= 8'h10 ;
			data[61761] <= 8'h10 ;
			data[61762] <= 8'h10 ;
			data[61763] <= 8'h10 ;
			data[61764] <= 8'h10 ;
			data[61765] <= 8'h10 ;
			data[61766] <= 8'h10 ;
			data[61767] <= 8'h10 ;
			data[61768] <= 8'h10 ;
			data[61769] <= 8'h10 ;
			data[61770] <= 8'h10 ;
			data[61771] <= 8'h10 ;
			data[61772] <= 8'h10 ;
			data[61773] <= 8'h10 ;
			data[61774] <= 8'h10 ;
			data[61775] <= 8'h10 ;
			data[61776] <= 8'h10 ;
			data[61777] <= 8'h10 ;
			data[61778] <= 8'h10 ;
			data[61779] <= 8'h10 ;
			data[61780] <= 8'h10 ;
			data[61781] <= 8'h10 ;
			data[61782] <= 8'h10 ;
			data[61783] <= 8'h10 ;
			data[61784] <= 8'h10 ;
			data[61785] <= 8'h10 ;
			data[61786] <= 8'h10 ;
			data[61787] <= 8'h10 ;
			data[61788] <= 8'h10 ;
			data[61789] <= 8'h10 ;
			data[61790] <= 8'h10 ;
			data[61791] <= 8'h10 ;
			data[61792] <= 8'h10 ;
			data[61793] <= 8'h10 ;
			data[61794] <= 8'h10 ;
			data[61795] <= 8'h10 ;
			data[61796] <= 8'h10 ;
			data[61797] <= 8'h10 ;
			data[61798] <= 8'h10 ;
			data[61799] <= 8'h10 ;
			data[61800] <= 8'h10 ;
			data[61801] <= 8'h10 ;
			data[61802] <= 8'h10 ;
			data[61803] <= 8'h10 ;
			data[61804] <= 8'h10 ;
			data[61805] <= 8'h10 ;
			data[61806] <= 8'h10 ;
			data[61807] <= 8'h10 ;
			data[61808] <= 8'h10 ;
			data[61809] <= 8'h10 ;
			data[61810] <= 8'h10 ;
			data[61811] <= 8'h10 ;
			data[61812] <= 8'h10 ;
			data[61813] <= 8'h10 ;
			data[61814] <= 8'h10 ;
			data[61815] <= 8'h10 ;
			data[61816] <= 8'h10 ;
			data[61817] <= 8'h10 ;
			data[61818] <= 8'h10 ;
			data[61819] <= 8'h10 ;
			data[61820] <= 8'h10 ;
			data[61821] <= 8'h10 ;
			data[61822] <= 8'h10 ;
			data[61823] <= 8'h10 ;
			data[61824] <= 8'h10 ;
			data[61825] <= 8'h10 ;
			data[61826] <= 8'h10 ;
			data[61827] <= 8'h10 ;
			data[61828] <= 8'h10 ;
			data[61829] <= 8'h10 ;
			data[61830] <= 8'h10 ;
			data[61831] <= 8'h10 ;
			data[61832] <= 8'h10 ;
			data[61833] <= 8'h10 ;
			data[61834] <= 8'h10 ;
			data[61835] <= 8'h10 ;
			data[61836] <= 8'h10 ;
			data[61837] <= 8'h10 ;
			data[61838] <= 8'h10 ;
			data[61839] <= 8'h10 ;
			data[61840] <= 8'h10 ;
			data[61841] <= 8'h10 ;
			data[61842] <= 8'h10 ;
			data[61843] <= 8'h10 ;
			data[61844] <= 8'h10 ;
			data[61845] <= 8'h10 ;
			data[61846] <= 8'h10 ;
			data[61847] <= 8'h10 ;
			data[61848] <= 8'h10 ;
			data[61849] <= 8'h10 ;
			data[61850] <= 8'h10 ;
			data[61851] <= 8'h10 ;
			data[61852] <= 8'h10 ;
			data[61853] <= 8'h10 ;
			data[61854] <= 8'h10 ;
			data[61855] <= 8'h10 ;
			data[61856] <= 8'h10 ;
			data[61857] <= 8'h10 ;
			data[61858] <= 8'h10 ;
			data[61859] <= 8'h10 ;
			data[61860] <= 8'h10 ;
			data[61861] <= 8'h10 ;
			data[61862] <= 8'h10 ;
			data[61863] <= 8'h10 ;
			data[61864] <= 8'h10 ;
			data[61865] <= 8'h10 ;
			data[61866] <= 8'h10 ;
			data[61867] <= 8'h10 ;
			data[61868] <= 8'h10 ;
			data[61869] <= 8'h10 ;
			data[61870] <= 8'h10 ;
			data[61871] <= 8'h10 ;
			data[61872] <= 8'h10 ;
			data[61873] <= 8'h10 ;
			data[61874] <= 8'h10 ;
			data[61875] <= 8'h10 ;
			data[61876] <= 8'h10 ;
			data[61877] <= 8'h10 ;
			data[61878] <= 8'h10 ;
			data[61879] <= 8'h10 ;
			data[61880] <= 8'h10 ;
			data[61881] <= 8'h10 ;
			data[61882] <= 8'h10 ;
			data[61883] <= 8'h10 ;
			data[61884] <= 8'h10 ;
			data[61885] <= 8'h10 ;
			data[61886] <= 8'h10 ;
			data[61887] <= 8'h10 ;
			data[61888] <= 8'h10 ;
			data[61889] <= 8'h10 ;
			data[61890] <= 8'h10 ;
			data[61891] <= 8'h10 ;
			data[61892] <= 8'h10 ;
			data[61893] <= 8'h10 ;
			data[61894] <= 8'h10 ;
			data[61895] <= 8'h10 ;
			data[61896] <= 8'h10 ;
			data[61897] <= 8'h10 ;
			data[61898] <= 8'h10 ;
			data[61899] <= 8'h10 ;
			data[61900] <= 8'h10 ;
			data[61901] <= 8'h10 ;
			data[61902] <= 8'h10 ;
			data[61903] <= 8'h10 ;
			data[61904] <= 8'h10 ;
			data[61905] <= 8'h10 ;
			data[61906] <= 8'h10 ;
			data[61907] <= 8'h10 ;
			data[61908] <= 8'h10 ;
			data[61909] <= 8'h10 ;
			data[61910] <= 8'h10 ;
			data[61911] <= 8'h10 ;
			data[61912] <= 8'h10 ;
			data[61913] <= 8'h10 ;
			data[61914] <= 8'h10 ;
			data[61915] <= 8'h10 ;
			data[61916] <= 8'h10 ;
			data[61917] <= 8'h10 ;
			data[61918] <= 8'h10 ;
			data[61919] <= 8'h10 ;
			data[61920] <= 8'h10 ;
			data[61921] <= 8'h10 ;
			data[61922] <= 8'h10 ;
			data[61923] <= 8'h10 ;
			data[61924] <= 8'h10 ;
			data[61925] <= 8'h10 ;
			data[61926] <= 8'h10 ;
			data[61927] <= 8'h10 ;
			data[61928] <= 8'h10 ;
			data[61929] <= 8'h10 ;
			data[61930] <= 8'h10 ;
			data[61931] <= 8'h10 ;
			data[61932] <= 8'h10 ;
			data[61933] <= 8'h10 ;
			data[61934] <= 8'h10 ;
			data[61935] <= 8'h10 ;
			data[61936] <= 8'h10 ;
			data[61937] <= 8'h10 ;
			data[61938] <= 8'h10 ;
			data[61939] <= 8'h10 ;
			data[61940] <= 8'h10 ;
			data[61941] <= 8'h10 ;
			data[61942] <= 8'h10 ;
			data[61943] <= 8'h10 ;
			data[61944] <= 8'h10 ;
			data[61945] <= 8'h10 ;
			data[61946] <= 8'h10 ;
			data[61947] <= 8'h10 ;
			data[61948] <= 8'h10 ;
			data[61949] <= 8'h10 ;
			data[61950] <= 8'h10 ;
			data[61951] <= 8'h10 ;
			data[61952] <= 8'h10 ;
			data[61953] <= 8'h10 ;
			data[61954] <= 8'h10 ;
			data[61955] <= 8'h10 ;
			data[61956] <= 8'h10 ;
			data[61957] <= 8'h10 ;
			data[61958] <= 8'h10 ;
			data[61959] <= 8'h10 ;
			data[61960] <= 8'h10 ;
			data[61961] <= 8'h10 ;
			data[61962] <= 8'h10 ;
			data[61963] <= 8'h10 ;
			data[61964] <= 8'h10 ;
			data[61965] <= 8'h10 ;
			data[61966] <= 8'h10 ;
			data[61967] <= 8'h10 ;
			data[61968] <= 8'h10 ;
			data[61969] <= 8'h10 ;
			data[61970] <= 8'h10 ;
			data[61971] <= 8'h10 ;
			data[61972] <= 8'h10 ;
			data[61973] <= 8'h10 ;
			data[61974] <= 8'h10 ;
			data[61975] <= 8'h10 ;
			data[61976] <= 8'h10 ;
			data[61977] <= 8'h10 ;
			data[61978] <= 8'h10 ;
			data[61979] <= 8'h10 ;
			data[61980] <= 8'h10 ;
			data[61981] <= 8'h10 ;
			data[61982] <= 8'h10 ;
			data[61983] <= 8'h10 ;
			data[61984] <= 8'h10 ;
			data[61985] <= 8'h10 ;
			data[61986] <= 8'h10 ;
			data[61987] <= 8'h10 ;
			data[61988] <= 8'h10 ;
			data[61989] <= 8'h10 ;
			data[61990] <= 8'h10 ;
			data[61991] <= 8'h10 ;
			data[61992] <= 8'h10 ;
			data[61993] <= 8'h10 ;
			data[61994] <= 8'h10 ;
			data[61995] <= 8'h10 ;
			data[61996] <= 8'h10 ;
			data[61997] <= 8'h10 ;
			data[61998] <= 8'h10 ;
			data[61999] <= 8'h10 ;
			data[62000] <= 8'h10 ;
			data[62001] <= 8'h10 ;
			data[62002] <= 8'h10 ;
			data[62003] <= 8'h10 ;
			data[62004] <= 8'h10 ;
			data[62005] <= 8'h10 ;
			data[62006] <= 8'h10 ;
			data[62007] <= 8'h10 ;
			data[62008] <= 8'h10 ;
			data[62009] <= 8'h10 ;
			data[62010] <= 8'h10 ;
			data[62011] <= 8'h10 ;
			data[62012] <= 8'h10 ;
			data[62013] <= 8'h10 ;
			data[62014] <= 8'h10 ;
			data[62015] <= 8'h10 ;
			data[62016] <= 8'h10 ;
			data[62017] <= 8'h10 ;
			data[62018] <= 8'h10 ;
			data[62019] <= 8'h10 ;
			data[62020] <= 8'h10 ;
			data[62021] <= 8'h10 ;
			data[62022] <= 8'h10 ;
			data[62023] <= 8'h10 ;
			data[62024] <= 8'h10 ;
			data[62025] <= 8'h10 ;
			data[62026] <= 8'h10 ;
			data[62027] <= 8'h10 ;
			data[62028] <= 8'h10 ;
			data[62029] <= 8'h10 ;
			data[62030] <= 8'h10 ;
			data[62031] <= 8'h10 ;
			data[62032] <= 8'h10 ;
			data[62033] <= 8'h10 ;
			data[62034] <= 8'h10 ;
			data[62035] <= 8'h10 ;
			data[62036] <= 8'h10 ;
			data[62037] <= 8'h10 ;
			data[62038] <= 8'h10 ;
			data[62039] <= 8'h10 ;
			data[62040] <= 8'h10 ;
			data[62041] <= 8'h10 ;
			data[62042] <= 8'h10 ;
			data[62043] <= 8'h10 ;
			data[62044] <= 8'h10 ;
			data[62045] <= 8'h10 ;
			data[62046] <= 8'h10 ;
			data[62047] <= 8'h10 ;
			data[62048] <= 8'h10 ;
			data[62049] <= 8'h10 ;
			data[62050] <= 8'h10 ;
			data[62051] <= 8'h10 ;
			data[62052] <= 8'h10 ;
			data[62053] <= 8'h10 ;
			data[62054] <= 8'h10 ;
			data[62055] <= 8'h10 ;
			data[62056] <= 8'h10 ;
			data[62057] <= 8'h10 ;
			data[62058] <= 8'h10 ;
			data[62059] <= 8'h10 ;
			data[62060] <= 8'h10 ;
			data[62061] <= 8'h10 ;
			data[62062] <= 8'h10 ;
			data[62063] <= 8'h10 ;
			data[62064] <= 8'h10 ;
			data[62065] <= 8'h10 ;
			data[62066] <= 8'h10 ;
			data[62067] <= 8'h10 ;
			data[62068] <= 8'h10 ;
			data[62069] <= 8'h10 ;
			data[62070] <= 8'h10 ;
			data[62071] <= 8'h10 ;
			data[62072] <= 8'h10 ;
			data[62073] <= 8'h10 ;
			data[62074] <= 8'h10 ;
			data[62075] <= 8'h10 ;
			data[62076] <= 8'h10 ;
			data[62077] <= 8'h10 ;
			data[62078] <= 8'h10 ;
			data[62079] <= 8'h10 ;
			data[62080] <= 8'h10 ;
			data[62081] <= 8'h10 ;
			data[62082] <= 8'h10 ;
			data[62083] <= 8'h10 ;
			data[62084] <= 8'h10 ;
			data[62085] <= 8'h10 ;
			data[62086] <= 8'h10 ;
			data[62087] <= 8'h10 ;
			data[62088] <= 8'h10 ;
			data[62089] <= 8'h10 ;
			data[62090] <= 8'h10 ;
			data[62091] <= 8'h10 ;
			data[62092] <= 8'h10 ;
			data[62093] <= 8'h10 ;
			data[62094] <= 8'h10 ;
			data[62095] <= 8'h10 ;
			data[62096] <= 8'h10 ;
			data[62097] <= 8'h10 ;
			data[62098] <= 8'h10 ;
			data[62099] <= 8'h10 ;
			data[62100] <= 8'h10 ;
			data[62101] <= 8'h10 ;
			data[62102] <= 8'h10 ;
			data[62103] <= 8'h10 ;
			data[62104] <= 8'h10 ;
			data[62105] <= 8'h10 ;
			data[62106] <= 8'h10 ;
			data[62107] <= 8'h10 ;
			data[62108] <= 8'h10 ;
			data[62109] <= 8'h10 ;
			data[62110] <= 8'h10 ;
			data[62111] <= 8'h10 ;
			data[62112] <= 8'h10 ;
			data[62113] <= 8'h10 ;
			data[62114] <= 8'h10 ;
			data[62115] <= 8'h10 ;
			data[62116] <= 8'h10 ;
			data[62117] <= 8'h10 ;
			data[62118] <= 8'h10 ;
			data[62119] <= 8'h10 ;
			data[62120] <= 8'h10 ;
			data[62121] <= 8'h10 ;
			data[62122] <= 8'h10 ;
			data[62123] <= 8'h10 ;
			data[62124] <= 8'h10 ;
			data[62125] <= 8'h10 ;
			data[62126] <= 8'h10 ;
			data[62127] <= 8'h10 ;
			data[62128] <= 8'h10 ;
			data[62129] <= 8'h10 ;
			data[62130] <= 8'h10 ;
			data[62131] <= 8'h10 ;
			data[62132] <= 8'h10 ;
			data[62133] <= 8'h10 ;
			data[62134] <= 8'h10 ;
			data[62135] <= 8'h10 ;
			data[62136] <= 8'h10 ;
			data[62137] <= 8'h10 ;
			data[62138] <= 8'h10 ;
			data[62139] <= 8'h10 ;
			data[62140] <= 8'h10 ;
			data[62141] <= 8'h10 ;
			data[62142] <= 8'h10 ;
			data[62143] <= 8'h10 ;
			data[62144] <= 8'h10 ;
			data[62145] <= 8'h10 ;
			data[62146] <= 8'h10 ;
			data[62147] <= 8'h10 ;
			data[62148] <= 8'h10 ;
			data[62149] <= 8'h10 ;
			data[62150] <= 8'h10 ;
			data[62151] <= 8'h10 ;
			data[62152] <= 8'h10 ;
			data[62153] <= 8'h10 ;
			data[62154] <= 8'h10 ;
			data[62155] <= 8'h10 ;
			data[62156] <= 8'h10 ;
			data[62157] <= 8'h10 ;
			data[62158] <= 8'h10 ;
			data[62159] <= 8'h10 ;
			data[62160] <= 8'h10 ;
			data[62161] <= 8'h10 ;
			data[62162] <= 8'h10 ;
			data[62163] <= 8'h10 ;
			data[62164] <= 8'h10 ;
			data[62165] <= 8'h10 ;
			data[62166] <= 8'h10 ;
			data[62167] <= 8'h10 ;
			data[62168] <= 8'h10 ;
			data[62169] <= 8'h10 ;
			data[62170] <= 8'h10 ;
			data[62171] <= 8'h10 ;
			data[62172] <= 8'h10 ;
			data[62173] <= 8'h10 ;
			data[62174] <= 8'h10 ;
			data[62175] <= 8'h10 ;
			data[62176] <= 8'h10 ;
			data[62177] <= 8'h10 ;
			data[62178] <= 8'h10 ;
			data[62179] <= 8'h10 ;
			data[62180] <= 8'h10 ;
			data[62181] <= 8'h10 ;
			data[62182] <= 8'h10 ;
			data[62183] <= 8'h10 ;
			data[62184] <= 8'h10 ;
			data[62185] <= 8'h10 ;
			data[62186] <= 8'h10 ;
			data[62187] <= 8'h10 ;
			data[62188] <= 8'h10 ;
			data[62189] <= 8'h10 ;
			data[62190] <= 8'h10 ;
			data[62191] <= 8'h10 ;
			data[62192] <= 8'h10 ;
			data[62193] <= 8'h10 ;
			data[62194] <= 8'h10 ;
			data[62195] <= 8'h10 ;
			data[62196] <= 8'h10 ;
			data[62197] <= 8'h10 ;
			data[62198] <= 8'h10 ;
			data[62199] <= 8'h10 ;
			data[62200] <= 8'h10 ;
			data[62201] <= 8'h10 ;
			data[62202] <= 8'h10 ;
			data[62203] <= 8'h10 ;
			data[62204] <= 8'h10 ;
			data[62205] <= 8'h10 ;
			data[62206] <= 8'h10 ;
			data[62207] <= 8'h10 ;
			data[62208] <= 8'h10 ;
			data[62209] <= 8'h10 ;
			data[62210] <= 8'h10 ;
			data[62211] <= 8'h10 ;
			data[62212] <= 8'h10 ;
			data[62213] <= 8'h10 ;
			data[62214] <= 8'h10 ;
			data[62215] <= 8'h10 ;
			data[62216] <= 8'h10 ;
			data[62217] <= 8'h10 ;
			data[62218] <= 8'h10 ;
			data[62219] <= 8'h10 ;
			data[62220] <= 8'h10 ;
			data[62221] <= 8'h10 ;
			data[62222] <= 8'h10 ;
			data[62223] <= 8'h10 ;
			data[62224] <= 8'h10 ;
			data[62225] <= 8'h10 ;
			data[62226] <= 8'h10 ;
			data[62227] <= 8'h10 ;
			data[62228] <= 8'h10 ;
			data[62229] <= 8'h10 ;
			data[62230] <= 8'h10 ;
			data[62231] <= 8'h10 ;
			data[62232] <= 8'h10 ;
			data[62233] <= 8'h10 ;
			data[62234] <= 8'h10 ;
			data[62235] <= 8'h10 ;
			data[62236] <= 8'h10 ;
			data[62237] <= 8'h10 ;
			data[62238] <= 8'h10 ;
			data[62239] <= 8'h10 ;
			data[62240] <= 8'h10 ;
			data[62241] <= 8'h10 ;
			data[62242] <= 8'h10 ;
			data[62243] <= 8'h10 ;
			data[62244] <= 8'h10 ;
			data[62245] <= 8'h10 ;
			data[62246] <= 8'h10 ;
			data[62247] <= 8'h10 ;
			data[62248] <= 8'h10 ;
			data[62249] <= 8'h10 ;
			data[62250] <= 8'h10 ;
			data[62251] <= 8'h10 ;
			data[62252] <= 8'h10 ;
			data[62253] <= 8'h10 ;
			data[62254] <= 8'h10 ;
			data[62255] <= 8'h10 ;
			data[62256] <= 8'h10 ;
			data[62257] <= 8'h10 ;
			data[62258] <= 8'h10 ;
			data[62259] <= 8'h10 ;
			data[62260] <= 8'h10 ;
			data[62261] <= 8'h10 ;
			data[62262] <= 8'h10 ;
			data[62263] <= 8'h10 ;
			data[62264] <= 8'h10 ;
			data[62265] <= 8'h10 ;
			data[62266] <= 8'h10 ;
			data[62267] <= 8'h10 ;
			data[62268] <= 8'h10 ;
			data[62269] <= 8'h10 ;
			data[62270] <= 8'h10 ;
			data[62271] <= 8'h10 ;
			data[62272] <= 8'h10 ;
			data[62273] <= 8'h10 ;
			data[62274] <= 8'h10 ;
			data[62275] <= 8'h10 ;
			data[62276] <= 8'h10 ;
			data[62277] <= 8'h10 ;
			data[62278] <= 8'h10 ;
			data[62279] <= 8'h10 ;
			data[62280] <= 8'h10 ;
			data[62281] <= 8'h10 ;
			data[62282] <= 8'h10 ;
			data[62283] <= 8'h10 ;
			data[62284] <= 8'h10 ;
			data[62285] <= 8'h10 ;
			data[62286] <= 8'h10 ;
			data[62287] <= 8'h10 ;
			data[62288] <= 8'h10 ;
			data[62289] <= 8'h10 ;
			data[62290] <= 8'h10 ;
			data[62291] <= 8'h10 ;
			data[62292] <= 8'h10 ;
			data[62293] <= 8'h10 ;
			data[62294] <= 8'h10 ;
			data[62295] <= 8'h10 ;
			data[62296] <= 8'h10 ;
			data[62297] <= 8'h10 ;
			data[62298] <= 8'h10 ;
			data[62299] <= 8'h10 ;
			data[62300] <= 8'h10 ;
			data[62301] <= 8'h10 ;
			data[62302] <= 8'h10 ;
			data[62303] <= 8'h10 ;
			data[62304] <= 8'h10 ;
			data[62305] <= 8'h10 ;
			data[62306] <= 8'h10 ;
			data[62307] <= 8'h10 ;
			data[62308] <= 8'h10 ;
			data[62309] <= 8'h10 ;
			data[62310] <= 8'h10 ;
			data[62311] <= 8'h10 ;
			data[62312] <= 8'h10 ;
			data[62313] <= 8'h10 ;
			data[62314] <= 8'h10 ;
			data[62315] <= 8'h10 ;
			data[62316] <= 8'h10 ;
			data[62317] <= 8'h10 ;
			data[62318] <= 8'h10 ;
			data[62319] <= 8'h10 ;
			data[62320] <= 8'h10 ;
			data[62321] <= 8'h10 ;
			data[62322] <= 8'h10 ;
			data[62323] <= 8'h10 ;
			data[62324] <= 8'h10 ;
			data[62325] <= 8'h10 ;
			data[62326] <= 8'h10 ;
			data[62327] <= 8'h10 ;
			data[62328] <= 8'h10 ;
			data[62329] <= 8'h10 ;
			data[62330] <= 8'h10 ;
			data[62331] <= 8'h10 ;
			data[62332] <= 8'h10 ;
			data[62333] <= 8'h10 ;
			data[62334] <= 8'h10 ;
			data[62335] <= 8'h10 ;
			data[62336] <= 8'h10 ;
			data[62337] <= 8'h10 ;
			data[62338] <= 8'h10 ;
			data[62339] <= 8'h10 ;
			data[62340] <= 8'h10 ;
			data[62341] <= 8'h10 ;
			data[62342] <= 8'h10 ;
			data[62343] <= 8'h10 ;
			data[62344] <= 8'h10 ;
			data[62345] <= 8'h10 ;
			data[62346] <= 8'h10 ;
			data[62347] <= 8'h10 ;
			data[62348] <= 8'h10 ;
			data[62349] <= 8'h10 ;
			data[62350] <= 8'h10 ;
			data[62351] <= 8'h10 ;
			data[62352] <= 8'h10 ;
			data[62353] <= 8'h10 ;
			data[62354] <= 8'h10 ;
			data[62355] <= 8'h10 ;
			data[62356] <= 8'h10 ;
			data[62357] <= 8'h10 ;
			data[62358] <= 8'h10 ;
			data[62359] <= 8'h10 ;
			data[62360] <= 8'h10 ;
			data[62361] <= 8'h10 ;
			data[62362] <= 8'h10 ;
			data[62363] <= 8'h10 ;
			data[62364] <= 8'h10 ;
			data[62365] <= 8'h10 ;
			data[62366] <= 8'h10 ;
			data[62367] <= 8'h10 ;
			data[62368] <= 8'h10 ;
			data[62369] <= 8'h10 ;
			data[62370] <= 8'h10 ;
			data[62371] <= 8'h10 ;
			data[62372] <= 8'h10 ;
			data[62373] <= 8'h10 ;
			data[62374] <= 8'h10 ;
			data[62375] <= 8'h10 ;
			data[62376] <= 8'h10 ;
			data[62377] <= 8'h10 ;
			data[62378] <= 8'h10 ;
			data[62379] <= 8'h10 ;
			data[62380] <= 8'h10 ;
			data[62381] <= 8'h10 ;
			data[62382] <= 8'h10 ;
			data[62383] <= 8'h10 ;
			data[62384] <= 8'h10 ;
			data[62385] <= 8'h10 ;
			data[62386] <= 8'h10 ;
			data[62387] <= 8'h10 ;
			data[62388] <= 8'h10 ;
			data[62389] <= 8'h10 ;
			data[62390] <= 8'h10 ;
			data[62391] <= 8'h10 ;
			data[62392] <= 8'h10 ;
			data[62393] <= 8'h10 ;
			data[62394] <= 8'h10 ;
			data[62395] <= 8'h10 ;
			data[62396] <= 8'h10 ;
			data[62397] <= 8'h10 ;
			data[62398] <= 8'h10 ;
			data[62399] <= 8'h10 ;
			data[62400] <= 8'h10 ;
			data[62401] <= 8'h10 ;
			data[62402] <= 8'h10 ;
			data[62403] <= 8'h10 ;
			data[62404] <= 8'h10 ;
			data[62405] <= 8'h10 ;
			data[62406] <= 8'h10 ;
			data[62407] <= 8'h10 ;
			data[62408] <= 8'h10 ;
			data[62409] <= 8'h10 ;
			data[62410] <= 8'h10 ;
			data[62411] <= 8'h10 ;
			data[62412] <= 8'h10 ;
			data[62413] <= 8'h10 ;
			data[62414] <= 8'h10 ;
			data[62415] <= 8'h10 ;
			data[62416] <= 8'h10 ;
			data[62417] <= 8'h10 ;
			data[62418] <= 8'h10 ;
			data[62419] <= 8'h10 ;
			data[62420] <= 8'h10 ;
			data[62421] <= 8'h10 ;
			data[62422] <= 8'h10 ;
			data[62423] <= 8'h10 ;
			data[62424] <= 8'h10 ;
			data[62425] <= 8'h10 ;
			data[62426] <= 8'h10 ;
			data[62427] <= 8'h10 ;
			data[62428] <= 8'h10 ;
			data[62429] <= 8'h10 ;
			data[62430] <= 8'h10 ;
			data[62431] <= 8'h10 ;
			data[62432] <= 8'h10 ;
			data[62433] <= 8'h10 ;
			data[62434] <= 8'h10 ;
			data[62435] <= 8'h10 ;
			data[62436] <= 8'h10 ;
			data[62437] <= 8'h10 ;
			data[62438] <= 8'h10 ;
			data[62439] <= 8'h10 ;
			data[62440] <= 8'h10 ;
			data[62441] <= 8'h10 ;
			data[62442] <= 8'h10 ;
			data[62443] <= 8'h10 ;
			data[62444] <= 8'h10 ;
			data[62445] <= 8'h10 ;
			data[62446] <= 8'h10 ;
			data[62447] <= 8'h10 ;
			data[62448] <= 8'h10 ;
			data[62449] <= 8'h10 ;
			data[62450] <= 8'h10 ;
			data[62451] <= 8'h10 ;
			data[62452] <= 8'h10 ;
			data[62453] <= 8'h10 ;
			data[62454] <= 8'h10 ;
			data[62455] <= 8'h10 ;
			data[62456] <= 8'h10 ;
			data[62457] <= 8'h10 ;
			data[62458] <= 8'h10 ;
			data[62459] <= 8'h10 ;
			data[62460] <= 8'h10 ;
			data[62461] <= 8'h10 ;
			data[62462] <= 8'h10 ;
			data[62463] <= 8'h10 ;
			data[62464] <= 8'h10 ;
			data[62465] <= 8'h10 ;
			data[62466] <= 8'h10 ;
			data[62467] <= 8'h10 ;
			data[62468] <= 8'h10 ;
			data[62469] <= 8'h10 ;
			data[62470] <= 8'h10 ;
			data[62471] <= 8'h10 ;
			data[62472] <= 8'h10 ;
			data[62473] <= 8'h10 ;
			data[62474] <= 8'h10 ;
			data[62475] <= 8'h10 ;
			data[62476] <= 8'h10 ;
			data[62477] <= 8'h10 ;
			data[62478] <= 8'h10 ;
			data[62479] <= 8'h10 ;
			data[62480] <= 8'h10 ;
			data[62481] <= 8'h10 ;
			data[62482] <= 8'h10 ;
			data[62483] <= 8'h10 ;
			data[62484] <= 8'h10 ;
			data[62485] <= 8'h10 ;
			data[62486] <= 8'h10 ;
			data[62487] <= 8'h10 ;
			data[62488] <= 8'h10 ;
			data[62489] <= 8'h10 ;
			data[62490] <= 8'h10 ;
			data[62491] <= 8'h10 ;
			data[62492] <= 8'h10 ;
			data[62493] <= 8'h10 ;
			data[62494] <= 8'h10 ;
			data[62495] <= 8'h10 ;
			data[62496] <= 8'h10 ;
			data[62497] <= 8'h10 ;
			data[62498] <= 8'h10 ;
			data[62499] <= 8'h10 ;
			data[62500] <= 8'h10 ;
			data[62501] <= 8'h10 ;
			data[62502] <= 8'h10 ;
			data[62503] <= 8'h10 ;
			data[62504] <= 8'h10 ;
			data[62505] <= 8'h10 ;
			data[62506] <= 8'h10 ;
			data[62507] <= 8'h10 ;
			data[62508] <= 8'h10 ;
			data[62509] <= 8'h10 ;
			data[62510] <= 8'h10 ;
			data[62511] <= 8'h10 ;
			data[62512] <= 8'h10 ;
			data[62513] <= 8'h10 ;
			data[62514] <= 8'h10 ;
			data[62515] <= 8'h10 ;
			data[62516] <= 8'h10 ;
			data[62517] <= 8'h10 ;
			data[62518] <= 8'h10 ;
			data[62519] <= 8'h10 ;
			data[62520] <= 8'h10 ;
			data[62521] <= 8'h10 ;
			data[62522] <= 8'h10 ;
			data[62523] <= 8'h10 ;
			data[62524] <= 8'h10 ;
			data[62525] <= 8'h10 ;
			data[62526] <= 8'h10 ;
			data[62527] <= 8'h10 ;
			data[62528] <= 8'h10 ;
			data[62529] <= 8'h10 ;
			data[62530] <= 8'h10 ;
			data[62531] <= 8'h10 ;
			data[62532] <= 8'h10 ;
			data[62533] <= 8'h10 ;
			data[62534] <= 8'h10 ;
			data[62535] <= 8'h10 ;
			data[62536] <= 8'h10 ;
			data[62537] <= 8'h10 ;
			data[62538] <= 8'h10 ;
			data[62539] <= 8'h10 ;
			data[62540] <= 8'h10 ;
			data[62541] <= 8'h10 ;
			data[62542] <= 8'h10 ;
			data[62543] <= 8'h10 ;
			data[62544] <= 8'h10 ;
			data[62545] <= 8'h10 ;
			data[62546] <= 8'h10 ;
			data[62547] <= 8'h10 ;
			data[62548] <= 8'h10 ;
			data[62549] <= 8'h10 ;
			data[62550] <= 8'h10 ;
			data[62551] <= 8'h10 ;
			data[62552] <= 8'h10 ;
			data[62553] <= 8'h10 ;
			data[62554] <= 8'h10 ;
			data[62555] <= 8'h10 ;
			data[62556] <= 8'h10 ;
			data[62557] <= 8'h10 ;
			data[62558] <= 8'h10 ;
			data[62559] <= 8'h10 ;
			data[62560] <= 8'h10 ;
			data[62561] <= 8'h10 ;
			data[62562] <= 8'h10 ;
			data[62563] <= 8'h10 ;
			data[62564] <= 8'h10 ;
			data[62565] <= 8'h10 ;
			data[62566] <= 8'h10 ;
			data[62567] <= 8'h10 ;
			data[62568] <= 8'h10 ;
			data[62569] <= 8'h10 ;
			data[62570] <= 8'h10 ;
			data[62571] <= 8'h10 ;
			data[62572] <= 8'h10 ;
			data[62573] <= 8'h10 ;
			data[62574] <= 8'h10 ;
			data[62575] <= 8'h10 ;
			data[62576] <= 8'h10 ;
			data[62577] <= 8'h10 ;
			data[62578] <= 8'h10 ;
			data[62579] <= 8'h10 ;
			data[62580] <= 8'h10 ;
			data[62581] <= 8'h10 ;
			data[62582] <= 8'h10 ;
			data[62583] <= 8'h10 ;
			data[62584] <= 8'h10 ;
			data[62585] <= 8'h10 ;
			data[62586] <= 8'h10 ;
			data[62587] <= 8'h10 ;
			data[62588] <= 8'h10 ;
			data[62589] <= 8'h10 ;
			data[62590] <= 8'h10 ;
			data[62591] <= 8'h10 ;
			data[62592] <= 8'h10 ;
			data[62593] <= 8'h10 ;
			data[62594] <= 8'h10 ;
			data[62595] <= 8'h10 ;
			data[62596] <= 8'h10 ;
			data[62597] <= 8'h10 ;
			data[62598] <= 8'h10 ;
			data[62599] <= 8'h10 ;
			data[62600] <= 8'h10 ;
			data[62601] <= 8'h10 ;
			data[62602] <= 8'h10 ;
			data[62603] <= 8'h10 ;
			data[62604] <= 8'h10 ;
			data[62605] <= 8'h10 ;
			data[62606] <= 8'h10 ;
			data[62607] <= 8'h10 ;
			data[62608] <= 8'h10 ;
			data[62609] <= 8'h10 ;
			data[62610] <= 8'h10 ;
			data[62611] <= 8'h10 ;
			data[62612] <= 8'h10 ;
			data[62613] <= 8'h10 ;
			data[62614] <= 8'h10 ;
			data[62615] <= 8'h10 ;
			data[62616] <= 8'h10 ;
			data[62617] <= 8'h10 ;
			data[62618] <= 8'h10 ;
			data[62619] <= 8'h10 ;
			data[62620] <= 8'h10 ;
			data[62621] <= 8'h10 ;
			data[62622] <= 8'h10 ;
			data[62623] <= 8'h10 ;
			data[62624] <= 8'h10 ;
			data[62625] <= 8'h10 ;
			data[62626] <= 8'h10 ;
			data[62627] <= 8'h10 ;
			data[62628] <= 8'h10 ;
			data[62629] <= 8'h10 ;
			data[62630] <= 8'h10 ;
			data[62631] <= 8'h10 ;
			data[62632] <= 8'h10 ;
			data[62633] <= 8'h10 ;
			data[62634] <= 8'h10 ;
			data[62635] <= 8'h10 ;
			data[62636] <= 8'h10 ;
			data[62637] <= 8'h10 ;
			data[62638] <= 8'h10 ;
			data[62639] <= 8'h10 ;
			data[62640] <= 8'h10 ;
			data[62641] <= 8'h10 ;
			data[62642] <= 8'h10 ;
			data[62643] <= 8'h10 ;
			data[62644] <= 8'h10 ;
			data[62645] <= 8'h10 ;
			data[62646] <= 8'h10 ;
			data[62647] <= 8'h10 ;
			data[62648] <= 8'h10 ;
			data[62649] <= 8'h10 ;
			data[62650] <= 8'h10 ;
			data[62651] <= 8'h10 ;
			data[62652] <= 8'h10 ;
			data[62653] <= 8'h10 ;
			data[62654] <= 8'h10 ;
			data[62655] <= 8'h10 ;
			data[62656] <= 8'h10 ;
			data[62657] <= 8'h10 ;
			data[62658] <= 8'h10 ;
			data[62659] <= 8'h10 ;
			data[62660] <= 8'h10 ;
			data[62661] <= 8'h10 ;
			data[62662] <= 8'h10 ;
			data[62663] <= 8'h10 ;
			data[62664] <= 8'h10 ;
			data[62665] <= 8'h10 ;
			data[62666] <= 8'h10 ;
			data[62667] <= 8'h10 ;
			data[62668] <= 8'h10 ;
			data[62669] <= 8'h10 ;
			data[62670] <= 8'h10 ;
			data[62671] <= 8'h10 ;
			data[62672] <= 8'h10 ;
			data[62673] <= 8'h10 ;
			data[62674] <= 8'h10 ;
			data[62675] <= 8'h10 ;
			data[62676] <= 8'h10 ;
			data[62677] <= 8'h10 ;
			data[62678] <= 8'h10 ;
			data[62679] <= 8'h10 ;
			data[62680] <= 8'h10 ;
			data[62681] <= 8'h10 ;
			data[62682] <= 8'h10 ;
			data[62683] <= 8'h10 ;
			data[62684] <= 8'h10 ;
			data[62685] <= 8'h10 ;
			data[62686] <= 8'h10 ;
			data[62687] <= 8'h10 ;
			data[62688] <= 8'h10 ;
			data[62689] <= 8'h10 ;
			data[62690] <= 8'h10 ;
			data[62691] <= 8'h10 ;
			data[62692] <= 8'h10 ;
			data[62693] <= 8'h10 ;
			data[62694] <= 8'h10 ;
			data[62695] <= 8'h10 ;
			data[62696] <= 8'h10 ;
			data[62697] <= 8'h10 ;
			data[62698] <= 8'h10 ;
			data[62699] <= 8'h10 ;
			data[62700] <= 8'h10 ;
			data[62701] <= 8'h10 ;
			data[62702] <= 8'h10 ;
			data[62703] <= 8'h10 ;
			data[62704] <= 8'h10 ;
			data[62705] <= 8'h10 ;
			data[62706] <= 8'h10 ;
			data[62707] <= 8'h10 ;
			data[62708] <= 8'h10 ;
			data[62709] <= 8'h10 ;
			data[62710] <= 8'h10 ;
			data[62711] <= 8'h10 ;
			data[62712] <= 8'h10 ;
			data[62713] <= 8'h10 ;
			data[62714] <= 8'h10 ;
			data[62715] <= 8'h10 ;
			data[62716] <= 8'h10 ;
			data[62717] <= 8'h10 ;
			data[62718] <= 8'h10 ;
			data[62719] <= 8'h10 ;
			data[62720] <= 8'h10 ;
			data[62721] <= 8'h10 ;
			data[62722] <= 8'h10 ;
			data[62723] <= 8'h10 ;
			data[62724] <= 8'h10 ;
			data[62725] <= 8'h10 ;
			data[62726] <= 8'h10 ;
			data[62727] <= 8'h10 ;
			data[62728] <= 8'h10 ;
			data[62729] <= 8'h10 ;
			data[62730] <= 8'h10 ;
			data[62731] <= 8'h10 ;
			data[62732] <= 8'h10 ;
			data[62733] <= 8'h10 ;
			data[62734] <= 8'h10 ;
			data[62735] <= 8'h10 ;
			data[62736] <= 8'h10 ;
			data[62737] <= 8'h10 ;
			data[62738] <= 8'h10 ;
			data[62739] <= 8'h10 ;
			data[62740] <= 8'h10 ;
			data[62741] <= 8'h10 ;
			data[62742] <= 8'h10 ;
			data[62743] <= 8'h10 ;
			data[62744] <= 8'h10 ;
			data[62745] <= 8'h10 ;
			data[62746] <= 8'h10 ;
			data[62747] <= 8'h10 ;
			data[62748] <= 8'h10 ;
			data[62749] <= 8'h10 ;
			data[62750] <= 8'h10 ;
			data[62751] <= 8'h10 ;
			data[62752] <= 8'h10 ;
			data[62753] <= 8'h10 ;
			data[62754] <= 8'h10 ;
			data[62755] <= 8'h10 ;
			data[62756] <= 8'h10 ;
			data[62757] <= 8'h10 ;
			data[62758] <= 8'h10 ;
			data[62759] <= 8'h10 ;
			data[62760] <= 8'h10 ;
			data[62761] <= 8'h10 ;
			data[62762] <= 8'h10 ;
			data[62763] <= 8'h10 ;
			data[62764] <= 8'h10 ;
			data[62765] <= 8'h10 ;
			data[62766] <= 8'h10 ;
			data[62767] <= 8'h10 ;
			data[62768] <= 8'h10 ;
			data[62769] <= 8'h10 ;
			data[62770] <= 8'h10 ;
			data[62771] <= 8'h10 ;
			data[62772] <= 8'h10 ;
			data[62773] <= 8'h10 ;
			data[62774] <= 8'h10 ;
			data[62775] <= 8'h10 ;
			data[62776] <= 8'h10 ;
			data[62777] <= 8'h10 ;
			data[62778] <= 8'h10 ;
			data[62779] <= 8'h10 ;
			data[62780] <= 8'h10 ;
			data[62781] <= 8'h10 ;
			data[62782] <= 8'h10 ;
			data[62783] <= 8'h10 ;
			data[62784] <= 8'h10 ;
			data[62785] <= 8'h10 ;
			data[62786] <= 8'h10 ;
			data[62787] <= 8'h10 ;
			data[62788] <= 8'h10 ;
			data[62789] <= 8'h10 ;
			data[62790] <= 8'h10 ;
			data[62791] <= 8'h10 ;
			data[62792] <= 8'h10 ;
			data[62793] <= 8'h10 ;
			data[62794] <= 8'h10 ;
			data[62795] <= 8'h10 ;
			data[62796] <= 8'h10 ;
			data[62797] <= 8'h10 ;
			data[62798] <= 8'h10 ;
			data[62799] <= 8'h10 ;
			data[62800] <= 8'h10 ;
			data[62801] <= 8'h10 ;
			data[62802] <= 8'h10 ;
			data[62803] <= 8'h10 ;
			data[62804] <= 8'h10 ;
			data[62805] <= 8'h10 ;
			data[62806] <= 8'h10 ;
			data[62807] <= 8'h10 ;
			data[62808] <= 8'h10 ;
			data[62809] <= 8'h10 ;
			data[62810] <= 8'h10 ;
			data[62811] <= 8'h10 ;
			data[62812] <= 8'h10 ;
			data[62813] <= 8'h10 ;
			data[62814] <= 8'h10 ;
			data[62815] <= 8'h10 ;
			data[62816] <= 8'h10 ;
			data[62817] <= 8'h10 ;
			data[62818] <= 8'h10 ;
			data[62819] <= 8'h10 ;
			data[62820] <= 8'h10 ;
			data[62821] <= 8'h10 ;
			data[62822] <= 8'h10 ;
			data[62823] <= 8'h10 ;
			data[62824] <= 8'h10 ;
			data[62825] <= 8'h10 ;
			data[62826] <= 8'h10 ;
			data[62827] <= 8'h10 ;
			data[62828] <= 8'h10 ;
			data[62829] <= 8'h10 ;
			data[62830] <= 8'h10 ;
			data[62831] <= 8'h10 ;
			data[62832] <= 8'h10 ;
			data[62833] <= 8'h10 ;
			data[62834] <= 8'h10 ;
			data[62835] <= 8'h10 ;
			data[62836] <= 8'h10 ;
			data[62837] <= 8'h10 ;
			data[62838] <= 8'h10 ;
			data[62839] <= 8'h10 ;
			data[62840] <= 8'h10 ;
			data[62841] <= 8'h10 ;
			data[62842] <= 8'h10 ;
			data[62843] <= 8'h10 ;
			data[62844] <= 8'h10 ;
			data[62845] <= 8'h10 ;
			data[62846] <= 8'h10 ;
			data[62847] <= 8'h10 ;
			data[62848] <= 8'h10 ;
			data[62849] <= 8'h10 ;
			data[62850] <= 8'h10 ;
			data[62851] <= 8'h10 ;
			data[62852] <= 8'h10 ;
			data[62853] <= 8'h10 ;
			data[62854] <= 8'h10 ;
			data[62855] <= 8'h10 ;
			data[62856] <= 8'h10 ;
			data[62857] <= 8'h10 ;
			data[62858] <= 8'h10 ;
			data[62859] <= 8'h10 ;
			data[62860] <= 8'h10 ;
			data[62861] <= 8'h10 ;
			data[62862] <= 8'h10 ;
			data[62863] <= 8'h10 ;
			data[62864] <= 8'h10 ;
			data[62865] <= 8'h10 ;
			data[62866] <= 8'h10 ;
			data[62867] <= 8'h10 ;
			data[62868] <= 8'h10 ;
			data[62869] <= 8'h10 ;
			data[62870] <= 8'h10 ;
			data[62871] <= 8'h10 ;
			data[62872] <= 8'h10 ;
			data[62873] <= 8'h10 ;
			data[62874] <= 8'h10 ;
			data[62875] <= 8'h10 ;
			data[62876] <= 8'h10 ;
			data[62877] <= 8'h10 ;
			data[62878] <= 8'h10 ;
			data[62879] <= 8'h10 ;
			data[62880] <= 8'h10 ;
			data[62881] <= 8'h10 ;
			data[62882] <= 8'h10 ;
			data[62883] <= 8'h10 ;
			data[62884] <= 8'h10 ;
			data[62885] <= 8'h10 ;
			data[62886] <= 8'h10 ;
			data[62887] <= 8'h10 ;
			data[62888] <= 8'h10 ;
			data[62889] <= 8'h10 ;
			data[62890] <= 8'h10 ;
			data[62891] <= 8'h10 ;
			data[62892] <= 8'h10 ;
			data[62893] <= 8'h10 ;
			data[62894] <= 8'h10 ;
			data[62895] <= 8'h10 ;
			data[62896] <= 8'h10 ;
			data[62897] <= 8'h10 ;
			data[62898] <= 8'h10 ;
			data[62899] <= 8'h10 ;
			data[62900] <= 8'h10 ;
			data[62901] <= 8'h10 ;
			data[62902] <= 8'h10 ;
			data[62903] <= 8'h10 ;
			data[62904] <= 8'h10 ;
			data[62905] <= 8'h10 ;
			data[62906] <= 8'h10 ;
			data[62907] <= 8'h10 ;
			data[62908] <= 8'h10 ;
			data[62909] <= 8'h10 ;
			data[62910] <= 8'h10 ;
			data[62911] <= 8'h10 ;
			data[62912] <= 8'h10 ;
			data[62913] <= 8'h10 ;
			data[62914] <= 8'h10 ;
			data[62915] <= 8'h10 ;
			data[62916] <= 8'h10 ;
			data[62917] <= 8'h10 ;
			data[62918] <= 8'h10 ;
			data[62919] <= 8'h10 ;
			data[62920] <= 8'h10 ;
			data[62921] <= 8'h10 ;
			data[62922] <= 8'h10 ;
			data[62923] <= 8'h10 ;
			data[62924] <= 8'h10 ;
			data[62925] <= 8'h10 ;
			data[62926] <= 8'h10 ;
			data[62927] <= 8'h10 ;
			data[62928] <= 8'h10 ;
			data[62929] <= 8'h10 ;
			data[62930] <= 8'h10 ;
			data[62931] <= 8'h10 ;
			data[62932] <= 8'h10 ;
			data[62933] <= 8'h10 ;
			data[62934] <= 8'h10 ;
			data[62935] <= 8'h10 ;
			data[62936] <= 8'h10 ;
			data[62937] <= 8'h10 ;
			data[62938] <= 8'h10 ;
			data[62939] <= 8'h10 ;
			data[62940] <= 8'h10 ;
			data[62941] <= 8'h10 ;
			data[62942] <= 8'h10 ;
			data[62943] <= 8'h10 ;
			data[62944] <= 8'h10 ;
			data[62945] <= 8'h10 ;
			data[62946] <= 8'h10 ;
			data[62947] <= 8'h10 ;
			data[62948] <= 8'h10 ;
			data[62949] <= 8'h10 ;
			data[62950] <= 8'h10 ;
			data[62951] <= 8'h10 ;
			data[62952] <= 8'h10 ;
			data[62953] <= 8'h10 ;
			data[62954] <= 8'h10 ;
			data[62955] <= 8'h10 ;
			data[62956] <= 8'h10 ;
			data[62957] <= 8'h10 ;
			data[62958] <= 8'h10 ;
			data[62959] <= 8'h10 ;
			data[62960] <= 8'h10 ;
			data[62961] <= 8'h10 ;
			data[62962] <= 8'h10 ;
			data[62963] <= 8'h10 ;
			data[62964] <= 8'h10 ;
			data[62965] <= 8'h10 ;
			data[62966] <= 8'h10 ;
			data[62967] <= 8'h10 ;
			data[62968] <= 8'h10 ;
			data[62969] <= 8'h10 ;
			data[62970] <= 8'h10 ;
			data[62971] <= 8'h10 ;
			data[62972] <= 8'h10 ;
			data[62973] <= 8'h10 ;
			data[62974] <= 8'h10 ;
			data[62975] <= 8'h10 ;
			data[62976] <= 8'h10 ;
			data[62977] <= 8'h10 ;
			data[62978] <= 8'h10 ;
			data[62979] <= 8'h10 ;
			data[62980] <= 8'h10 ;
			data[62981] <= 8'h10 ;
			data[62982] <= 8'h10 ;
			data[62983] <= 8'h10 ;
			data[62984] <= 8'h10 ;
			data[62985] <= 8'h10 ;
			data[62986] <= 8'h10 ;
			data[62987] <= 8'h10 ;
			data[62988] <= 8'h10 ;
			data[62989] <= 8'h10 ;
			data[62990] <= 8'h10 ;
			data[62991] <= 8'h10 ;
			data[62992] <= 8'h10 ;
			data[62993] <= 8'h10 ;
			data[62994] <= 8'h10 ;
			data[62995] <= 8'h10 ;
			data[62996] <= 8'h10 ;
			data[62997] <= 8'h10 ;
			data[62998] <= 8'h10 ;
			data[62999] <= 8'h10 ;
			data[63000] <= 8'h10 ;
			data[63001] <= 8'h10 ;
			data[63002] <= 8'h10 ;
			data[63003] <= 8'h10 ;
			data[63004] <= 8'h10 ;
			data[63005] <= 8'h10 ;
			data[63006] <= 8'h10 ;
			data[63007] <= 8'h10 ;
			data[63008] <= 8'h10 ;
			data[63009] <= 8'h10 ;
			data[63010] <= 8'h10 ;
			data[63011] <= 8'h10 ;
			data[63012] <= 8'h10 ;
			data[63013] <= 8'h10 ;
			data[63014] <= 8'h10 ;
			data[63015] <= 8'h10 ;
			data[63016] <= 8'h10 ;
			data[63017] <= 8'h10 ;
			data[63018] <= 8'h10 ;
			data[63019] <= 8'h10 ;
			data[63020] <= 8'h10 ;
			data[63021] <= 8'h10 ;
			data[63022] <= 8'h10 ;
			data[63023] <= 8'h10 ;
			data[63024] <= 8'h10 ;
			data[63025] <= 8'h10 ;
			data[63026] <= 8'h10 ;
			data[63027] <= 8'h10 ;
			data[63028] <= 8'h10 ;
			data[63029] <= 8'h10 ;
			data[63030] <= 8'h10 ;
			data[63031] <= 8'h10 ;
			data[63032] <= 8'h10 ;
			data[63033] <= 8'h10 ;
			data[63034] <= 8'h10 ;
			data[63035] <= 8'h10 ;
			data[63036] <= 8'h10 ;
			data[63037] <= 8'h10 ;
			data[63038] <= 8'h10 ;
			data[63039] <= 8'h10 ;
			data[63040] <= 8'h10 ;
			data[63041] <= 8'h10 ;
			data[63042] <= 8'h10 ;
			data[63043] <= 8'h10 ;
			data[63044] <= 8'h10 ;
			data[63045] <= 8'h10 ;
			data[63046] <= 8'h10 ;
			data[63047] <= 8'h10 ;
			data[63048] <= 8'h10 ;
			data[63049] <= 8'h10 ;
			data[63050] <= 8'h10 ;
			data[63051] <= 8'h10 ;
			data[63052] <= 8'h10 ;
			data[63053] <= 8'h10 ;
			data[63054] <= 8'h10 ;
			data[63055] <= 8'h10 ;
			data[63056] <= 8'h10 ;
			data[63057] <= 8'h10 ;
			data[63058] <= 8'h10 ;
			data[63059] <= 8'h10 ;
			data[63060] <= 8'h10 ;
			data[63061] <= 8'h10 ;
			data[63062] <= 8'h10 ;
			data[63063] <= 8'h10 ;
			data[63064] <= 8'h10 ;
			data[63065] <= 8'h10 ;
			data[63066] <= 8'h10 ;
			data[63067] <= 8'h10 ;
			data[63068] <= 8'h10 ;
			data[63069] <= 8'h10 ;
			data[63070] <= 8'h10 ;
			data[63071] <= 8'h10 ;
			data[63072] <= 8'h10 ;
			data[63073] <= 8'h10 ;
			data[63074] <= 8'h10 ;
			data[63075] <= 8'h10 ;
			data[63076] <= 8'h10 ;
			data[63077] <= 8'h10 ;
			data[63078] <= 8'h10 ;
			data[63079] <= 8'h10 ;
			data[63080] <= 8'h10 ;
			data[63081] <= 8'h10 ;
			data[63082] <= 8'h10 ;
			data[63083] <= 8'h10 ;
			data[63084] <= 8'h10 ;
			data[63085] <= 8'h10 ;
			data[63086] <= 8'h10 ;
			data[63087] <= 8'h10 ;
			data[63088] <= 8'h10 ;
			data[63089] <= 8'h10 ;
			data[63090] <= 8'h10 ;
			data[63091] <= 8'h10 ;
			data[63092] <= 8'h10 ;
			data[63093] <= 8'h10 ;
			data[63094] <= 8'h10 ;
			data[63095] <= 8'h10 ;
			data[63096] <= 8'h10 ;
			data[63097] <= 8'h10 ;
			data[63098] <= 8'h10 ;
			data[63099] <= 8'h10 ;
			data[63100] <= 8'h10 ;
			data[63101] <= 8'h10 ;
			data[63102] <= 8'h10 ;
			data[63103] <= 8'h10 ;
			data[63104] <= 8'h10 ;
			data[63105] <= 8'h10 ;
			data[63106] <= 8'h10 ;
			data[63107] <= 8'h10 ;
			data[63108] <= 8'h10 ;
			data[63109] <= 8'h10 ;
			data[63110] <= 8'h10 ;
			data[63111] <= 8'h10 ;
			data[63112] <= 8'h10 ;
			data[63113] <= 8'h10 ;
			data[63114] <= 8'h10 ;
			data[63115] <= 8'h10 ;
			data[63116] <= 8'h10 ;
			data[63117] <= 8'h10 ;
			data[63118] <= 8'h10 ;
			data[63119] <= 8'h10 ;
			data[63120] <= 8'h10 ;
			data[63121] <= 8'h10 ;
			data[63122] <= 8'h10 ;
			data[63123] <= 8'h10 ;
			data[63124] <= 8'h10 ;
			data[63125] <= 8'h10 ;
			data[63126] <= 8'h10 ;
			data[63127] <= 8'h10 ;
			data[63128] <= 8'h10 ;
			data[63129] <= 8'h10 ;
			data[63130] <= 8'h10 ;
			data[63131] <= 8'h10 ;
			data[63132] <= 8'h10 ;
			data[63133] <= 8'h10 ;
			data[63134] <= 8'h10 ;
			data[63135] <= 8'h10 ;
			data[63136] <= 8'h10 ;
			data[63137] <= 8'h10 ;
			data[63138] <= 8'h10 ;
			data[63139] <= 8'h10 ;
			data[63140] <= 8'h10 ;
			data[63141] <= 8'h10 ;
			data[63142] <= 8'h10 ;
			data[63143] <= 8'h10 ;
			data[63144] <= 8'h10 ;
			data[63145] <= 8'h10 ;
			data[63146] <= 8'h10 ;
			data[63147] <= 8'h10 ;
			data[63148] <= 8'h10 ;
			data[63149] <= 8'h10 ;
			data[63150] <= 8'h10 ;
			data[63151] <= 8'h10 ;
			data[63152] <= 8'h10 ;
			data[63153] <= 8'h10 ;
			data[63154] <= 8'h10 ;
			data[63155] <= 8'h10 ;
			data[63156] <= 8'h10 ;
			data[63157] <= 8'h10 ;
			data[63158] <= 8'h10 ;
			data[63159] <= 8'h10 ;
			data[63160] <= 8'h10 ;
			data[63161] <= 8'h10 ;
			data[63162] <= 8'h10 ;
			data[63163] <= 8'h10 ;
			data[63164] <= 8'h10 ;
			data[63165] <= 8'h10 ;
			data[63166] <= 8'h10 ;
			data[63167] <= 8'h10 ;
			data[63168] <= 8'h10 ;
			data[63169] <= 8'h10 ;
			data[63170] <= 8'h10 ;
			data[63171] <= 8'h10 ;
			data[63172] <= 8'h10 ;
			data[63173] <= 8'h10 ;
			data[63174] <= 8'h10 ;
			data[63175] <= 8'h10 ;
			data[63176] <= 8'h10 ;
			data[63177] <= 8'h10 ;
			data[63178] <= 8'h10 ;
			data[63179] <= 8'h10 ;
			data[63180] <= 8'h10 ;
			data[63181] <= 8'h10 ;
			data[63182] <= 8'h10 ;
			data[63183] <= 8'h10 ;
			data[63184] <= 8'h10 ;
			data[63185] <= 8'h10 ;
			data[63186] <= 8'h10 ;
			data[63187] <= 8'h10 ;
			data[63188] <= 8'h10 ;
			data[63189] <= 8'h10 ;
			data[63190] <= 8'h10 ;
			data[63191] <= 8'h10 ;
			data[63192] <= 8'h10 ;
			data[63193] <= 8'h10 ;
			data[63194] <= 8'h10 ;
			data[63195] <= 8'h10 ;
			data[63196] <= 8'h10 ;
			data[63197] <= 8'h10 ;
			data[63198] <= 8'h10 ;
			data[63199] <= 8'h10 ;
			data[63200] <= 8'h10 ;
			data[63201] <= 8'h10 ;
			data[63202] <= 8'h10 ;
			data[63203] <= 8'h10 ;
			data[63204] <= 8'h10 ;
			data[63205] <= 8'h10 ;
			data[63206] <= 8'h10 ;
			data[63207] <= 8'h10 ;
			data[63208] <= 8'h10 ;
			data[63209] <= 8'h10 ;
			data[63210] <= 8'h10 ;
			data[63211] <= 8'h10 ;
			data[63212] <= 8'h10 ;
			data[63213] <= 8'h10 ;
			data[63214] <= 8'h10 ;
			data[63215] <= 8'h10 ;
			data[63216] <= 8'h10 ;
			data[63217] <= 8'h10 ;
			data[63218] <= 8'h10 ;
			data[63219] <= 8'h10 ;
			data[63220] <= 8'h10 ;
			data[63221] <= 8'h10 ;
			data[63222] <= 8'h10 ;
			data[63223] <= 8'h10 ;
			data[63224] <= 8'h10 ;
			data[63225] <= 8'h10 ;
			data[63226] <= 8'h10 ;
			data[63227] <= 8'h10 ;
			data[63228] <= 8'h10 ;
			data[63229] <= 8'h10 ;
			data[63230] <= 8'h10 ;
			data[63231] <= 8'h10 ;
			data[63232] <= 8'h10 ;
			data[63233] <= 8'h10 ;
			data[63234] <= 8'h10 ;
			data[63235] <= 8'h10 ;
			data[63236] <= 8'h10 ;
			data[63237] <= 8'h10 ;
			data[63238] <= 8'h10 ;
			data[63239] <= 8'h10 ;
			data[63240] <= 8'h10 ;
			data[63241] <= 8'h10 ;
			data[63242] <= 8'h10 ;
			data[63243] <= 8'h10 ;
			data[63244] <= 8'h10 ;
			data[63245] <= 8'h10 ;
			data[63246] <= 8'h10 ;
			data[63247] <= 8'h10 ;
			data[63248] <= 8'h10 ;
			data[63249] <= 8'h10 ;
			data[63250] <= 8'h10 ;
			data[63251] <= 8'h10 ;
			data[63252] <= 8'h10 ;
			data[63253] <= 8'h10 ;
			data[63254] <= 8'h10 ;
			data[63255] <= 8'h10 ;
			data[63256] <= 8'h10 ;
			data[63257] <= 8'h10 ;
			data[63258] <= 8'h10 ;
			data[63259] <= 8'h10 ;
			data[63260] <= 8'h10 ;
			data[63261] <= 8'h10 ;
			data[63262] <= 8'h10 ;
			data[63263] <= 8'h10 ;
			data[63264] <= 8'h10 ;
			data[63265] <= 8'h10 ;
			data[63266] <= 8'h10 ;
			data[63267] <= 8'h10 ;
			data[63268] <= 8'h10 ;
			data[63269] <= 8'h10 ;
			data[63270] <= 8'h10 ;
			data[63271] <= 8'h10 ;
			data[63272] <= 8'h10 ;
			data[63273] <= 8'h10 ;
			data[63274] <= 8'h10 ;
			data[63275] <= 8'h10 ;
			data[63276] <= 8'h10 ;
			data[63277] <= 8'h10 ;
			data[63278] <= 8'h10 ;
			data[63279] <= 8'h10 ;
			data[63280] <= 8'h10 ;
			data[63281] <= 8'h10 ;
			data[63282] <= 8'h10 ;
			data[63283] <= 8'h10 ;
			data[63284] <= 8'h10 ;
			data[63285] <= 8'h10 ;
			data[63286] <= 8'h10 ;
			data[63287] <= 8'h10 ;
			data[63288] <= 8'h10 ;
			data[63289] <= 8'h10 ;
			data[63290] <= 8'h10 ;
			data[63291] <= 8'h10 ;
			data[63292] <= 8'h10 ;
			data[63293] <= 8'h10 ;
			data[63294] <= 8'h10 ;
			data[63295] <= 8'h10 ;
			data[63296] <= 8'h10 ;
			data[63297] <= 8'h10 ;
			data[63298] <= 8'h10 ;
			data[63299] <= 8'h10 ;
			data[63300] <= 8'h10 ;
			data[63301] <= 8'h10 ;
			data[63302] <= 8'h10 ;
			data[63303] <= 8'h10 ;
			data[63304] <= 8'h10 ;
			data[63305] <= 8'h10 ;
			data[63306] <= 8'h10 ;
			data[63307] <= 8'h10 ;
			data[63308] <= 8'h10 ;
			data[63309] <= 8'h10 ;
			data[63310] <= 8'h10 ;
			data[63311] <= 8'h10 ;
			data[63312] <= 8'h10 ;
			data[63313] <= 8'h10 ;
			data[63314] <= 8'h10 ;
			data[63315] <= 8'h10 ;
			data[63316] <= 8'h10 ;
			data[63317] <= 8'h10 ;
			data[63318] <= 8'h10 ;
			data[63319] <= 8'h10 ;
			data[63320] <= 8'h10 ;
			data[63321] <= 8'h10 ;
			data[63322] <= 8'h10 ;
			data[63323] <= 8'h10 ;
			data[63324] <= 8'h10 ;
			data[63325] <= 8'h10 ;
			data[63326] <= 8'h10 ;
			data[63327] <= 8'h10 ;
			data[63328] <= 8'h10 ;
			data[63329] <= 8'h10 ;
			data[63330] <= 8'h10 ;
			data[63331] <= 8'h10 ;
			data[63332] <= 8'h10 ;
			data[63333] <= 8'h10 ;
			data[63334] <= 8'h10 ;
			data[63335] <= 8'h10 ;
			data[63336] <= 8'h10 ;
			data[63337] <= 8'h10 ;
			data[63338] <= 8'h10 ;
			data[63339] <= 8'h10 ;
			data[63340] <= 8'h10 ;
			data[63341] <= 8'h10 ;
			data[63342] <= 8'h10 ;
			data[63343] <= 8'h10 ;
			data[63344] <= 8'h10 ;
			data[63345] <= 8'h10 ;
			data[63346] <= 8'h10 ;
			data[63347] <= 8'h10 ;
			data[63348] <= 8'h10 ;
			data[63349] <= 8'h10 ;
			data[63350] <= 8'h10 ;
			data[63351] <= 8'h10 ;
			data[63352] <= 8'h10 ;
			data[63353] <= 8'h10 ;
			data[63354] <= 8'h10 ;
			data[63355] <= 8'h10 ;
			data[63356] <= 8'h10 ;
			data[63357] <= 8'h10 ;
			data[63358] <= 8'h10 ;
			data[63359] <= 8'h10 ;
			data[63360] <= 8'h10 ;
			data[63361] <= 8'h10 ;
			data[63362] <= 8'h10 ;
			data[63363] <= 8'h10 ;
			data[63364] <= 8'h10 ;
			data[63365] <= 8'h10 ;
			data[63366] <= 8'h10 ;
			data[63367] <= 8'h10 ;
			data[63368] <= 8'h10 ;
			data[63369] <= 8'h10 ;
			data[63370] <= 8'h10 ;
			data[63371] <= 8'h10 ;
			data[63372] <= 8'h10 ;
			data[63373] <= 8'h10 ;
			data[63374] <= 8'h10 ;
			data[63375] <= 8'h10 ;
			data[63376] <= 8'h10 ;
			data[63377] <= 8'h10 ;
			data[63378] <= 8'h10 ;
			data[63379] <= 8'h10 ;
			data[63380] <= 8'h10 ;
			data[63381] <= 8'h10 ;
			data[63382] <= 8'h10 ;
			data[63383] <= 8'h10 ;
			data[63384] <= 8'h10 ;
			data[63385] <= 8'h10 ;
			data[63386] <= 8'h10 ;
			data[63387] <= 8'h10 ;
			data[63388] <= 8'h10 ;
			data[63389] <= 8'h10 ;
			data[63390] <= 8'h10 ;
			data[63391] <= 8'h10 ;
			data[63392] <= 8'h10 ;
			data[63393] <= 8'h10 ;
			data[63394] <= 8'h10 ;
			data[63395] <= 8'h10 ;
			data[63396] <= 8'h10 ;
			data[63397] <= 8'h10 ;
			data[63398] <= 8'h10 ;
			data[63399] <= 8'h10 ;
			data[63400] <= 8'h10 ;
			data[63401] <= 8'h10 ;
			data[63402] <= 8'h10 ;
			data[63403] <= 8'h10 ;
			data[63404] <= 8'h10 ;
			data[63405] <= 8'h10 ;
			data[63406] <= 8'h10 ;
			data[63407] <= 8'h10 ;
			data[63408] <= 8'h10 ;
			data[63409] <= 8'h10 ;
			data[63410] <= 8'h10 ;
			data[63411] <= 8'h10 ;
			data[63412] <= 8'h10 ;
			data[63413] <= 8'h10 ;
			data[63414] <= 8'h10 ;
			data[63415] <= 8'h10 ;
			data[63416] <= 8'h10 ;
			data[63417] <= 8'h10 ;
			data[63418] <= 8'h10 ;
			data[63419] <= 8'h10 ;
			data[63420] <= 8'h10 ;
			data[63421] <= 8'h10 ;
			data[63422] <= 8'h10 ;
			data[63423] <= 8'h10 ;
			data[63424] <= 8'h10 ;
			data[63425] <= 8'h10 ;
			data[63426] <= 8'h10 ;
			data[63427] <= 8'h10 ;
			data[63428] <= 8'h10 ;
			data[63429] <= 8'h10 ;
			data[63430] <= 8'h10 ;
			data[63431] <= 8'h10 ;
			data[63432] <= 8'h10 ;
			data[63433] <= 8'h10 ;
			data[63434] <= 8'h10 ;
			data[63435] <= 8'h10 ;
			data[63436] <= 8'h10 ;
			data[63437] <= 8'h10 ;
			data[63438] <= 8'h10 ;
			data[63439] <= 8'h10 ;
			data[63440] <= 8'h10 ;
			data[63441] <= 8'h10 ;
			data[63442] <= 8'h10 ;
			data[63443] <= 8'h10 ;
			data[63444] <= 8'h10 ;
			data[63445] <= 8'h10 ;
			data[63446] <= 8'h10 ;
			data[63447] <= 8'h10 ;
			data[63448] <= 8'h10 ;
			data[63449] <= 8'h10 ;
			data[63450] <= 8'h10 ;
			data[63451] <= 8'h10 ;
			data[63452] <= 8'h10 ;
			data[63453] <= 8'h10 ;
			data[63454] <= 8'h10 ;
			data[63455] <= 8'h10 ;
			data[63456] <= 8'h10 ;
			data[63457] <= 8'h10 ;
			data[63458] <= 8'h10 ;
			data[63459] <= 8'h10 ;
			data[63460] <= 8'h10 ;
			data[63461] <= 8'h10 ;
			data[63462] <= 8'h10 ;
			data[63463] <= 8'h10 ;
			data[63464] <= 8'h10 ;
			data[63465] <= 8'h10 ;
			data[63466] <= 8'h10 ;
			data[63467] <= 8'h10 ;
			data[63468] <= 8'h10 ;
			data[63469] <= 8'h10 ;
			data[63470] <= 8'h10 ;
			data[63471] <= 8'h10 ;
			data[63472] <= 8'h10 ;
			data[63473] <= 8'h10 ;
			data[63474] <= 8'h10 ;
			data[63475] <= 8'h10 ;
			data[63476] <= 8'h10 ;
			data[63477] <= 8'h10 ;
			data[63478] <= 8'h10 ;
			data[63479] <= 8'h10 ;
			data[63480] <= 8'h10 ;
			data[63481] <= 8'h10 ;
			data[63482] <= 8'h10 ;
			data[63483] <= 8'h10 ;
			data[63484] <= 8'h10 ;
			data[63485] <= 8'h10 ;
			data[63486] <= 8'h10 ;
			data[63487] <= 8'h10 ;
			data[63488] <= 8'h10 ;
			data[63489] <= 8'h10 ;
			data[63490] <= 8'h10 ;
			data[63491] <= 8'h10 ;
			data[63492] <= 8'h10 ;
			data[63493] <= 8'h10 ;
			data[63494] <= 8'h10 ;
			data[63495] <= 8'h10 ;
			data[63496] <= 8'h10 ;
			data[63497] <= 8'h10 ;
			data[63498] <= 8'h10 ;
			data[63499] <= 8'h10 ;
			data[63500] <= 8'h10 ;
			data[63501] <= 8'h10 ;
			data[63502] <= 8'h10 ;
			data[63503] <= 8'h10 ;
			data[63504] <= 8'h10 ;
			data[63505] <= 8'h10 ;
			data[63506] <= 8'h10 ;
			data[63507] <= 8'h10 ;
			data[63508] <= 8'h10 ;
			data[63509] <= 8'h10 ;
			data[63510] <= 8'h10 ;
			data[63511] <= 8'h10 ;
			data[63512] <= 8'h10 ;
			data[63513] <= 8'h10 ;
			data[63514] <= 8'h10 ;
			data[63515] <= 8'h10 ;
			data[63516] <= 8'h10 ;
			data[63517] <= 8'h10 ;
			data[63518] <= 8'h10 ;
			data[63519] <= 8'h10 ;
			data[63520] <= 8'h10 ;
			data[63521] <= 8'h10 ;
			data[63522] <= 8'h10 ;
			data[63523] <= 8'h10 ;
			data[63524] <= 8'h10 ;
			data[63525] <= 8'h10 ;
			data[63526] <= 8'h10 ;
			data[63527] <= 8'h10 ;
			data[63528] <= 8'h10 ;
			data[63529] <= 8'h10 ;
			data[63530] <= 8'h10 ;
			data[63531] <= 8'h10 ;
			data[63532] <= 8'h10 ;
			data[63533] <= 8'h10 ;
			data[63534] <= 8'h10 ;
			data[63535] <= 8'h10 ;
			data[63536] <= 8'h10 ;
			data[63537] <= 8'h10 ;
			data[63538] <= 8'h10 ;
			data[63539] <= 8'h10 ;
			data[63540] <= 8'h10 ;
			data[63541] <= 8'h10 ;
			data[63542] <= 8'h10 ;
			data[63543] <= 8'h10 ;
			data[63544] <= 8'h10 ;
			data[63545] <= 8'h10 ;
			data[63546] <= 8'h10 ;
			data[63547] <= 8'h10 ;
			data[63548] <= 8'h10 ;
			data[63549] <= 8'h10 ;
			data[63550] <= 8'h10 ;
			data[63551] <= 8'h10 ;
			data[63552] <= 8'h10 ;
			data[63553] <= 8'h10 ;
			data[63554] <= 8'h10 ;
			data[63555] <= 8'h10 ;
			data[63556] <= 8'h10 ;
			data[63557] <= 8'h10 ;
			data[63558] <= 8'h10 ;
			data[63559] <= 8'h10 ;
			data[63560] <= 8'h10 ;
			data[63561] <= 8'h10 ;
			data[63562] <= 8'h10 ;
			data[63563] <= 8'h10 ;
			data[63564] <= 8'h10 ;
			data[63565] <= 8'h10 ;
			data[63566] <= 8'h10 ;
			data[63567] <= 8'h10 ;
			data[63568] <= 8'h10 ;
			data[63569] <= 8'h10 ;
			data[63570] <= 8'h10 ;
			data[63571] <= 8'h10 ;
			data[63572] <= 8'h10 ;
			data[63573] <= 8'h10 ;
			data[63574] <= 8'h10 ;
			data[63575] <= 8'h10 ;
			data[63576] <= 8'h10 ;
			data[63577] <= 8'h10 ;
			data[63578] <= 8'h10 ;
			data[63579] <= 8'h10 ;
			data[63580] <= 8'h10 ;
			data[63581] <= 8'h10 ;
			data[63582] <= 8'h10 ;
			data[63583] <= 8'h10 ;
			data[63584] <= 8'h10 ;
			data[63585] <= 8'h10 ;
			data[63586] <= 8'h10 ;
			data[63587] <= 8'h10 ;
			data[63588] <= 8'h10 ;
			data[63589] <= 8'h10 ;
			data[63590] <= 8'h10 ;
			data[63591] <= 8'h10 ;
			data[63592] <= 8'h10 ;
			data[63593] <= 8'h10 ;
			data[63594] <= 8'h10 ;
			data[63595] <= 8'h10 ;
			data[63596] <= 8'h10 ;
			data[63597] <= 8'h10 ;
			data[63598] <= 8'h10 ;
			data[63599] <= 8'h10 ;
			data[63600] <= 8'h10 ;
			data[63601] <= 8'h10 ;
			data[63602] <= 8'h10 ;
			data[63603] <= 8'h10 ;
			data[63604] <= 8'h10 ;
			data[63605] <= 8'h10 ;
			data[63606] <= 8'h10 ;
			data[63607] <= 8'h10 ;
			data[63608] <= 8'h10 ;
			data[63609] <= 8'h10 ;
			data[63610] <= 8'h10 ;
			data[63611] <= 8'h10 ;
			data[63612] <= 8'h10 ;
			data[63613] <= 8'h10 ;
			data[63614] <= 8'h10 ;
			data[63615] <= 8'h10 ;
			data[63616] <= 8'h10 ;
			data[63617] <= 8'h10 ;
			data[63618] <= 8'h10 ;
			data[63619] <= 8'h10 ;
			data[63620] <= 8'h10 ;
			data[63621] <= 8'h10 ;
			data[63622] <= 8'h10 ;
			data[63623] <= 8'h10 ;
			data[63624] <= 8'h10 ;
			data[63625] <= 8'h10 ;
			data[63626] <= 8'h10 ;
			data[63627] <= 8'h10 ;
			data[63628] <= 8'h10 ;
			data[63629] <= 8'h10 ;
			data[63630] <= 8'h10 ;
			data[63631] <= 8'h10 ;
			data[63632] <= 8'h10 ;
			data[63633] <= 8'h10 ;
			data[63634] <= 8'h10 ;
			data[63635] <= 8'h10 ;
			data[63636] <= 8'h10 ;
			data[63637] <= 8'h10 ;
			data[63638] <= 8'h10 ;
			data[63639] <= 8'h10 ;
			data[63640] <= 8'h10 ;
			data[63641] <= 8'h10 ;
			data[63642] <= 8'h10 ;
			data[63643] <= 8'h10 ;
			data[63644] <= 8'h10 ;
			data[63645] <= 8'h10 ;
			data[63646] <= 8'h10 ;
			data[63647] <= 8'h10 ;
			data[63648] <= 8'h10 ;
			data[63649] <= 8'h10 ;
			data[63650] <= 8'h10 ;
			data[63651] <= 8'h10 ;
			data[63652] <= 8'h10 ;
			data[63653] <= 8'h10 ;
			data[63654] <= 8'h10 ;
			data[63655] <= 8'h10 ;
			data[63656] <= 8'h10 ;
			data[63657] <= 8'h10 ;
			data[63658] <= 8'h10 ;
			data[63659] <= 8'h10 ;
			data[63660] <= 8'h10 ;
			data[63661] <= 8'h10 ;
			data[63662] <= 8'h10 ;
			data[63663] <= 8'h10 ;
			data[63664] <= 8'h10 ;
			data[63665] <= 8'h10 ;
			data[63666] <= 8'h10 ;
			data[63667] <= 8'h10 ;
			data[63668] <= 8'h10 ;
			data[63669] <= 8'h10 ;
			data[63670] <= 8'h10 ;
			data[63671] <= 8'h10 ;
			data[63672] <= 8'h10 ;
			data[63673] <= 8'h10 ;
			data[63674] <= 8'h10 ;
			data[63675] <= 8'h10 ;
			data[63676] <= 8'h10 ;
			data[63677] <= 8'h10 ;
			data[63678] <= 8'h10 ;
			data[63679] <= 8'h10 ;
			data[63680] <= 8'h10 ;
			data[63681] <= 8'h10 ;
			data[63682] <= 8'h10 ;
			data[63683] <= 8'h10 ;
			data[63684] <= 8'h10 ;
			data[63685] <= 8'h10 ;
			data[63686] <= 8'h10 ;
			data[63687] <= 8'h10 ;
			data[63688] <= 8'h10 ;
			data[63689] <= 8'h10 ;
			data[63690] <= 8'h10 ;
			data[63691] <= 8'h10 ;
			data[63692] <= 8'h10 ;
			data[63693] <= 8'h10 ;
			data[63694] <= 8'h10 ;
			data[63695] <= 8'h10 ;
			data[63696] <= 8'h10 ;
			data[63697] <= 8'h10 ;
			data[63698] <= 8'h10 ;
			data[63699] <= 8'h10 ;
			data[63700] <= 8'h10 ;
			data[63701] <= 8'h10 ;
			data[63702] <= 8'h10 ;
			data[63703] <= 8'h10 ;
			data[63704] <= 8'h10 ;
			data[63705] <= 8'h10 ;
			data[63706] <= 8'h10 ;
			data[63707] <= 8'h10 ;
			data[63708] <= 8'h10 ;
			data[63709] <= 8'h10 ;
			data[63710] <= 8'h10 ;
			data[63711] <= 8'h10 ;
			data[63712] <= 8'h10 ;
			data[63713] <= 8'h10 ;
			data[63714] <= 8'h10 ;
			data[63715] <= 8'h10 ;
			data[63716] <= 8'h10 ;
			data[63717] <= 8'h10 ;
			data[63718] <= 8'h10 ;
			data[63719] <= 8'h10 ;
			data[63720] <= 8'h10 ;
			data[63721] <= 8'h10 ;
			data[63722] <= 8'h10 ;
			data[63723] <= 8'h10 ;
			data[63724] <= 8'h10 ;
			data[63725] <= 8'h10 ;
			data[63726] <= 8'h10 ;
			data[63727] <= 8'h10 ;
			data[63728] <= 8'h10 ;
			data[63729] <= 8'h10 ;
			data[63730] <= 8'h10 ;
			data[63731] <= 8'h10 ;
			data[63732] <= 8'h10 ;
			data[63733] <= 8'h10 ;
			data[63734] <= 8'h10 ;
			data[63735] <= 8'h10 ;
			data[63736] <= 8'h10 ;
			data[63737] <= 8'h10 ;
			data[63738] <= 8'h10 ;
			data[63739] <= 8'h10 ;
			data[63740] <= 8'h10 ;
			data[63741] <= 8'h10 ;
			data[63742] <= 8'h10 ;
			data[63743] <= 8'h10 ;
			data[63744] <= 8'h10 ;
			data[63745] <= 8'h10 ;
			data[63746] <= 8'h10 ;
			data[63747] <= 8'h10 ;
			data[63748] <= 8'h10 ;
			data[63749] <= 8'h10 ;
			data[63750] <= 8'h10 ;
			data[63751] <= 8'h10 ;
			data[63752] <= 8'h10 ;
			data[63753] <= 8'h10 ;
			data[63754] <= 8'h10 ;
			data[63755] <= 8'h10 ;
			data[63756] <= 8'h10 ;
			data[63757] <= 8'h10 ;
			data[63758] <= 8'h10 ;
			data[63759] <= 8'h10 ;
			data[63760] <= 8'h10 ;
			data[63761] <= 8'h10 ;
			data[63762] <= 8'h10 ;
			data[63763] <= 8'h10 ;
			data[63764] <= 8'h10 ;
			data[63765] <= 8'h10 ;
			data[63766] <= 8'h10 ;
			data[63767] <= 8'h10 ;
			data[63768] <= 8'h10 ;
			data[63769] <= 8'h10 ;
			data[63770] <= 8'h10 ;
			data[63771] <= 8'h10 ;
			data[63772] <= 8'h10 ;
			data[63773] <= 8'h10 ;
			data[63774] <= 8'h10 ;
			data[63775] <= 8'h10 ;
			data[63776] <= 8'h10 ;
			data[63777] <= 8'h10 ;
			data[63778] <= 8'h10 ;
			data[63779] <= 8'h10 ;
			data[63780] <= 8'h10 ;
			data[63781] <= 8'h10 ;
			data[63782] <= 8'h10 ;
			data[63783] <= 8'h10 ;
			data[63784] <= 8'h10 ;
			data[63785] <= 8'h10 ;
			data[63786] <= 8'h10 ;
			data[63787] <= 8'h10 ;
			data[63788] <= 8'h10 ;
			data[63789] <= 8'h10 ;
			data[63790] <= 8'h10 ;
			data[63791] <= 8'h10 ;
			data[63792] <= 8'h10 ;
			data[63793] <= 8'h10 ;
			data[63794] <= 8'h10 ;
			data[63795] <= 8'h10 ;
			data[63796] <= 8'h10 ;
			data[63797] <= 8'h10 ;
			data[63798] <= 8'h10 ;
			data[63799] <= 8'h10 ;
			data[63800] <= 8'h10 ;
			data[63801] <= 8'h10 ;
			data[63802] <= 8'h10 ;
			data[63803] <= 8'h10 ;
			data[63804] <= 8'h10 ;
			data[63805] <= 8'h10 ;
			data[63806] <= 8'h10 ;
			data[63807] <= 8'h10 ;
			data[63808] <= 8'h10 ;
			data[63809] <= 8'h10 ;
			data[63810] <= 8'h10 ;
			data[63811] <= 8'h10 ;
			data[63812] <= 8'h10 ;
			data[63813] <= 8'h10 ;
			data[63814] <= 8'h10 ;
			data[63815] <= 8'h10 ;
			data[63816] <= 8'h10 ;
			data[63817] <= 8'h10 ;
			data[63818] <= 8'h10 ;
			data[63819] <= 8'h10 ;
			data[63820] <= 8'h10 ;
			data[63821] <= 8'h10 ;
			data[63822] <= 8'h10 ;
			data[63823] <= 8'h10 ;
			data[63824] <= 8'h10 ;
			data[63825] <= 8'h10 ;
			data[63826] <= 8'h10 ;
			data[63827] <= 8'h10 ;
			data[63828] <= 8'h10 ;
			data[63829] <= 8'h10 ;
			data[63830] <= 8'h10 ;
			data[63831] <= 8'h10 ;
			data[63832] <= 8'h10 ;
			data[63833] <= 8'h10 ;
			data[63834] <= 8'h10 ;
			data[63835] <= 8'h10 ;
			data[63836] <= 8'h10 ;
			data[63837] <= 8'h10 ;
			data[63838] <= 8'h10 ;
			data[63839] <= 8'h10 ;
			data[63840] <= 8'h10 ;
			data[63841] <= 8'h10 ;
			data[63842] <= 8'h10 ;
			data[63843] <= 8'h10 ;
			data[63844] <= 8'h10 ;
			data[63845] <= 8'h10 ;
			data[63846] <= 8'h10 ;
			data[63847] <= 8'h10 ;
			data[63848] <= 8'h10 ;
			data[63849] <= 8'h10 ;
			data[63850] <= 8'h10 ;
			data[63851] <= 8'h10 ;
			data[63852] <= 8'h10 ;
			data[63853] <= 8'h10 ;
			data[63854] <= 8'h10 ;
			data[63855] <= 8'h10 ;
			data[63856] <= 8'h10 ;
			data[63857] <= 8'h10 ;
			data[63858] <= 8'h10 ;
			data[63859] <= 8'h10 ;
			data[63860] <= 8'h10 ;
			data[63861] <= 8'h10 ;
			data[63862] <= 8'h10 ;
			data[63863] <= 8'h10 ;
			data[63864] <= 8'h10 ;
			data[63865] <= 8'h10 ;
			data[63866] <= 8'h10 ;
			data[63867] <= 8'h10 ;
			data[63868] <= 8'h10 ;
			data[63869] <= 8'h10 ;
			data[63870] <= 8'h10 ;
			data[63871] <= 8'h10 ;
			data[63872] <= 8'h10 ;
			data[63873] <= 8'h10 ;
			data[63874] <= 8'h10 ;
			data[63875] <= 8'h10 ;
			data[63876] <= 8'h10 ;
			data[63877] <= 8'h10 ;
			data[63878] <= 8'h10 ;
			data[63879] <= 8'h10 ;
			data[63880] <= 8'h10 ;
			data[63881] <= 8'h10 ;
			data[63882] <= 8'h10 ;
			data[63883] <= 8'h10 ;
			data[63884] <= 8'h10 ;
			data[63885] <= 8'h10 ;
			data[63886] <= 8'h10 ;
			data[63887] <= 8'h10 ;
			data[63888] <= 8'h10 ;
			data[63889] <= 8'h10 ;
			data[63890] <= 8'h10 ;
			data[63891] <= 8'h10 ;
			data[63892] <= 8'h10 ;
			data[63893] <= 8'h10 ;
			data[63894] <= 8'h10 ;
			data[63895] <= 8'h10 ;
			data[63896] <= 8'h10 ;
			data[63897] <= 8'h10 ;
			data[63898] <= 8'h10 ;
			data[63899] <= 8'h10 ;
			data[63900] <= 8'h10 ;
			data[63901] <= 8'h10 ;
			data[63902] <= 8'h10 ;
			data[63903] <= 8'h10 ;
			data[63904] <= 8'h10 ;
			data[63905] <= 8'h10 ;
			data[63906] <= 8'h10 ;
			data[63907] <= 8'h10 ;
			data[63908] <= 8'h10 ;
			data[63909] <= 8'h10 ;
			data[63910] <= 8'h10 ;
			data[63911] <= 8'h10 ;
			data[63912] <= 8'h10 ;
			data[63913] <= 8'h10 ;
			data[63914] <= 8'h10 ;
			data[63915] <= 8'h10 ;
			data[63916] <= 8'h10 ;
			data[63917] <= 8'h10 ;
			data[63918] <= 8'h10 ;
			data[63919] <= 8'h10 ;
			data[63920] <= 8'h10 ;
			data[63921] <= 8'h10 ;
			data[63922] <= 8'h10 ;
			data[63923] <= 8'h10 ;
			data[63924] <= 8'h10 ;
			data[63925] <= 8'h10 ;
			data[63926] <= 8'h10 ;
			data[63927] <= 8'h10 ;
			data[63928] <= 8'h10 ;
			data[63929] <= 8'h10 ;
			data[63930] <= 8'h10 ;
			data[63931] <= 8'h10 ;
			data[63932] <= 8'h10 ;
			data[63933] <= 8'h10 ;
			data[63934] <= 8'h10 ;
			data[63935] <= 8'h10 ;
			data[63936] <= 8'h10 ;
			data[63937] <= 8'h10 ;
			data[63938] <= 8'h10 ;
			data[63939] <= 8'h10 ;
			data[63940] <= 8'h10 ;
			data[63941] <= 8'h10 ;
			data[63942] <= 8'h10 ;
			data[63943] <= 8'h10 ;
			data[63944] <= 8'h10 ;
			data[63945] <= 8'h10 ;
			data[63946] <= 8'h10 ;
			data[63947] <= 8'h10 ;
			data[63948] <= 8'h10 ;
			data[63949] <= 8'h10 ;
			data[63950] <= 8'h10 ;
			data[63951] <= 8'h10 ;
			data[63952] <= 8'h10 ;
			data[63953] <= 8'h10 ;
			data[63954] <= 8'h10 ;
			data[63955] <= 8'h10 ;
			data[63956] <= 8'h10 ;
			data[63957] <= 8'h10 ;
			data[63958] <= 8'h10 ;
			data[63959] <= 8'h10 ;
			data[63960] <= 8'h10 ;
			data[63961] <= 8'h10 ;
			data[63962] <= 8'h10 ;
			data[63963] <= 8'h10 ;
			data[63964] <= 8'h10 ;
			data[63965] <= 8'h10 ;
			data[63966] <= 8'h10 ;
			data[63967] <= 8'h10 ;
			data[63968] <= 8'h10 ;
			data[63969] <= 8'h10 ;
			data[63970] <= 8'h10 ;
			data[63971] <= 8'h10 ;
			data[63972] <= 8'h10 ;
			data[63973] <= 8'h10 ;
			data[63974] <= 8'h10 ;
			data[63975] <= 8'h10 ;
			data[63976] <= 8'h10 ;
			data[63977] <= 8'h10 ;
			data[63978] <= 8'h10 ;
			data[63979] <= 8'h10 ;
			data[63980] <= 8'h10 ;
			data[63981] <= 8'h10 ;
			data[63982] <= 8'h10 ;
			data[63983] <= 8'h10 ;
			data[63984] <= 8'h10 ;
			data[63985] <= 8'h10 ;
			data[63986] <= 8'h10 ;
			data[63987] <= 8'h10 ;
			data[63988] <= 8'h10 ;
			data[63989] <= 8'h10 ;
			data[63990] <= 8'h10 ;
			data[63991] <= 8'h10 ;
			data[63992] <= 8'h10 ;
			data[63993] <= 8'h10 ;
			data[63994] <= 8'h10 ;
			data[63995] <= 8'h10 ;
			data[63996] <= 8'h10 ;
			data[63997] <= 8'h10 ;
			data[63998] <= 8'h10 ;
			data[63999] <= 8'h10 ;
			data[64000] <= 8'h10 ;
			data[64001] <= 8'h10 ;
			data[64002] <= 8'h10 ;
			data[64003] <= 8'h10 ;
			data[64004] <= 8'h10 ;
			data[64005] <= 8'h10 ;
			data[64006] <= 8'h10 ;
			data[64007] <= 8'h10 ;
			data[64008] <= 8'h10 ;
			data[64009] <= 8'h10 ;
			data[64010] <= 8'h10 ;
			data[64011] <= 8'h10 ;
			data[64012] <= 8'h10 ;
			data[64013] <= 8'h10 ;
			data[64014] <= 8'h10 ;
			data[64015] <= 8'h10 ;
			data[64016] <= 8'h10 ;
			data[64017] <= 8'h10 ;
			data[64018] <= 8'h10 ;
			data[64019] <= 8'h10 ;
			data[64020] <= 8'h10 ;
			data[64021] <= 8'h10 ;
			data[64022] <= 8'h10 ;
			data[64023] <= 8'h10 ;
			data[64024] <= 8'h10 ;
			data[64025] <= 8'h10 ;
			data[64026] <= 8'h10 ;
			data[64027] <= 8'h10 ;
			data[64028] <= 8'h10 ;
			data[64029] <= 8'h10 ;
			data[64030] <= 8'h10 ;
			data[64031] <= 8'h10 ;
			data[64032] <= 8'h10 ;
			data[64033] <= 8'h10 ;
			data[64034] <= 8'h10 ;
			data[64035] <= 8'h10 ;
			data[64036] <= 8'h10 ;
			data[64037] <= 8'h10 ;
			data[64038] <= 8'h10 ;
			data[64039] <= 8'h10 ;
			data[64040] <= 8'h10 ;
			data[64041] <= 8'h10 ;
			data[64042] <= 8'h10 ;
			data[64043] <= 8'h10 ;
			data[64044] <= 8'h10 ;
			data[64045] <= 8'h10 ;
			data[64046] <= 8'h10 ;
			data[64047] <= 8'h10 ;
			data[64048] <= 8'h10 ;
			data[64049] <= 8'h10 ;
			data[64050] <= 8'h10 ;
			data[64051] <= 8'h10 ;
			data[64052] <= 8'h10 ;
			data[64053] <= 8'h10 ;
			data[64054] <= 8'h10 ;
			data[64055] <= 8'h10 ;
			data[64056] <= 8'h10 ;
			data[64057] <= 8'h10 ;
			data[64058] <= 8'h10 ;
			data[64059] <= 8'h10 ;
			data[64060] <= 8'h10 ;
			data[64061] <= 8'h10 ;
			data[64062] <= 8'h10 ;
			data[64063] <= 8'h10 ;
			data[64064] <= 8'h10 ;
			data[64065] <= 8'h10 ;
			data[64066] <= 8'h10 ;
			data[64067] <= 8'h10 ;
			data[64068] <= 8'h10 ;
			data[64069] <= 8'h10 ;
			data[64070] <= 8'h10 ;
			data[64071] <= 8'h10 ;
			data[64072] <= 8'h10 ;
			data[64073] <= 8'h10 ;
			data[64074] <= 8'h10 ;
			data[64075] <= 8'h10 ;
			data[64076] <= 8'h10 ;
			data[64077] <= 8'h10 ;
			data[64078] <= 8'h10 ;
			data[64079] <= 8'h10 ;
			data[64080] <= 8'h10 ;
			data[64081] <= 8'h10 ;
			data[64082] <= 8'h10 ;
			data[64083] <= 8'h10 ;
			data[64084] <= 8'h10 ;
			data[64085] <= 8'h10 ;
			data[64086] <= 8'h10 ;
			data[64087] <= 8'h10 ;
			data[64088] <= 8'h10 ;
			data[64089] <= 8'h10 ;
			data[64090] <= 8'h10 ;
			data[64091] <= 8'h10 ;
			data[64092] <= 8'h10 ;
			data[64093] <= 8'h10 ;
			data[64094] <= 8'h10 ;
			data[64095] <= 8'h10 ;
			data[64096] <= 8'h10 ;
			data[64097] <= 8'h10 ;
			data[64098] <= 8'h10 ;
			data[64099] <= 8'h10 ;
			data[64100] <= 8'h10 ;
			data[64101] <= 8'h10 ;
			data[64102] <= 8'h10 ;
			data[64103] <= 8'h10 ;
			data[64104] <= 8'h10 ;
			data[64105] <= 8'h10 ;
			data[64106] <= 8'h10 ;
			data[64107] <= 8'h10 ;
			data[64108] <= 8'h10 ;
			data[64109] <= 8'h10 ;
			data[64110] <= 8'h10 ;
			data[64111] <= 8'h10 ;
			data[64112] <= 8'h10 ;
			data[64113] <= 8'h10 ;
			data[64114] <= 8'h10 ;
			data[64115] <= 8'h10 ;
			data[64116] <= 8'h10 ;
			data[64117] <= 8'h10 ;
			data[64118] <= 8'h10 ;
			data[64119] <= 8'h10 ;
			data[64120] <= 8'h10 ;
			data[64121] <= 8'h10 ;
			data[64122] <= 8'h10 ;
			data[64123] <= 8'h10 ;
			data[64124] <= 8'h10 ;
			data[64125] <= 8'h10 ;
			data[64126] <= 8'h10 ;
			data[64127] <= 8'h10 ;
			data[64128] <= 8'h10 ;
			data[64129] <= 8'h10 ;
			data[64130] <= 8'h10 ;
			data[64131] <= 8'h10 ;
			data[64132] <= 8'h10 ;
			data[64133] <= 8'h10 ;
			data[64134] <= 8'h10 ;
			data[64135] <= 8'h10 ;
			data[64136] <= 8'h10 ;
			data[64137] <= 8'h10 ;
			data[64138] <= 8'h10 ;
			data[64139] <= 8'h10 ;
			data[64140] <= 8'h10 ;
			data[64141] <= 8'h10 ;
			data[64142] <= 8'h10 ;
			data[64143] <= 8'h10 ;
			data[64144] <= 8'h10 ;
			data[64145] <= 8'h10 ;
			data[64146] <= 8'h10 ;
			data[64147] <= 8'h10 ;
			data[64148] <= 8'h10 ;
			data[64149] <= 8'h10 ;
			data[64150] <= 8'h10 ;
			data[64151] <= 8'h10 ;
			data[64152] <= 8'h10 ;
			data[64153] <= 8'h10 ;
			data[64154] <= 8'h10 ;
			data[64155] <= 8'h10 ;
			data[64156] <= 8'h10 ;
			data[64157] <= 8'h10 ;
			data[64158] <= 8'h10 ;
			data[64159] <= 8'h10 ;
			data[64160] <= 8'h10 ;
			data[64161] <= 8'h10 ;
			data[64162] <= 8'h10 ;
			data[64163] <= 8'h10 ;
			data[64164] <= 8'h10 ;
			data[64165] <= 8'h10 ;
			data[64166] <= 8'h10 ;
			data[64167] <= 8'h10 ;
			data[64168] <= 8'h10 ;
			data[64169] <= 8'h10 ;
			data[64170] <= 8'h10 ;
			data[64171] <= 8'h10 ;
			data[64172] <= 8'h10 ;
			data[64173] <= 8'h10 ;
			data[64174] <= 8'h10 ;
			data[64175] <= 8'h10 ;
			data[64176] <= 8'h10 ;
			data[64177] <= 8'h10 ;
			data[64178] <= 8'h10 ;
			data[64179] <= 8'h10 ;
			data[64180] <= 8'h10 ;
			data[64181] <= 8'h10 ;
			data[64182] <= 8'h10 ;
			data[64183] <= 8'h10 ;
			data[64184] <= 8'h10 ;
			data[64185] <= 8'h10 ;
			data[64186] <= 8'h10 ;
			data[64187] <= 8'h10 ;
			data[64188] <= 8'h10 ;
			data[64189] <= 8'h10 ;
			data[64190] <= 8'h10 ;
			data[64191] <= 8'h10 ;
			data[64192] <= 8'h10 ;
			data[64193] <= 8'h10 ;
			data[64194] <= 8'h10 ;
			data[64195] <= 8'h10 ;
			data[64196] <= 8'h10 ;
			data[64197] <= 8'h10 ;
			data[64198] <= 8'h10 ;
			data[64199] <= 8'h10 ;
			data[64200] <= 8'h10 ;
			data[64201] <= 8'h10 ;
			data[64202] <= 8'h10 ;
			data[64203] <= 8'h10 ;
			data[64204] <= 8'h10 ;
			data[64205] <= 8'h10 ;
			data[64206] <= 8'h10 ;
			data[64207] <= 8'h10 ;
			data[64208] <= 8'h10 ;
			data[64209] <= 8'h10 ;
			data[64210] <= 8'h10 ;
			data[64211] <= 8'h10 ;
			data[64212] <= 8'h10 ;
			data[64213] <= 8'h10 ;
			data[64214] <= 8'h10 ;
			data[64215] <= 8'h10 ;
			data[64216] <= 8'h10 ;
			data[64217] <= 8'h10 ;
			data[64218] <= 8'h10 ;
			data[64219] <= 8'h10 ;
			data[64220] <= 8'h10 ;
			data[64221] <= 8'h10 ;
			data[64222] <= 8'h10 ;
			data[64223] <= 8'h10 ;
			data[64224] <= 8'h10 ;
			data[64225] <= 8'h10 ;
			data[64226] <= 8'h10 ;
			data[64227] <= 8'h10 ;
			data[64228] <= 8'h10 ;
			data[64229] <= 8'h10 ;
			data[64230] <= 8'h10 ;
			data[64231] <= 8'h10 ;
			data[64232] <= 8'h10 ;
			data[64233] <= 8'h10 ;
			data[64234] <= 8'h10 ;
			data[64235] <= 8'h10 ;
			data[64236] <= 8'h10 ;
			data[64237] <= 8'h10 ;
			data[64238] <= 8'h10 ;
			data[64239] <= 8'h10 ;
			data[64240] <= 8'h10 ;
			data[64241] <= 8'h10 ;
			data[64242] <= 8'h10 ;
			data[64243] <= 8'h10 ;
			data[64244] <= 8'h10 ;
			data[64245] <= 8'h10 ;
			data[64246] <= 8'h10 ;
			data[64247] <= 8'h10 ;
			data[64248] <= 8'h10 ;
			data[64249] <= 8'h10 ;
			data[64250] <= 8'h10 ;
			data[64251] <= 8'h10 ;
			data[64252] <= 8'h10 ;
			data[64253] <= 8'h10 ;
			data[64254] <= 8'h10 ;
			data[64255] <= 8'h10 ;
			data[64256] <= 8'h10 ;
			data[64257] <= 8'h10 ;
			data[64258] <= 8'h10 ;
			data[64259] <= 8'h10 ;
			data[64260] <= 8'h10 ;
			data[64261] <= 8'h10 ;
			data[64262] <= 8'h10 ;
			data[64263] <= 8'h10 ;
			data[64264] <= 8'h10 ;
			data[64265] <= 8'h10 ;
			data[64266] <= 8'h10 ;
			data[64267] <= 8'h10 ;
			data[64268] <= 8'h10 ;
			data[64269] <= 8'h10 ;
			data[64270] <= 8'h10 ;
			data[64271] <= 8'h10 ;
			data[64272] <= 8'h10 ;
			data[64273] <= 8'h10 ;
			data[64274] <= 8'h10 ;
			data[64275] <= 8'h10 ;
			data[64276] <= 8'h10 ;
			data[64277] <= 8'h10 ;
			data[64278] <= 8'h10 ;
			data[64279] <= 8'h10 ;
			data[64280] <= 8'h10 ;
			data[64281] <= 8'h10 ;
			data[64282] <= 8'h10 ;
			data[64283] <= 8'h10 ;
			data[64284] <= 8'h10 ;
			data[64285] <= 8'h10 ;
			data[64286] <= 8'h10 ;
			data[64287] <= 8'h10 ;
			data[64288] <= 8'h10 ;
			data[64289] <= 8'h10 ;
			data[64290] <= 8'h10 ;
			data[64291] <= 8'h10 ;
			data[64292] <= 8'h10 ;
			data[64293] <= 8'h10 ;
			data[64294] <= 8'h10 ;
			data[64295] <= 8'h10 ;
			data[64296] <= 8'h10 ;
			data[64297] <= 8'h10 ;
			data[64298] <= 8'h10 ;
			data[64299] <= 8'h10 ;
			data[64300] <= 8'h10 ;
			data[64301] <= 8'h10 ;
			data[64302] <= 8'h10 ;
			data[64303] <= 8'h10 ;
			data[64304] <= 8'h10 ;
			data[64305] <= 8'h10 ;
			data[64306] <= 8'h10 ;
			data[64307] <= 8'h10 ;
			data[64308] <= 8'h10 ;
			data[64309] <= 8'h10 ;
			data[64310] <= 8'h10 ;
			data[64311] <= 8'h10 ;
			data[64312] <= 8'h10 ;
			data[64313] <= 8'h10 ;
			data[64314] <= 8'h10 ;
			data[64315] <= 8'h10 ;
			data[64316] <= 8'h10 ;
			data[64317] <= 8'h10 ;
			data[64318] <= 8'h10 ;
			data[64319] <= 8'h10 ;
			data[64320] <= 8'h10 ;
			data[64321] <= 8'h10 ;
			data[64322] <= 8'h10 ;
			data[64323] <= 8'h10 ;
			data[64324] <= 8'h10 ;
			data[64325] <= 8'h10 ;
			data[64326] <= 8'h10 ;
			data[64327] <= 8'h10 ;
			data[64328] <= 8'h10 ;
			data[64329] <= 8'h10 ;
			data[64330] <= 8'h10 ;
			data[64331] <= 8'h10 ;
			data[64332] <= 8'h10 ;
			data[64333] <= 8'h10 ;
			data[64334] <= 8'h10 ;
			data[64335] <= 8'h10 ;
			data[64336] <= 8'h10 ;
			data[64337] <= 8'h10 ;
			data[64338] <= 8'h10 ;
			data[64339] <= 8'h10 ;
			data[64340] <= 8'h10 ;
			data[64341] <= 8'h10 ;
			data[64342] <= 8'h10 ;
			data[64343] <= 8'h10 ;
			data[64344] <= 8'h10 ;
			data[64345] <= 8'h10 ;
			data[64346] <= 8'h10 ;
			data[64347] <= 8'h10 ;
			data[64348] <= 8'h10 ;
			data[64349] <= 8'h10 ;
			data[64350] <= 8'h10 ;
			data[64351] <= 8'h10 ;
			data[64352] <= 8'h10 ;
			data[64353] <= 8'h10 ;
			data[64354] <= 8'h10 ;
			data[64355] <= 8'h10 ;
			data[64356] <= 8'h10 ;
			data[64357] <= 8'h10 ;
			data[64358] <= 8'h10 ;
			data[64359] <= 8'h10 ;
			data[64360] <= 8'h10 ;
			data[64361] <= 8'h10 ;
			data[64362] <= 8'h10 ;
			data[64363] <= 8'h10 ;
			data[64364] <= 8'h10 ;
			data[64365] <= 8'h10 ;
			data[64366] <= 8'h10 ;
			data[64367] <= 8'h10 ;
			data[64368] <= 8'h10 ;
			data[64369] <= 8'h10 ;
			data[64370] <= 8'h10 ;
			data[64371] <= 8'h10 ;
			data[64372] <= 8'h10 ;
			data[64373] <= 8'h10 ;
			data[64374] <= 8'h10 ;
			data[64375] <= 8'h10 ;
			data[64376] <= 8'h10 ;
			data[64377] <= 8'h10 ;
			data[64378] <= 8'h10 ;
			data[64379] <= 8'h10 ;
			data[64380] <= 8'h10 ;
			data[64381] <= 8'h10 ;
			data[64382] <= 8'h10 ;
			data[64383] <= 8'h10 ;
			data[64384] <= 8'h10 ;
			data[64385] <= 8'h10 ;
			data[64386] <= 8'h10 ;
			data[64387] <= 8'h10 ;
			data[64388] <= 8'h10 ;
			data[64389] <= 8'h10 ;
			data[64390] <= 8'h10 ;
			data[64391] <= 8'h10 ;
			data[64392] <= 8'h10 ;
			data[64393] <= 8'h10 ;
			data[64394] <= 8'h10 ;
			data[64395] <= 8'h10 ;
			data[64396] <= 8'h10 ;
			data[64397] <= 8'h10 ;
			data[64398] <= 8'h10 ;
			data[64399] <= 8'h10 ;
			data[64400] <= 8'h10 ;
			data[64401] <= 8'h10 ;
			data[64402] <= 8'h10 ;
			data[64403] <= 8'h10 ;
			data[64404] <= 8'h10 ;
			data[64405] <= 8'h10 ;
			data[64406] <= 8'h10 ;
			data[64407] <= 8'h10 ;
			data[64408] <= 8'h10 ;
			data[64409] <= 8'h10 ;
			data[64410] <= 8'h10 ;
			data[64411] <= 8'h10 ;
			data[64412] <= 8'h10 ;
			data[64413] <= 8'h10 ;
			data[64414] <= 8'h10 ;
			data[64415] <= 8'h10 ;
			data[64416] <= 8'h10 ;
			data[64417] <= 8'h10 ;
			data[64418] <= 8'h10 ;
			data[64419] <= 8'h10 ;
			data[64420] <= 8'h10 ;
			data[64421] <= 8'h10 ;
			data[64422] <= 8'h10 ;
			data[64423] <= 8'h10 ;
			data[64424] <= 8'h10 ;
			data[64425] <= 8'h10 ;
			data[64426] <= 8'h10 ;
			data[64427] <= 8'h10 ;
			data[64428] <= 8'h10 ;
			data[64429] <= 8'h10 ;
			data[64430] <= 8'h10 ;
			data[64431] <= 8'h10 ;
			data[64432] <= 8'h10 ;
			data[64433] <= 8'h10 ;
			data[64434] <= 8'h10 ;
			data[64435] <= 8'h10 ;
			data[64436] <= 8'h10 ;
			data[64437] <= 8'h10 ;
			data[64438] <= 8'h10 ;
			data[64439] <= 8'h10 ;
			data[64440] <= 8'h10 ;
			data[64441] <= 8'h10 ;
			data[64442] <= 8'h10 ;
			data[64443] <= 8'h10 ;
			data[64444] <= 8'h10 ;
			data[64445] <= 8'h10 ;
			data[64446] <= 8'h10 ;
			data[64447] <= 8'h10 ;
			data[64448] <= 8'h10 ;
			data[64449] <= 8'h10 ;
			data[64450] <= 8'h10 ;
			data[64451] <= 8'h10 ;
			data[64452] <= 8'h10 ;
			data[64453] <= 8'h10 ;
			data[64454] <= 8'h10 ;
			data[64455] <= 8'h10 ;
			data[64456] <= 8'h10 ;
			data[64457] <= 8'h10 ;
			data[64458] <= 8'h10 ;
			data[64459] <= 8'h10 ;
			data[64460] <= 8'h10 ;
			data[64461] <= 8'h10 ;
			data[64462] <= 8'h10 ;
			data[64463] <= 8'h10 ;
			data[64464] <= 8'h10 ;
			data[64465] <= 8'h10 ;
			data[64466] <= 8'h10 ;
			data[64467] <= 8'h10 ;
			data[64468] <= 8'h10 ;
			data[64469] <= 8'h10 ;
			data[64470] <= 8'h10 ;
			data[64471] <= 8'h10 ;
			data[64472] <= 8'h10 ;
			data[64473] <= 8'h10 ;
			data[64474] <= 8'h10 ;
			data[64475] <= 8'h10 ;
			data[64476] <= 8'h10 ;
			data[64477] <= 8'h10 ;
			data[64478] <= 8'h10 ;
			data[64479] <= 8'h10 ;
			data[64480] <= 8'h10 ;
			data[64481] <= 8'h10 ;
			data[64482] <= 8'h10 ;
			data[64483] <= 8'h10 ;
			data[64484] <= 8'h10 ;
			data[64485] <= 8'h10 ;
			data[64486] <= 8'h10 ;
			data[64487] <= 8'h10 ;
			data[64488] <= 8'h10 ;
			data[64489] <= 8'h10 ;
			data[64490] <= 8'h10 ;
			data[64491] <= 8'h10 ;
			data[64492] <= 8'h10 ;
			data[64493] <= 8'h10 ;
			data[64494] <= 8'h10 ;
			data[64495] <= 8'h10 ;
			data[64496] <= 8'h10 ;
			data[64497] <= 8'h10 ;
			data[64498] <= 8'h10 ;
			data[64499] <= 8'h10 ;
			data[64500] <= 8'h10 ;
			data[64501] <= 8'h10 ;
			data[64502] <= 8'h10 ;
			data[64503] <= 8'h10 ;
			data[64504] <= 8'h10 ;
			data[64505] <= 8'h10 ;
			data[64506] <= 8'h10 ;
			data[64507] <= 8'h10 ;
			data[64508] <= 8'h10 ;
			data[64509] <= 8'h10 ;
			data[64510] <= 8'h10 ;
			data[64511] <= 8'h10 ;
			data[64512] <= 8'h10 ;
			data[64513] <= 8'h10 ;
			data[64514] <= 8'h10 ;
			data[64515] <= 8'h10 ;
			data[64516] <= 8'h10 ;
			data[64517] <= 8'h10 ;
			data[64518] <= 8'h10 ;
			data[64519] <= 8'h10 ;
			data[64520] <= 8'h10 ;
			data[64521] <= 8'h10 ;
			data[64522] <= 8'h10 ;
			data[64523] <= 8'h10 ;
			data[64524] <= 8'h10 ;
			data[64525] <= 8'h10 ;
			data[64526] <= 8'h10 ;
			data[64527] <= 8'h10 ;
			data[64528] <= 8'h10 ;
			data[64529] <= 8'h10 ;
			data[64530] <= 8'h10 ;
			data[64531] <= 8'h10 ;
			data[64532] <= 8'h10 ;
			data[64533] <= 8'h10 ;
			data[64534] <= 8'h10 ;
			data[64535] <= 8'h10 ;
			data[64536] <= 8'h10 ;
			data[64537] <= 8'h10 ;
			data[64538] <= 8'h10 ;
			data[64539] <= 8'h10 ;
			data[64540] <= 8'h10 ;
			data[64541] <= 8'h10 ;
			data[64542] <= 8'h10 ;
			data[64543] <= 8'h10 ;
			data[64544] <= 8'h10 ;
			data[64545] <= 8'h10 ;
			data[64546] <= 8'h10 ;
			data[64547] <= 8'h10 ;
			data[64548] <= 8'h10 ;
			data[64549] <= 8'h10 ;
			data[64550] <= 8'h10 ;
			data[64551] <= 8'h10 ;
			data[64552] <= 8'h10 ;
			data[64553] <= 8'h10 ;
			data[64554] <= 8'h10 ;
			data[64555] <= 8'h10 ;
			data[64556] <= 8'h10 ;
			data[64557] <= 8'h10 ;
			data[64558] <= 8'h10 ;
			data[64559] <= 8'h10 ;
			data[64560] <= 8'h10 ;
			data[64561] <= 8'h10 ;
			data[64562] <= 8'h10 ;
			data[64563] <= 8'h10 ;
			data[64564] <= 8'h10 ;
			data[64565] <= 8'h10 ;
			data[64566] <= 8'h10 ;
			data[64567] <= 8'h10 ;
			data[64568] <= 8'h10 ;
			data[64569] <= 8'h10 ;
			data[64570] <= 8'h10 ;
			data[64571] <= 8'h10 ;
			data[64572] <= 8'h10 ;
			data[64573] <= 8'h10 ;
			data[64574] <= 8'h10 ;
			data[64575] <= 8'h10 ;
			data[64576] <= 8'h10 ;
			data[64577] <= 8'h10 ;
			data[64578] <= 8'h10 ;
			data[64579] <= 8'h10 ;
			data[64580] <= 8'h10 ;
			data[64581] <= 8'h10 ;
			data[64582] <= 8'h10 ;
			data[64583] <= 8'h10 ;
			data[64584] <= 8'h10 ;
			data[64585] <= 8'h10 ;
			data[64586] <= 8'h10 ;
			data[64587] <= 8'h10 ;
			data[64588] <= 8'h10 ;
			data[64589] <= 8'h10 ;
			data[64590] <= 8'h10 ;
			data[64591] <= 8'h10 ;
			data[64592] <= 8'h10 ;
			data[64593] <= 8'h10 ;
			data[64594] <= 8'h10 ;
			data[64595] <= 8'h10 ;
			data[64596] <= 8'h10 ;
			data[64597] <= 8'h10 ;
			data[64598] <= 8'h10 ;
			data[64599] <= 8'h10 ;
			data[64600] <= 8'h10 ;
			data[64601] <= 8'h10 ;
			data[64602] <= 8'h10 ;
			data[64603] <= 8'h10 ;
			data[64604] <= 8'h10 ;
			data[64605] <= 8'h10 ;
			data[64606] <= 8'h10 ;
			data[64607] <= 8'h10 ;
			data[64608] <= 8'h10 ;
			data[64609] <= 8'h10 ;
			data[64610] <= 8'h10 ;
			data[64611] <= 8'h10 ;
			data[64612] <= 8'h10 ;
			data[64613] <= 8'h10 ;
			data[64614] <= 8'h10 ;
			data[64615] <= 8'h10 ;
			data[64616] <= 8'h10 ;
			data[64617] <= 8'h10 ;
			data[64618] <= 8'h10 ;
			data[64619] <= 8'h10 ;
			data[64620] <= 8'h10 ;
			data[64621] <= 8'h10 ;
			data[64622] <= 8'h10 ;
			data[64623] <= 8'h10 ;
			data[64624] <= 8'h10 ;
			data[64625] <= 8'h10 ;
			data[64626] <= 8'h10 ;
			data[64627] <= 8'h10 ;
			data[64628] <= 8'h10 ;
			data[64629] <= 8'h10 ;
			data[64630] <= 8'h10 ;
			data[64631] <= 8'h10 ;
			data[64632] <= 8'h10 ;
			data[64633] <= 8'h10 ;
			data[64634] <= 8'h10 ;
			data[64635] <= 8'h10 ;
			data[64636] <= 8'h10 ;
			data[64637] <= 8'h10 ;
			data[64638] <= 8'h10 ;
			data[64639] <= 8'h10 ;
			data[64640] <= 8'h10 ;
			data[64641] <= 8'h10 ;
			data[64642] <= 8'h10 ;
			data[64643] <= 8'h10 ;
			data[64644] <= 8'h10 ;
			data[64645] <= 8'h10 ;
			data[64646] <= 8'h10 ;
			data[64647] <= 8'h10 ;
			data[64648] <= 8'h10 ;
			data[64649] <= 8'h10 ;
			data[64650] <= 8'h10 ;
			data[64651] <= 8'h10 ;
			data[64652] <= 8'h10 ;
			data[64653] <= 8'h10 ;
			data[64654] <= 8'h10 ;
			data[64655] <= 8'h10 ;
			data[64656] <= 8'h10 ;
			data[64657] <= 8'h10 ;
			data[64658] <= 8'h10 ;
			data[64659] <= 8'h10 ;
			data[64660] <= 8'h10 ;
			data[64661] <= 8'h10 ;
			data[64662] <= 8'h10 ;
			data[64663] <= 8'h10 ;
			data[64664] <= 8'h10 ;
			data[64665] <= 8'h10 ;
			data[64666] <= 8'h10 ;
			data[64667] <= 8'h10 ;
			data[64668] <= 8'h10 ;
			data[64669] <= 8'h10 ;
			data[64670] <= 8'h10 ;
			data[64671] <= 8'h10 ;
			data[64672] <= 8'h10 ;
			data[64673] <= 8'h10 ;
			data[64674] <= 8'h10 ;
			data[64675] <= 8'h10 ;
			data[64676] <= 8'h10 ;
			data[64677] <= 8'h10 ;
			data[64678] <= 8'h10 ;
			data[64679] <= 8'h10 ;
			data[64680] <= 8'h10 ;
			data[64681] <= 8'h10 ;
			data[64682] <= 8'h10 ;
			data[64683] <= 8'h10 ;
			data[64684] <= 8'h10 ;
			data[64685] <= 8'h10 ;
			data[64686] <= 8'h10 ;
			data[64687] <= 8'h10 ;
			data[64688] <= 8'h10 ;
			data[64689] <= 8'h10 ;
			data[64690] <= 8'h10 ;
			data[64691] <= 8'h10 ;
			data[64692] <= 8'h10 ;
			data[64693] <= 8'h10 ;
			data[64694] <= 8'h10 ;
			data[64695] <= 8'h10 ;
			data[64696] <= 8'h10 ;
			data[64697] <= 8'h10 ;
			data[64698] <= 8'h10 ;
			data[64699] <= 8'h10 ;
			data[64700] <= 8'h10 ;
			data[64701] <= 8'h10 ;
			data[64702] <= 8'h10 ;
			data[64703] <= 8'h10 ;
			data[64704] <= 8'h10 ;
			data[64705] <= 8'h10 ;
			data[64706] <= 8'h10 ;
			data[64707] <= 8'h10 ;
			data[64708] <= 8'h10 ;
			data[64709] <= 8'h10 ;
			data[64710] <= 8'h10 ;
			data[64711] <= 8'h10 ;
			data[64712] <= 8'h10 ;
			data[64713] <= 8'h10 ;
			data[64714] <= 8'h10 ;
			data[64715] <= 8'h10 ;
			data[64716] <= 8'h10 ;
			data[64717] <= 8'h10 ;
			data[64718] <= 8'h10 ;
			data[64719] <= 8'h10 ;
			data[64720] <= 8'h10 ;
			data[64721] <= 8'h10 ;
			data[64722] <= 8'h10 ;
			data[64723] <= 8'h10 ;
			data[64724] <= 8'h10 ;
			data[64725] <= 8'h10 ;
			data[64726] <= 8'h10 ;
			data[64727] <= 8'h10 ;
			data[64728] <= 8'h10 ;
			data[64729] <= 8'h10 ;
			data[64730] <= 8'h10 ;
			data[64731] <= 8'h10 ;
			data[64732] <= 8'h10 ;
			data[64733] <= 8'h10 ;
			data[64734] <= 8'h10 ;
			data[64735] <= 8'h10 ;
			data[64736] <= 8'h10 ;
			data[64737] <= 8'h10 ;
			data[64738] <= 8'h10 ;
			data[64739] <= 8'h10 ;
			data[64740] <= 8'h10 ;
			data[64741] <= 8'h10 ;
			data[64742] <= 8'h10 ;
			data[64743] <= 8'h10 ;
			data[64744] <= 8'h10 ;
			data[64745] <= 8'h10 ;
			data[64746] <= 8'h10 ;
			data[64747] <= 8'h10 ;
			data[64748] <= 8'h10 ;
			data[64749] <= 8'h10 ;
			data[64750] <= 8'h10 ;
			data[64751] <= 8'h10 ;
			data[64752] <= 8'h10 ;
			data[64753] <= 8'h10 ;
			data[64754] <= 8'h10 ;
			data[64755] <= 8'h10 ;
			data[64756] <= 8'h10 ;
			data[64757] <= 8'h10 ;
			data[64758] <= 8'h10 ;
			data[64759] <= 8'h10 ;
			data[64760] <= 8'h10 ;
			data[64761] <= 8'h10 ;
			data[64762] <= 8'h10 ;
			data[64763] <= 8'h10 ;
			data[64764] <= 8'h10 ;
			data[64765] <= 8'h10 ;
			data[64766] <= 8'h10 ;
			data[64767] <= 8'h10 ;
			data[64768] <= 8'h10 ;
			data[64769] <= 8'h10 ;
			data[64770] <= 8'h10 ;
			data[64771] <= 8'h10 ;
			data[64772] <= 8'h10 ;
			data[64773] <= 8'h10 ;
			data[64774] <= 8'h10 ;
			data[64775] <= 8'h10 ;
			data[64776] <= 8'h10 ;
			data[64777] <= 8'h10 ;
			data[64778] <= 8'h10 ;
			data[64779] <= 8'h10 ;
			data[64780] <= 8'h10 ;
			data[64781] <= 8'h10 ;
			data[64782] <= 8'h10 ;
			data[64783] <= 8'h10 ;
			data[64784] <= 8'h10 ;
			data[64785] <= 8'h10 ;
			data[64786] <= 8'h10 ;
			data[64787] <= 8'h10 ;
			data[64788] <= 8'h10 ;
			data[64789] <= 8'h10 ;
			data[64790] <= 8'h10 ;
			data[64791] <= 8'h10 ;
			data[64792] <= 8'h10 ;
			data[64793] <= 8'h10 ;
			data[64794] <= 8'h10 ;
			data[64795] <= 8'h10 ;
			data[64796] <= 8'h10 ;
			data[64797] <= 8'h10 ;
			data[64798] <= 8'h10 ;
			data[64799] <= 8'h10 ;
			data[64800] <= 8'h10 ;
			data[64801] <= 8'h10 ;
			data[64802] <= 8'h10 ;
			data[64803] <= 8'h10 ;
			data[64804] <= 8'h10 ;
			data[64805] <= 8'h10 ;
			data[64806] <= 8'h10 ;
			data[64807] <= 8'h10 ;
			data[64808] <= 8'h10 ;
			data[64809] <= 8'h10 ;
			data[64810] <= 8'h10 ;
			data[64811] <= 8'h10 ;
			data[64812] <= 8'h10 ;
			data[64813] <= 8'h10 ;
			data[64814] <= 8'h10 ;
			data[64815] <= 8'h10 ;
			data[64816] <= 8'h10 ;
			data[64817] <= 8'h10 ;
			data[64818] <= 8'h10 ;
			data[64819] <= 8'h10 ;
			data[64820] <= 8'h10 ;
			data[64821] <= 8'h10 ;
			data[64822] <= 8'h10 ;
			data[64823] <= 8'h10 ;
			data[64824] <= 8'h10 ;
			data[64825] <= 8'h10 ;
			data[64826] <= 8'h10 ;
			data[64827] <= 8'h10 ;
			data[64828] <= 8'h10 ;
			data[64829] <= 8'h10 ;
			data[64830] <= 8'h10 ;
			data[64831] <= 8'h10 ;
			data[64832] <= 8'h10 ;
			data[64833] <= 8'h10 ;
			data[64834] <= 8'h10 ;
			data[64835] <= 8'h10 ;
			data[64836] <= 8'h10 ;
			data[64837] <= 8'h10 ;
			data[64838] <= 8'h10 ;
			data[64839] <= 8'h10 ;
			data[64840] <= 8'h10 ;
			data[64841] <= 8'h10 ;
			data[64842] <= 8'h10 ;
			data[64843] <= 8'h10 ;
			data[64844] <= 8'h10 ;
			data[64845] <= 8'h10 ;
			data[64846] <= 8'h10 ;
			data[64847] <= 8'h10 ;
			data[64848] <= 8'h10 ;
			data[64849] <= 8'h10 ;
			data[64850] <= 8'h10 ;
			data[64851] <= 8'h10 ;
			data[64852] <= 8'h10 ;
			data[64853] <= 8'h10 ;
			data[64854] <= 8'h10 ;
			data[64855] <= 8'h10 ;
			data[64856] <= 8'h10 ;
			data[64857] <= 8'h10 ;
			data[64858] <= 8'h10 ;
			data[64859] <= 8'h10 ;
			data[64860] <= 8'h10 ;
			data[64861] <= 8'h10 ;
			data[64862] <= 8'h10 ;
			data[64863] <= 8'h10 ;
			data[64864] <= 8'h10 ;
			data[64865] <= 8'h10 ;
			data[64866] <= 8'h10 ;
			data[64867] <= 8'h10 ;
			data[64868] <= 8'h10 ;
			data[64869] <= 8'h10 ;
			data[64870] <= 8'h10 ;
			data[64871] <= 8'h10 ;
			data[64872] <= 8'h10 ;
			data[64873] <= 8'h10 ;
			data[64874] <= 8'h10 ;
			data[64875] <= 8'h10 ;
			data[64876] <= 8'h10 ;
			data[64877] <= 8'h10 ;
			data[64878] <= 8'h10 ;
			data[64879] <= 8'h10 ;
			data[64880] <= 8'h10 ;
			data[64881] <= 8'h10 ;
			data[64882] <= 8'h10 ;
			data[64883] <= 8'h10 ;
			data[64884] <= 8'h10 ;
			data[64885] <= 8'h10 ;
			data[64886] <= 8'h10 ;
			data[64887] <= 8'h10 ;
			data[64888] <= 8'h10 ;
			data[64889] <= 8'h10 ;
			data[64890] <= 8'h10 ;
			data[64891] <= 8'h10 ;
			data[64892] <= 8'h10 ;
			data[64893] <= 8'h10 ;
			data[64894] <= 8'h10 ;
			data[64895] <= 8'h10 ;
			data[64896] <= 8'h10 ;
			data[64897] <= 8'h10 ;
			data[64898] <= 8'h10 ;
			data[64899] <= 8'h10 ;
			data[64900] <= 8'h10 ;
			data[64901] <= 8'h10 ;
			data[64902] <= 8'h10 ;
			data[64903] <= 8'h10 ;
			data[64904] <= 8'h10 ;
			data[64905] <= 8'h10 ;
			data[64906] <= 8'h10 ;
			data[64907] <= 8'h10 ;
			data[64908] <= 8'h10 ;
			data[64909] <= 8'h10 ;
			data[64910] <= 8'h10 ;
			data[64911] <= 8'h10 ;
			data[64912] <= 8'h10 ;
			data[64913] <= 8'h10 ;
			data[64914] <= 8'h10 ;
			data[64915] <= 8'h10 ;
			data[64916] <= 8'h10 ;
			data[64917] <= 8'h10 ;
			data[64918] <= 8'h10 ;
			data[64919] <= 8'h10 ;
			data[64920] <= 8'h10 ;
			data[64921] <= 8'h10 ;
			data[64922] <= 8'h10 ;
			data[64923] <= 8'h10 ;
			data[64924] <= 8'h10 ;
			data[64925] <= 8'h10 ;
			data[64926] <= 8'h10 ;
			data[64927] <= 8'h10 ;
			data[64928] <= 8'h10 ;
			data[64929] <= 8'h10 ;
			data[64930] <= 8'h10 ;
			data[64931] <= 8'h10 ;
			data[64932] <= 8'h10 ;
			data[64933] <= 8'h10 ;
			data[64934] <= 8'h10 ;
			data[64935] <= 8'h10 ;
			data[64936] <= 8'h10 ;
			data[64937] <= 8'h10 ;
			data[64938] <= 8'h10 ;
			data[64939] <= 8'h10 ;
			data[64940] <= 8'h10 ;
			data[64941] <= 8'h10 ;
			data[64942] <= 8'h10 ;
			data[64943] <= 8'h10 ;
			data[64944] <= 8'h10 ;
			data[64945] <= 8'h10 ;
			data[64946] <= 8'h10 ;
			data[64947] <= 8'h10 ;
			data[64948] <= 8'h10 ;
			data[64949] <= 8'h10 ;
			data[64950] <= 8'h10 ;
			data[64951] <= 8'h10 ;
			data[64952] <= 8'h10 ;
			data[64953] <= 8'h10 ;
			data[64954] <= 8'h10 ;
			data[64955] <= 8'h10 ;
			data[64956] <= 8'h10 ;
			data[64957] <= 8'h10 ;
			data[64958] <= 8'h10 ;
			data[64959] <= 8'h10 ;
			data[64960] <= 8'h10 ;
			data[64961] <= 8'h10 ;
			data[64962] <= 8'h10 ;
			data[64963] <= 8'h10 ;
			data[64964] <= 8'h10 ;
			data[64965] <= 8'h10 ;
			data[64966] <= 8'h10 ;
			data[64967] <= 8'h10 ;
			data[64968] <= 8'h10 ;
			data[64969] <= 8'h10 ;
			data[64970] <= 8'h10 ;
			data[64971] <= 8'h10 ;
			data[64972] <= 8'h10 ;
			data[64973] <= 8'h10 ;
			data[64974] <= 8'h10 ;
			data[64975] <= 8'h10 ;
			data[64976] <= 8'h10 ;
			data[64977] <= 8'h10 ;
			data[64978] <= 8'h10 ;
			data[64979] <= 8'h10 ;
			data[64980] <= 8'h10 ;
			data[64981] <= 8'h10 ;
			data[64982] <= 8'h10 ;
			data[64983] <= 8'h10 ;
			data[64984] <= 8'h10 ;
			data[64985] <= 8'h10 ;
			data[64986] <= 8'h10 ;
			data[64987] <= 8'h10 ;
			data[64988] <= 8'h10 ;
			data[64989] <= 8'h10 ;
			data[64990] <= 8'h10 ;
			data[64991] <= 8'h10 ;
			data[64992] <= 8'h10 ;
			data[64993] <= 8'h10 ;
			data[64994] <= 8'h10 ;
			data[64995] <= 8'h10 ;
			data[64996] <= 8'h10 ;
			data[64997] <= 8'h10 ;
			data[64998] <= 8'h10 ;
			data[64999] <= 8'h10 ;
			data[65000] <= 8'h10 ;
			data[65001] <= 8'h10 ;
			data[65002] <= 8'h10 ;
			data[65003] <= 8'h10 ;
			data[65004] <= 8'h10 ;
			data[65005] <= 8'h10 ;
			data[65006] <= 8'h10 ;
			data[65007] <= 8'h10 ;
			data[65008] <= 8'h10 ;
			data[65009] <= 8'h10 ;
			data[65010] <= 8'h10 ;
			data[65011] <= 8'h10 ;
			data[65012] <= 8'h10 ;
			data[65013] <= 8'h10 ;
			data[65014] <= 8'h10 ;
			data[65015] <= 8'h10 ;
			data[65016] <= 8'h10 ;
			data[65017] <= 8'h10 ;
			data[65018] <= 8'h10 ;
			data[65019] <= 8'h10 ;
			data[65020] <= 8'h10 ;
			data[65021] <= 8'h10 ;
			data[65022] <= 8'h10 ;
			data[65023] <= 8'h10 ;
			data[65024] <= 8'h10 ;
			data[65025] <= 8'h10 ;
			data[65026] <= 8'h10 ;
			data[65027] <= 8'h10 ;
			data[65028] <= 8'h10 ;
			data[65029] <= 8'h10 ;
			data[65030] <= 8'h10 ;
			data[65031] <= 8'h10 ;
			data[65032] <= 8'h10 ;
			data[65033] <= 8'h10 ;
			data[65034] <= 8'h10 ;
			data[65035] <= 8'h10 ;
			data[65036] <= 8'h10 ;
			data[65037] <= 8'h10 ;
			data[65038] <= 8'h10 ;
			data[65039] <= 8'h10 ;
			data[65040] <= 8'h10 ;
			data[65041] <= 8'h10 ;
			data[65042] <= 8'h10 ;
			data[65043] <= 8'h10 ;
			data[65044] <= 8'h10 ;
			data[65045] <= 8'h10 ;
			data[65046] <= 8'h10 ;
			data[65047] <= 8'h10 ;
			data[65048] <= 8'h10 ;
			data[65049] <= 8'h10 ;
			data[65050] <= 8'h10 ;
			data[65051] <= 8'h10 ;
			data[65052] <= 8'h10 ;
			data[65053] <= 8'h10 ;
			data[65054] <= 8'h10 ;
			data[65055] <= 8'h10 ;
			data[65056] <= 8'h10 ;
			data[65057] <= 8'h10 ;
			data[65058] <= 8'h10 ;
			data[65059] <= 8'h10 ;
			data[65060] <= 8'h10 ;
			data[65061] <= 8'h10 ;
			data[65062] <= 8'h10 ;
			data[65063] <= 8'h10 ;
			data[65064] <= 8'h10 ;
			data[65065] <= 8'h10 ;
			data[65066] <= 8'h10 ;
			data[65067] <= 8'h10 ;
			data[65068] <= 8'h10 ;
			data[65069] <= 8'h10 ;
			data[65070] <= 8'h10 ;
			data[65071] <= 8'h10 ;
			data[65072] <= 8'h10 ;
			data[65073] <= 8'h10 ;
			data[65074] <= 8'h10 ;
			data[65075] <= 8'h10 ;
			data[65076] <= 8'h10 ;
			data[65077] <= 8'h10 ;
			data[65078] <= 8'h10 ;
			data[65079] <= 8'h10 ;
			data[65080] <= 8'h10 ;
			data[65081] <= 8'h10 ;
			data[65082] <= 8'h10 ;
			data[65083] <= 8'h10 ;
			data[65084] <= 8'h10 ;
			data[65085] <= 8'h10 ;
			data[65086] <= 8'h10 ;
			data[65087] <= 8'h10 ;
			data[65088] <= 8'h10 ;
			data[65089] <= 8'h10 ;
			data[65090] <= 8'h10 ;
			data[65091] <= 8'h10 ;
			data[65092] <= 8'h10 ;
			data[65093] <= 8'h10 ;
			data[65094] <= 8'h10 ;
			data[65095] <= 8'h10 ;
			data[65096] <= 8'h10 ;
			data[65097] <= 8'h10 ;
			data[65098] <= 8'h10 ;
			data[65099] <= 8'h10 ;
			data[65100] <= 8'h10 ;
			data[65101] <= 8'h10 ;
			data[65102] <= 8'h10 ;
			data[65103] <= 8'h10 ;
			data[65104] <= 8'h10 ;
			data[65105] <= 8'h10 ;
			data[65106] <= 8'h10 ;
			data[65107] <= 8'h10 ;
			data[65108] <= 8'h10 ;
			data[65109] <= 8'h10 ;
			data[65110] <= 8'h10 ;
			data[65111] <= 8'h10 ;
			data[65112] <= 8'h10 ;
			data[65113] <= 8'h10 ;
			data[65114] <= 8'h10 ;
			data[65115] <= 8'h10 ;
			data[65116] <= 8'h10 ;
			data[65117] <= 8'h10 ;
			data[65118] <= 8'h10 ;
			data[65119] <= 8'h10 ;
			data[65120] <= 8'h10 ;
			data[65121] <= 8'h10 ;
			data[65122] <= 8'h10 ;
			data[65123] <= 8'h10 ;
			data[65124] <= 8'h10 ;
			data[65125] <= 8'h10 ;
			data[65126] <= 8'h10 ;
			data[65127] <= 8'h10 ;
			data[65128] <= 8'h10 ;
			data[65129] <= 8'h10 ;
			data[65130] <= 8'h10 ;
			data[65131] <= 8'h10 ;
			data[65132] <= 8'h10 ;
			data[65133] <= 8'h10 ;
			data[65134] <= 8'h10 ;
			data[65135] <= 8'h10 ;
			data[65136] <= 8'h10 ;
			data[65137] <= 8'h10 ;
			data[65138] <= 8'h10 ;
			data[65139] <= 8'h10 ;
			data[65140] <= 8'h10 ;
			data[65141] <= 8'h10 ;
			data[65142] <= 8'h10 ;
			data[65143] <= 8'h10 ;
			data[65144] <= 8'h10 ;
			data[65145] <= 8'h10 ;
			data[65146] <= 8'h10 ;
			data[65147] <= 8'h10 ;
			data[65148] <= 8'h10 ;
			data[65149] <= 8'h10 ;
			data[65150] <= 8'h10 ;
			data[65151] <= 8'h10 ;
			data[65152] <= 8'h10 ;
			data[65153] <= 8'h10 ;
			data[65154] <= 8'h10 ;
			data[65155] <= 8'h10 ;
			data[65156] <= 8'h10 ;
			data[65157] <= 8'h10 ;
			data[65158] <= 8'h10 ;
			data[65159] <= 8'h10 ;
			data[65160] <= 8'h10 ;
			data[65161] <= 8'h10 ;
			data[65162] <= 8'h10 ;
			data[65163] <= 8'h10 ;
			data[65164] <= 8'h10 ;
			data[65165] <= 8'h10 ;
			data[65166] <= 8'h10 ;
			data[65167] <= 8'h10 ;
			data[65168] <= 8'h10 ;
			data[65169] <= 8'h10 ;
			data[65170] <= 8'h10 ;
			data[65171] <= 8'h10 ;
			data[65172] <= 8'h10 ;
			data[65173] <= 8'h10 ;
			data[65174] <= 8'h10 ;
			data[65175] <= 8'h10 ;
			data[65176] <= 8'h10 ;
			data[65177] <= 8'h10 ;
			data[65178] <= 8'h10 ;
			data[65179] <= 8'h10 ;
			data[65180] <= 8'h10 ;
			data[65181] <= 8'h10 ;
			data[65182] <= 8'h10 ;
			data[65183] <= 8'h10 ;
			data[65184] <= 8'h10 ;
			data[65185] <= 8'h10 ;
			data[65186] <= 8'h10 ;
			data[65187] <= 8'h10 ;
			data[65188] <= 8'h10 ;
			data[65189] <= 8'h10 ;
			data[65190] <= 8'h10 ;
			data[65191] <= 8'h10 ;
			data[65192] <= 8'h10 ;
			data[65193] <= 8'h10 ;
			data[65194] <= 8'h10 ;
			data[65195] <= 8'h10 ;
			data[65196] <= 8'h10 ;
			data[65197] <= 8'h10 ;
			data[65198] <= 8'h10 ;
			data[65199] <= 8'h10 ;
			data[65200] <= 8'h10 ;
			data[65201] <= 8'h10 ;
			data[65202] <= 8'h10 ;
			data[65203] <= 8'h10 ;
			data[65204] <= 8'h10 ;
			data[65205] <= 8'h10 ;
			data[65206] <= 8'h10 ;
			data[65207] <= 8'h10 ;
			data[65208] <= 8'h10 ;
			data[65209] <= 8'h10 ;
			data[65210] <= 8'h10 ;
			data[65211] <= 8'h10 ;
			data[65212] <= 8'h10 ;
			data[65213] <= 8'h10 ;
			data[65214] <= 8'h10 ;
			data[65215] <= 8'h10 ;
			data[65216] <= 8'h10 ;
			data[65217] <= 8'h10 ;
			data[65218] <= 8'h10 ;
			data[65219] <= 8'h10 ;
			data[65220] <= 8'h10 ;
			data[65221] <= 8'h10 ;
			data[65222] <= 8'h10 ;
			data[65223] <= 8'h10 ;
			data[65224] <= 8'h10 ;
			data[65225] <= 8'h10 ;
			data[65226] <= 8'h10 ;
			data[65227] <= 8'h10 ;
			data[65228] <= 8'h10 ;
			data[65229] <= 8'h10 ;
			data[65230] <= 8'h10 ;
			data[65231] <= 8'h10 ;
			data[65232] <= 8'h10 ;
			data[65233] <= 8'h10 ;
			data[65234] <= 8'h10 ;
			data[65235] <= 8'h10 ;
			data[65236] <= 8'h10 ;
			data[65237] <= 8'h10 ;
			data[65238] <= 8'h10 ;
			data[65239] <= 8'h10 ;
			data[65240] <= 8'h10 ;
			data[65241] <= 8'h10 ;
			data[65242] <= 8'h10 ;
			data[65243] <= 8'h10 ;
			data[65244] <= 8'h10 ;
			data[65245] <= 8'h10 ;
			data[65246] <= 8'h10 ;
			data[65247] <= 8'h10 ;
			data[65248] <= 8'h10 ;
			data[65249] <= 8'h10 ;
			data[65250] <= 8'h10 ;
			data[65251] <= 8'h10 ;
			data[65252] <= 8'h10 ;
			data[65253] <= 8'h10 ;
			data[65254] <= 8'h10 ;
			data[65255] <= 8'h10 ;
			data[65256] <= 8'h10 ;
			data[65257] <= 8'h10 ;
			data[65258] <= 8'h10 ;
			data[65259] <= 8'h10 ;
			data[65260] <= 8'h10 ;
			data[65261] <= 8'h10 ;
			data[65262] <= 8'h10 ;
			data[65263] <= 8'h10 ;
			data[65264] <= 8'h10 ;
			data[65265] <= 8'h10 ;
			data[65266] <= 8'h10 ;
			data[65267] <= 8'h10 ;
			data[65268] <= 8'h10 ;
			data[65269] <= 8'h10 ;
			data[65270] <= 8'h10 ;
			data[65271] <= 8'h10 ;
			data[65272] <= 8'h10 ;
			data[65273] <= 8'h10 ;
			data[65274] <= 8'h10 ;
			data[65275] <= 8'h10 ;
			data[65276] <= 8'h10 ;
			data[65277] <= 8'h10 ;
			data[65278] <= 8'h10 ;
			data[65279] <= 8'h10 ;
			data[65280] <= 8'h10 ;
			data[65281] <= 8'h10 ;
			data[65282] <= 8'h10 ;
			data[65283] <= 8'h10 ;
			data[65284] <= 8'h10 ;
			data[65285] <= 8'h10 ;
			data[65286] <= 8'h10 ;
			data[65287] <= 8'h10 ;
			data[65288] <= 8'h10 ;
			data[65289] <= 8'h10 ;
			data[65290] <= 8'h10 ;
			data[65291] <= 8'h10 ;
			data[65292] <= 8'h10 ;
			data[65293] <= 8'h10 ;
			data[65294] <= 8'h10 ;
			data[65295] <= 8'h10 ;
			data[65296] <= 8'h10 ;
			data[65297] <= 8'h10 ;
			data[65298] <= 8'h10 ;
			data[65299] <= 8'h10 ;
			data[65300] <= 8'h10 ;
			data[65301] <= 8'h10 ;
			data[65302] <= 8'h10 ;
			data[65303] <= 8'h10 ;
			data[65304] <= 8'h10 ;
			data[65305] <= 8'h10 ;
			data[65306] <= 8'h10 ;
			data[65307] <= 8'h10 ;
			data[65308] <= 8'h10 ;
			data[65309] <= 8'h10 ;
			data[65310] <= 8'h10 ;
			data[65311] <= 8'h10 ;
			data[65312] <= 8'h10 ;
			data[65313] <= 8'h10 ;
			data[65314] <= 8'h10 ;
			data[65315] <= 8'h10 ;
			data[65316] <= 8'h10 ;
			data[65317] <= 8'h10 ;
			data[65318] <= 8'h10 ;
			data[65319] <= 8'h10 ;
			data[65320] <= 8'h10 ;
			data[65321] <= 8'h10 ;
			data[65322] <= 8'h10 ;
			data[65323] <= 8'h10 ;
			data[65324] <= 8'h10 ;
			data[65325] <= 8'h10 ;
			data[65326] <= 8'h10 ;
			data[65327] <= 8'h10 ;
			data[65328] <= 8'h10 ;
			data[65329] <= 8'h10 ;
			data[65330] <= 8'h10 ;
			data[65331] <= 8'h10 ;
			data[65332] <= 8'h10 ;
			data[65333] <= 8'h10 ;
			data[65334] <= 8'h10 ;
			data[65335] <= 8'h10 ;
			data[65336] <= 8'h10 ;
			data[65337] <= 8'h10 ;
			data[65338] <= 8'h10 ;
			data[65339] <= 8'h10 ;
			data[65340] <= 8'h10 ;
			data[65341] <= 8'h10 ;
			data[65342] <= 8'h10 ;
			data[65343] <= 8'h10 ;
			data[65344] <= 8'h10 ;
			data[65345] <= 8'h10 ;
			data[65346] <= 8'h10 ;
			data[65347] <= 8'h10 ;
			data[65348] <= 8'h10 ;
			data[65349] <= 8'h10 ;
			data[65350] <= 8'h10 ;
			data[65351] <= 8'h10 ;
			data[65352] <= 8'h10 ;
			data[65353] <= 8'h10 ;
			data[65354] <= 8'h10 ;
			data[65355] <= 8'h10 ;
			data[65356] <= 8'h10 ;
			data[65357] <= 8'h10 ;
			data[65358] <= 8'h10 ;
			data[65359] <= 8'h10 ;
			data[65360] <= 8'h10 ;
			data[65361] <= 8'h10 ;
			data[65362] <= 8'h10 ;
			data[65363] <= 8'h10 ;
			data[65364] <= 8'h10 ;
			data[65365] <= 8'h10 ;
			data[65366] <= 8'h10 ;
			data[65367] <= 8'h10 ;
			data[65368] <= 8'h10 ;
			data[65369] <= 8'h10 ;
			data[65370] <= 8'h10 ;
			data[65371] <= 8'h10 ;
			data[65372] <= 8'h10 ;
			data[65373] <= 8'h10 ;
			data[65374] <= 8'h10 ;
			data[65375] <= 8'h10 ;
			data[65376] <= 8'h10 ;
			data[65377] <= 8'h10 ;
			data[65378] <= 8'h10 ;
			data[65379] <= 8'h10 ;
			data[65380] <= 8'h10 ;
			data[65381] <= 8'h10 ;
			data[65382] <= 8'h10 ;
			data[65383] <= 8'h10 ;
			data[65384] <= 8'h10 ;
			data[65385] <= 8'h10 ;
			data[65386] <= 8'h10 ;
			data[65387] <= 8'h10 ;
			data[65388] <= 8'h10 ;
			data[65389] <= 8'h10 ;
			data[65390] <= 8'h10 ;
			data[65391] <= 8'h10 ;
			data[65392] <= 8'h10 ;
			data[65393] <= 8'h10 ;
			data[65394] <= 8'h10 ;
			data[65395] <= 8'h10 ;
			data[65396] <= 8'h10 ;
			data[65397] <= 8'h10 ;
			data[65398] <= 8'h10 ;
			data[65399] <= 8'h10 ;
			data[65400] <= 8'h10 ;
			data[65401] <= 8'h10 ;
			data[65402] <= 8'h10 ;
			data[65403] <= 8'h10 ;
			data[65404] <= 8'h10 ;
			data[65405] <= 8'h10 ;
			data[65406] <= 8'h10 ;
			data[65407] <= 8'h10 ;
			data[65408] <= 8'h10 ;
			data[65409] <= 8'h10 ;
			data[65410] <= 8'h10 ;
			data[65411] <= 8'h10 ;
			data[65412] <= 8'h10 ;
			data[65413] <= 8'h10 ;
			data[65414] <= 8'h10 ;
			data[65415] <= 8'h10 ;
			data[65416] <= 8'h10 ;
			data[65417] <= 8'h10 ;
			data[65418] <= 8'h10 ;
			data[65419] <= 8'h10 ;
			data[65420] <= 8'h10 ;
			data[65421] <= 8'h10 ;
			data[65422] <= 8'h10 ;
			data[65423] <= 8'h10 ;
			data[65424] <= 8'h10 ;
			data[65425] <= 8'h10 ;
			data[65426] <= 8'h10 ;
			data[65427] <= 8'h10 ;
			data[65428] <= 8'h10 ;
			data[65429] <= 8'h10 ;
			data[65430] <= 8'h10 ;
			data[65431] <= 8'h10 ;
			data[65432] <= 8'h10 ;
			data[65433] <= 8'h10 ;
			data[65434] <= 8'h10 ;
			data[65435] <= 8'h10 ;
			data[65436] <= 8'h10 ;
			data[65437] <= 8'h10 ;
			data[65438] <= 8'h10 ;
			data[65439] <= 8'h10 ;
			data[65440] <= 8'h10 ;
			data[65441] <= 8'h10 ;
			data[65442] <= 8'h10 ;
			data[65443] <= 8'h10 ;
			data[65444] <= 8'h10 ;
			data[65445] <= 8'h10 ;
			data[65446] <= 8'h10 ;
			data[65447] <= 8'h10 ;
			data[65448] <= 8'h10 ;
			data[65449] <= 8'h10 ;
			data[65450] <= 8'h10 ;
			data[65451] <= 8'h10 ;
			data[65452] <= 8'h10 ;
			data[65453] <= 8'h10 ;
			data[65454] <= 8'h10 ;
			data[65455] <= 8'h10 ;
			data[65456] <= 8'h10 ;
			data[65457] <= 8'h10 ;
			data[65458] <= 8'h10 ;
			data[65459] <= 8'h10 ;
			data[65460] <= 8'h10 ;
			data[65461] <= 8'h10 ;
			data[65462] <= 8'h10 ;
			data[65463] <= 8'h10 ;
			data[65464] <= 8'h10 ;
			data[65465] <= 8'h10 ;
			data[65466] <= 8'h10 ;
			data[65467] <= 8'h10 ;
			data[65468] <= 8'h10 ;
			data[65469] <= 8'h10 ;
			data[65470] <= 8'h10 ;
			data[65471] <= 8'h10 ;
			data[65472] <= 8'h10 ;
			data[65473] <= 8'h10 ;
			data[65474] <= 8'h10 ;
			data[65475] <= 8'h10 ;
			data[65476] <= 8'h10 ;
			data[65477] <= 8'h10 ;
			data[65478] <= 8'h10 ;
			data[65479] <= 8'h10 ;
			data[65480] <= 8'h10 ;
			data[65481] <= 8'h10 ;
			data[65482] <= 8'h10 ;
			data[65483] <= 8'h10 ;
			data[65484] <= 8'h10 ;
			data[65485] <= 8'h10 ;
			data[65486] <= 8'h10 ;
			data[65487] <= 8'h10 ;
			data[65488] <= 8'h10 ;
			data[65489] <= 8'h10 ;
			data[65490] <= 8'h10 ;
			data[65491] <= 8'h10 ;
			data[65492] <= 8'h10 ;
			data[65493] <= 8'h10 ;
			data[65494] <= 8'h10 ;
			data[65495] <= 8'h10 ;
			data[65496] <= 8'h10 ;
			data[65497] <= 8'h10 ;
			data[65498] <= 8'h10 ;
			data[65499] <= 8'h10 ;
			data[65500] <= 8'h10 ;
			data[65501] <= 8'h10 ;
			data[65502] <= 8'h10 ;
			data[65503] <= 8'h10 ;
			data[65504] <= 8'h10 ;
			data[65505] <= 8'h10 ;
			data[65506] <= 8'h10 ;
			data[65507] <= 8'h10 ;
			data[65508] <= 8'h10 ;
			data[65509] <= 8'h10 ;
			data[65510] <= 8'h10 ;
			data[65511] <= 8'h10 ;
			data[65512] <= 8'h10 ;
			data[65513] <= 8'h10 ;
			data[65514] <= 8'h10 ;
			data[65515] <= 8'h10 ;
			data[65516] <= 8'h10 ;
			data[65517] <= 8'h10 ;
			data[65518] <= 8'h10 ;
			data[65519] <= 8'h10 ;
			data[65520] <= 8'h10 ;
			data[65521] <= 8'h10 ;
			data[65522] <= 8'h10 ;
			data[65523] <= 8'h10 ;
			data[65524] <= 8'h10 ;
			data[65525] <= 8'h10 ;
			data[65526] <= 8'h10 ;
			data[65527] <= 8'h10 ;
			data[65528] <= 8'h10 ;
			data[65529] <= 8'h10 ;
			data[65530] <= 8'h10 ;
			data[65531] <= 8'h10 ;
			data[65532] <= 8'h10 ;
			data[65533] <= 8'h10 ;
			data[65534] <= 8'h10 ;
			data[65535] <= 8'h10 ;
			data[65536] <= 8'h10 ;
			data[65537] <= 8'h10 ;
			data[65538] <= 8'h10 ;
			data[65539] <= 8'h10 ;
			data[65540] <= 8'h10 ;
			data[65541] <= 8'h10 ;
			data[65542] <= 8'h10 ;
			data[65543] <= 8'h10 ;
			data[65544] <= 8'h10 ;
			data[65545] <= 8'h10 ;
			data[65546] <= 8'h10 ;
			data[65547] <= 8'h10 ;
			data[65548] <= 8'h10 ;
			data[65549] <= 8'h10 ;
			data[65550] <= 8'h10 ;
			data[65551] <= 8'h10 ;
			data[65552] <= 8'h10 ;
			data[65553] <= 8'h10 ;
			data[65554] <= 8'h10 ;
			data[65555] <= 8'h10 ;
			data[65556] <= 8'h10 ;
			data[65557] <= 8'h10 ;
			data[65558] <= 8'h10 ;
			data[65559] <= 8'h10 ;
			data[65560] <= 8'h10 ;
			data[65561] <= 8'h10 ;
			data[65562] <= 8'h10 ;
			data[65563] <= 8'h10 ;
			data[65564] <= 8'h10 ;
			data[65565] <= 8'h10 ;
			data[65566] <= 8'h10 ;
			data[65567] <= 8'h10 ;
			data[65568] <= 8'h10 ;
			data[65569] <= 8'h10 ;
			data[65570] <= 8'h10 ;
			data[65571] <= 8'h10 ;
			data[65572] <= 8'h10 ;
			data[65573] <= 8'h10 ;
			data[65574] <= 8'h10 ;
			data[65575] <= 8'h10 ;
			data[65576] <= 8'h10 ;
			data[65577] <= 8'h10 ;
			data[65578] <= 8'h10 ;
			data[65579] <= 8'h10 ;
			data[65580] <= 8'h10 ;
			data[65581] <= 8'h10 ;
			data[65582] <= 8'h10 ;
			data[65583] <= 8'h10 ;
			data[65584] <= 8'h10 ;
			data[65585] <= 8'h10 ;
			data[65586] <= 8'h10 ;
			data[65587] <= 8'h10 ;
			data[65588] <= 8'h10 ;
			data[65589] <= 8'h10 ;
			data[65590] <= 8'h10 ;
			data[65591] <= 8'h10 ;
			data[65592] <= 8'h10 ;
			data[65593] <= 8'h10 ;
			data[65594] <= 8'h10 ;
			data[65595] <= 8'h10 ;
			data[65596] <= 8'h10 ;
			data[65597] <= 8'h10 ;
			data[65598] <= 8'h10 ;
			data[65599] <= 8'h10 ;
			data[65600] <= 8'h10 ;
			data[65601] <= 8'h10 ;
			data[65602] <= 8'h10 ;
			data[65603] <= 8'h10 ;
			data[65604] <= 8'h10 ;
			data[65605] <= 8'h10 ;
			data[65606] <= 8'h10 ;
			data[65607] <= 8'h10 ;
			data[65608] <= 8'h10 ;
			data[65609] <= 8'h10 ;
			data[65610] <= 8'h10 ;
			data[65611] <= 8'h10 ;
			data[65612] <= 8'h10 ;
			data[65613] <= 8'h10 ;
			data[65614] <= 8'h10 ;
			data[65615] <= 8'h10 ;
			data[65616] <= 8'h10 ;
			data[65617] <= 8'h10 ;
			data[65618] <= 8'h10 ;
			data[65619] <= 8'h10 ;
			data[65620] <= 8'h10 ;
			data[65621] <= 8'h10 ;
			data[65622] <= 8'h10 ;
			data[65623] <= 8'h10 ;
			data[65624] <= 8'h10 ;
			data[65625] <= 8'h10 ;
			data[65626] <= 8'h10 ;
			data[65627] <= 8'h10 ;
			data[65628] <= 8'h10 ;
			data[65629] <= 8'h10 ;
			data[65630] <= 8'h10 ;
			data[65631] <= 8'h10 ;
			data[65632] <= 8'h10 ;
			data[65633] <= 8'h10 ;
			data[65634] <= 8'h10 ;
			data[65635] <= 8'h10 ;
			data[65636] <= 8'h10 ;
			data[65637] <= 8'h10 ;
			data[65638] <= 8'h10 ;
			data[65639] <= 8'h10 ;
			data[65640] <= 8'h10 ;
			data[65641] <= 8'h10 ;
			data[65642] <= 8'h10 ;
			data[65643] <= 8'h10 ;
			data[65644] <= 8'h10 ;
			data[65645] <= 8'h10 ;
			data[65646] <= 8'h10 ;
			data[65647] <= 8'h10 ;
			data[65648] <= 8'h10 ;
			data[65649] <= 8'h10 ;
			data[65650] <= 8'h10 ;
			data[65651] <= 8'h10 ;
			data[65652] <= 8'h10 ;
			data[65653] <= 8'h10 ;
			data[65654] <= 8'h10 ;
			data[65655] <= 8'h10 ;
			data[65656] <= 8'h10 ;
			data[65657] <= 8'h10 ;
			data[65658] <= 8'h10 ;
			data[65659] <= 8'h10 ;
			data[65660] <= 8'h10 ;
			data[65661] <= 8'h10 ;
			data[65662] <= 8'h10 ;
			data[65663] <= 8'h10 ;
			data[65664] <= 8'h10 ;
			data[65665] <= 8'h10 ;
			data[65666] <= 8'h10 ;
			data[65667] <= 8'h10 ;
			data[65668] <= 8'h10 ;
			data[65669] <= 8'h10 ;
			data[65670] <= 8'h10 ;
			data[65671] <= 8'h10 ;
			data[65672] <= 8'h10 ;
			data[65673] <= 8'h10 ;
			data[65674] <= 8'h10 ;
			data[65675] <= 8'h10 ;
			data[65676] <= 8'h10 ;
			data[65677] <= 8'h10 ;
			data[65678] <= 8'h10 ;
			data[65679] <= 8'h10 ;
			data[65680] <= 8'h10 ;
			data[65681] <= 8'h10 ;
			data[65682] <= 8'h10 ;
			data[65683] <= 8'h10 ;
			data[65684] <= 8'h10 ;
			data[65685] <= 8'h10 ;
			data[65686] <= 8'h10 ;
			data[65687] <= 8'h10 ;
			data[65688] <= 8'h10 ;
			data[65689] <= 8'h10 ;
			data[65690] <= 8'h10 ;
			data[65691] <= 8'h10 ;
			data[65692] <= 8'h10 ;
			data[65693] <= 8'h10 ;
			data[65694] <= 8'h10 ;
			data[65695] <= 8'h10 ;
			data[65696] <= 8'h10 ;
			data[65697] <= 8'h10 ;
			data[65698] <= 8'h10 ;
			data[65699] <= 8'h10 ;
			data[65700] <= 8'h10 ;
			data[65701] <= 8'h10 ;
			data[65702] <= 8'h10 ;
			data[65703] <= 8'h10 ;
			data[65704] <= 8'h10 ;
			data[65705] <= 8'h10 ;
			data[65706] <= 8'h10 ;
			data[65707] <= 8'h10 ;
			data[65708] <= 8'h10 ;
			data[65709] <= 8'h10 ;
			data[65710] <= 8'h10 ;
			data[65711] <= 8'h10 ;
			data[65712] <= 8'h10 ;
			data[65713] <= 8'h10 ;
			data[65714] <= 8'h10 ;
			data[65715] <= 8'h10 ;
			data[65716] <= 8'h10 ;
			data[65717] <= 8'h10 ;
			data[65718] <= 8'h10 ;
			data[65719] <= 8'h10 ;
			data[65720] <= 8'h10 ;
			data[65721] <= 8'h10 ;
			data[65722] <= 8'h10 ;
			data[65723] <= 8'h10 ;
			data[65724] <= 8'h10 ;
			data[65725] <= 8'h10 ;
			data[65726] <= 8'h10 ;
			data[65727] <= 8'h10 ;
			data[65728] <= 8'h10 ;
			data[65729] <= 8'h10 ;
			data[65730] <= 8'h10 ;
			data[65731] <= 8'h10 ;
			data[65732] <= 8'h10 ;
			data[65733] <= 8'h10 ;
			data[65734] <= 8'h10 ;
			data[65735] <= 8'h10 ;
			data[65736] <= 8'h10 ;
			data[65737] <= 8'h10 ;
			data[65738] <= 8'h10 ;
			data[65739] <= 8'h10 ;
			data[65740] <= 8'h10 ;
			data[65741] <= 8'h10 ;
			data[65742] <= 8'h10 ;
			data[65743] <= 8'h10 ;
			data[65744] <= 8'h10 ;
			data[65745] <= 8'h10 ;
			data[65746] <= 8'h10 ;
			data[65747] <= 8'h10 ;
			data[65748] <= 8'h10 ;
			data[65749] <= 8'h10 ;
			data[65750] <= 8'h10 ;
			data[65751] <= 8'h10 ;
			data[65752] <= 8'h10 ;
			data[65753] <= 8'h10 ;
			data[65754] <= 8'h10 ;
			data[65755] <= 8'h10 ;
			data[65756] <= 8'h10 ;
			data[65757] <= 8'h10 ;
			data[65758] <= 8'h10 ;
			data[65759] <= 8'h10 ;
			data[65760] <= 8'h10 ;
			data[65761] <= 8'h10 ;
			data[65762] <= 8'h10 ;
			data[65763] <= 8'h10 ;
			data[65764] <= 8'h10 ;
			data[65765] <= 8'h10 ;
			data[65766] <= 8'h10 ;
			data[65767] <= 8'h10 ;
			data[65768] <= 8'h10 ;
			data[65769] <= 8'h10 ;
			data[65770] <= 8'h10 ;
			data[65771] <= 8'h10 ;
			data[65772] <= 8'h10 ;
			data[65773] <= 8'h10 ;
			data[65774] <= 8'h10 ;
			data[65775] <= 8'h10 ;
			data[65776] <= 8'h10 ;
			data[65777] <= 8'h10 ;
			data[65778] <= 8'h10 ;
			data[65779] <= 8'h10 ;
			data[65780] <= 8'h10 ;
			data[65781] <= 8'h10 ;
			data[65782] <= 8'h10 ;
			data[65783] <= 8'h10 ;
			data[65784] <= 8'h10 ;
			data[65785] <= 8'h10 ;
			data[65786] <= 8'h10 ;
			data[65787] <= 8'h10 ;
			data[65788] <= 8'h10 ;
			data[65789] <= 8'h10 ;
			data[65790] <= 8'h10 ;
			data[65791] <= 8'h10 ;
			data[65792] <= 8'h10 ;
			data[65793] <= 8'h10 ;
			data[65794] <= 8'h10 ;
			data[65795] <= 8'h10 ;
			data[65796] <= 8'h10 ;
			data[65797] <= 8'h10 ;
			data[65798] <= 8'h10 ;
			data[65799] <= 8'h10 ;
			data[65800] <= 8'h10 ;
			data[65801] <= 8'h10 ;
			data[65802] <= 8'h10 ;
			data[65803] <= 8'h10 ;
			data[65804] <= 8'h10 ;
			data[65805] <= 8'h10 ;
			data[65806] <= 8'h10 ;
			data[65807] <= 8'h10 ;
			data[65808] <= 8'h10 ;
			data[65809] <= 8'h10 ;
			data[65810] <= 8'h10 ;
			data[65811] <= 8'h10 ;
			data[65812] <= 8'h10 ;
			data[65813] <= 8'h10 ;
			data[65814] <= 8'h10 ;
			data[65815] <= 8'h10 ;
			data[65816] <= 8'h10 ;
			data[65817] <= 8'h10 ;
			data[65818] <= 8'h10 ;
			data[65819] <= 8'h10 ;
			data[65820] <= 8'h10 ;
			data[65821] <= 8'h10 ;
			data[65822] <= 8'h10 ;
			data[65823] <= 8'h10 ;
			data[65824] <= 8'h10 ;
			data[65825] <= 8'h10 ;
			data[65826] <= 8'h10 ;
			data[65827] <= 8'h10 ;
			data[65828] <= 8'h10 ;
			data[65829] <= 8'h10 ;
			data[65830] <= 8'h10 ;
			data[65831] <= 8'h10 ;
			data[65832] <= 8'h10 ;
			data[65833] <= 8'h10 ;
			data[65834] <= 8'h10 ;
			data[65835] <= 8'h10 ;
			data[65836] <= 8'h10 ;
			data[65837] <= 8'h10 ;
			data[65838] <= 8'h10 ;
			data[65839] <= 8'h10 ;
			data[65840] <= 8'h10 ;
			data[65841] <= 8'h10 ;
			data[65842] <= 8'h10 ;
			data[65843] <= 8'h10 ;
			data[65844] <= 8'h10 ;
			data[65845] <= 8'h10 ;
			data[65846] <= 8'h10 ;
			data[65847] <= 8'h10 ;
			data[65848] <= 8'h10 ;
			data[65849] <= 8'h10 ;
			data[65850] <= 8'h10 ;
			data[65851] <= 8'h10 ;
			data[65852] <= 8'h10 ;
			data[65853] <= 8'h10 ;
			data[65854] <= 8'h10 ;
			data[65855] <= 8'h10 ;
			data[65856] <= 8'h10 ;
			data[65857] <= 8'h10 ;
			data[65858] <= 8'h10 ;
			data[65859] <= 8'h10 ;
			data[65860] <= 8'h10 ;
			data[65861] <= 8'h10 ;
			data[65862] <= 8'h10 ;
			data[65863] <= 8'h10 ;
			data[65864] <= 8'h10 ;
			data[65865] <= 8'h10 ;
			data[65866] <= 8'h10 ;
			data[65867] <= 8'h10 ;
			data[65868] <= 8'h10 ;
			data[65869] <= 8'h10 ;
			data[65870] <= 8'h10 ;
			data[65871] <= 8'h10 ;
			data[65872] <= 8'h10 ;
			data[65873] <= 8'h10 ;
			data[65874] <= 8'h10 ;
			data[65875] <= 8'h10 ;
			data[65876] <= 8'h10 ;
			data[65877] <= 8'h10 ;
			data[65878] <= 8'h10 ;
			data[65879] <= 8'h10 ;
			data[65880] <= 8'h10 ;
			data[65881] <= 8'h10 ;
			data[65882] <= 8'h10 ;
			data[65883] <= 8'h10 ;
			data[65884] <= 8'h10 ;
			data[65885] <= 8'h10 ;
			data[65886] <= 8'h10 ;
			data[65887] <= 8'h10 ;
			data[65888] <= 8'h10 ;
			data[65889] <= 8'h10 ;
			data[65890] <= 8'h10 ;
			data[65891] <= 8'h10 ;
			data[65892] <= 8'h10 ;
			data[65893] <= 8'h10 ;
			data[65894] <= 8'h10 ;
			data[65895] <= 8'h10 ;
			data[65896] <= 8'h10 ;
			data[65897] <= 8'h10 ;
			data[65898] <= 8'h10 ;
			data[65899] <= 8'h10 ;
			data[65900] <= 8'h10 ;
			data[65901] <= 8'h10 ;
			data[65902] <= 8'h10 ;
			data[65903] <= 8'h10 ;
			data[65904] <= 8'h10 ;
			data[65905] <= 8'h10 ;
			data[65906] <= 8'h10 ;
			data[65907] <= 8'h10 ;
			data[65908] <= 8'h10 ;
			data[65909] <= 8'h10 ;
			data[65910] <= 8'h10 ;
			data[65911] <= 8'h10 ;
			data[65912] <= 8'h10 ;
			data[65913] <= 8'h10 ;
			data[65914] <= 8'h10 ;
			data[65915] <= 8'h10 ;
			data[65916] <= 8'h10 ;
			data[65917] <= 8'h10 ;
			data[65918] <= 8'h10 ;
			data[65919] <= 8'h10 ;
			data[65920] <= 8'h10 ;
			data[65921] <= 8'h10 ;
			data[65922] <= 8'h10 ;
			data[65923] <= 8'h10 ;
			data[65924] <= 8'h10 ;
			data[65925] <= 8'h10 ;
			data[65926] <= 8'h10 ;
			data[65927] <= 8'h10 ;
			data[65928] <= 8'h10 ;
			data[65929] <= 8'h10 ;
			data[65930] <= 8'h10 ;
			data[65931] <= 8'h10 ;
			data[65932] <= 8'h10 ;
			data[65933] <= 8'h10 ;
			data[65934] <= 8'h10 ;
			data[65935] <= 8'h10 ;
			data[65936] <= 8'h10 ;
			data[65937] <= 8'h10 ;
			data[65938] <= 8'h10 ;
			data[65939] <= 8'h10 ;
			data[65940] <= 8'h10 ;
			data[65941] <= 8'h10 ;
			data[65942] <= 8'h10 ;
			data[65943] <= 8'h10 ;
			data[65944] <= 8'h10 ;
			data[65945] <= 8'h10 ;
			data[65946] <= 8'h10 ;
			data[65947] <= 8'h10 ;
			data[65948] <= 8'h10 ;
			data[65949] <= 8'h10 ;
			data[65950] <= 8'h10 ;
			data[65951] <= 8'h10 ;
			data[65952] <= 8'h10 ;
			data[65953] <= 8'h10 ;
			data[65954] <= 8'h10 ;
			data[65955] <= 8'h10 ;
			data[65956] <= 8'h10 ;
			data[65957] <= 8'h10 ;
			data[65958] <= 8'h10 ;
			data[65959] <= 8'h10 ;
			data[65960] <= 8'h10 ;
			data[65961] <= 8'h10 ;
			data[65962] <= 8'h10 ;
			data[65963] <= 8'h10 ;
			data[65964] <= 8'h10 ;
			data[65965] <= 8'h10 ;
			data[65966] <= 8'h10 ;
			data[65967] <= 8'h10 ;
			data[65968] <= 8'h10 ;
			data[65969] <= 8'h10 ;
			data[65970] <= 8'h10 ;
			data[65971] <= 8'h10 ;
			data[65972] <= 8'h10 ;
			data[65973] <= 8'h10 ;
			data[65974] <= 8'h10 ;
			data[65975] <= 8'h10 ;
			data[65976] <= 8'h10 ;
			data[65977] <= 8'h10 ;
			data[65978] <= 8'h10 ;
			data[65979] <= 8'h10 ;
			data[65980] <= 8'h10 ;
			data[65981] <= 8'h10 ;
			data[65982] <= 8'h10 ;
			data[65983] <= 8'h10 ;
			data[65984] <= 8'h10 ;
			data[65985] <= 8'h10 ;
			data[65986] <= 8'h10 ;
			data[65987] <= 8'h10 ;
			data[65988] <= 8'h10 ;
			data[65989] <= 8'h10 ;
			data[65990] <= 8'h10 ;
			data[65991] <= 8'h10 ;
			data[65992] <= 8'h10 ;
			data[65993] <= 8'h10 ;
			data[65994] <= 8'h10 ;
			data[65995] <= 8'h10 ;
			data[65996] <= 8'h10 ;
			data[65997] <= 8'h10 ;
			data[65998] <= 8'h10 ;
			data[65999] <= 8'h10 ;
			data[66000] <= 8'h10 ;
			data[66001] <= 8'h10 ;
			data[66002] <= 8'h10 ;
			data[66003] <= 8'h10 ;
			data[66004] <= 8'h10 ;
			data[66005] <= 8'h10 ;
			data[66006] <= 8'h10 ;
			data[66007] <= 8'h10 ;
			data[66008] <= 8'h10 ;
			data[66009] <= 8'h10 ;
			data[66010] <= 8'h10 ;
			data[66011] <= 8'h10 ;
			data[66012] <= 8'h10 ;
			data[66013] <= 8'h10 ;
			data[66014] <= 8'h10 ;
			data[66015] <= 8'h10 ;
			data[66016] <= 8'h10 ;
			data[66017] <= 8'h10 ;
			data[66018] <= 8'h10 ;
			data[66019] <= 8'h10 ;
			data[66020] <= 8'h10 ;
			data[66021] <= 8'h10 ;
			data[66022] <= 8'h10 ;
			data[66023] <= 8'h10 ;
			data[66024] <= 8'h10 ;
			data[66025] <= 8'h10 ;
			data[66026] <= 8'h10 ;
			data[66027] <= 8'h10 ;
			data[66028] <= 8'h10 ;
			data[66029] <= 8'h10 ;
			data[66030] <= 8'h10 ;
			data[66031] <= 8'h10 ;
			data[66032] <= 8'h10 ;
			data[66033] <= 8'h10 ;
			data[66034] <= 8'h10 ;
			data[66035] <= 8'h10 ;
			data[66036] <= 8'h10 ;
			data[66037] <= 8'h10 ;
			data[66038] <= 8'h10 ;
			data[66039] <= 8'h10 ;
			data[66040] <= 8'h10 ;
			data[66041] <= 8'h10 ;
			data[66042] <= 8'h10 ;
			data[66043] <= 8'h10 ;
			data[66044] <= 8'h10 ;
			data[66045] <= 8'h10 ;
			data[66046] <= 8'h10 ;
			data[66047] <= 8'h10 ;
			data[66048] <= 8'h10 ;
			data[66049] <= 8'h10 ;
			data[66050] <= 8'h10 ;
			data[66051] <= 8'h10 ;
			data[66052] <= 8'h10 ;
			data[66053] <= 8'h10 ;
			data[66054] <= 8'h10 ;
			data[66055] <= 8'h10 ;
			data[66056] <= 8'h10 ;
			data[66057] <= 8'h10 ;
			data[66058] <= 8'h10 ;
			data[66059] <= 8'h10 ;
			data[66060] <= 8'h10 ;
			data[66061] <= 8'h10 ;
			data[66062] <= 8'h10 ;
			data[66063] <= 8'h10 ;
			data[66064] <= 8'h10 ;
			data[66065] <= 8'h10 ;
			data[66066] <= 8'h10 ;
			data[66067] <= 8'h10 ;
			data[66068] <= 8'h10 ;
			data[66069] <= 8'h10 ;
			data[66070] <= 8'h10 ;
			data[66071] <= 8'h10 ;
			data[66072] <= 8'h10 ;
			data[66073] <= 8'h10 ;
			data[66074] <= 8'h10 ;
			data[66075] <= 8'h10 ;
			data[66076] <= 8'h10 ;
			data[66077] <= 8'h10 ;
			data[66078] <= 8'h10 ;
			data[66079] <= 8'h10 ;
			data[66080] <= 8'h10 ;
			data[66081] <= 8'h10 ;
			data[66082] <= 8'h10 ;
			data[66083] <= 8'h10 ;
			data[66084] <= 8'h10 ;
			data[66085] <= 8'h10 ;
			data[66086] <= 8'h10 ;
			data[66087] <= 8'h10 ;
			data[66088] <= 8'h10 ;
			data[66089] <= 8'h10 ;
			data[66090] <= 8'h10 ;
			data[66091] <= 8'h10 ;
			data[66092] <= 8'h10 ;
			data[66093] <= 8'h10 ;
			data[66094] <= 8'h10 ;
			data[66095] <= 8'h10 ;
			data[66096] <= 8'h10 ;
			data[66097] <= 8'h10 ;
			data[66098] <= 8'h10 ;
			data[66099] <= 8'h10 ;
			data[66100] <= 8'h10 ;
			data[66101] <= 8'h10 ;
			data[66102] <= 8'h10 ;
			data[66103] <= 8'h10 ;
			data[66104] <= 8'h10 ;
			data[66105] <= 8'h10 ;
			data[66106] <= 8'h10 ;
			data[66107] <= 8'h10 ;
			data[66108] <= 8'h10 ;
			data[66109] <= 8'h10 ;
			data[66110] <= 8'h10 ;
			data[66111] <= 8'h10 ;
			data[66112] <= 8'h10 ;
			data[66113] <= 8'h10 ;
			data[66114] <= 8'h10 ;
			data[66115] <= 8'h10 ;
			data[66116] <= 8'h10 ;
			data[66117] <= 8'h10 ;
			data[66118] <= 8'h10 ;
			data[66119] <= 8'h10 ;
			data[66120] <= 8'h10 ;
			data[66121] <= 8'h10 ;
			data[66122] <= 8'h10 ;
			data[66123] <= 8'h10 ;
			data[66124] <= 8'h10 ;
			data[66125] <= 8'h10 ;
			data[66126] <= 8'h10 ;
			data[66127] <= 8'h10 ;
			data[66128] <= 8'h10 ;
			data[66129] <= 8'h10 ;
			data[66130] <= 8'h10 ;
			data[66131] <= 8'h10 ;
			data[66132] <= 8'h10 ;
			data[66133] <= 8'h10 ;
			data[66134] <= 8'h10 ;
			data[66135] <= 8'h10 ;
			data[66136] <= 8'h10 ;
			data[66137] <= 8'h10 ;
			data[66138] <= 8'h10 ;
			data[66139] <= 8'h10 ;
			data[66140] <= 8'h10 ;
			data[66141] <= 8'h10 ;
			data[66142] <= 8'h10 ;
			data[66143] <= 8'h10 ;
			data[66144] <= 8'h10 ;
			data[66145] <= 8'h10 ;
			data[66146] <= 8'h10 ;
			data[66147] <= 8'h10 ;
			data[66148] <= 8'h10 ;
			data[66149] <= 8'h10 ;
			data[66150] <= 8'h10 ;
			data[66151] <= 8'h10 ;
			data[66152] <= 8'h10 ;
			data[66153] <= 8'h10 ;
			data[66154] <= 8'h10 ;
			data[66155] <= 8'h10 ;
			data[66156] <= 8'h10 ;
			data[66157] <= 8'h10 ;
			data[66158] <= 8'h10 ;
			data[66159] <= 8'h10 ;
			data[66160] <= 8'h10 ;
			data[66161] <= 8'h10 ;
			data[66162] <= 8'h10 ;
			data[66163] <= 8'h10 ;
			data[66164] <= 8'h10 ;
			data[66165] <= 8'h10 ;
			data[66166] <= 8'h10 ;
			data[66167] <= 8'h10 ;
			data[66168] <= 8'h10 ;
			data[66169] <= 8'h10 ;
			data[66170] <= 8'h10 ;
			data[66171] <= 8'h10 ;
			data[66172] <= 8'h10 ;
			data[66173] <= 8'h10 ;
			data[66174] <= 8'h10 ;
			data[66175] <= 8'h10 ;
			data[66176] <= 8'h10 ;
			data[66177] <= 8'h10 ;
			data[66178] <= 8'h10 ;
			data[66179] <= 8'h10 ;
			data[66180] <= 8'h10 ;
			data[66181] <= 8'h10 ;
			data[66182] <= 8'h10 ;
			data[66183] <= 8'h10 ;
			data[66184] <= 8'h10 ;
			data[66185] <= 8'h10 ;
			data[66186] <= 8'h10 ;
			data[66187] <= 8'h10 ;
			data[66188] <= 8'h10 ;
			data[66189] <= 8'h10 ;
			data[66190] <= 8'h10 ;
			data[66191] <= 8'h10 ;
			data[66192] <= 8'h10 ;
			data[66193] <= 8'h10 ;
			data[66194] <= 8'h10 ;
			data[66195] <= 8'h10 ;
			data[66196] <= 8'h10 ;
			data[66197] <= 8'h10 ;
			data[66198] <= 8'h10 ;
			data[66199] <= 8'h10 ;
			data[66200] <= 8'h10 ;
			data[66201] <= 8'h10 ;
			data[66202] <= 8'h10 ;
			data[66203] <= 8'h10 ;
			data[66204] <= 8'h10 ;
			data[66205] <= 8'h10 ;
			data[66206] <= 8'h10 ;
			data[66207] <= 8'h10 ;
			data[66208] <= 8'h10 ;
			data[66209] <= 8'h10 ;
			data[66210] <= 8'h10 ;
			data[66211] <= 8'h10 ;
			data[66212] <= 8'h10 ;
			data[66213] <= 8'h10 ;
			data[66214] <= 8'h10 ;
			data[66215] <= 8'h10 ;
			data[66216] <= 8'h10 ;
			data[66217] <= 8'h10 ;
			data[66218] <= 8'h10 ;
			data[66219] <= 8'h10 ;
			data[66220] <= 8'h10 ;
			data[66221] <= 8'h10 ;
			data[66222] <= 8'h10 ;
			data[66223] <= 8'h10 ;
			data[66224] <= 8'h10 ;
			data[66225] <= 8'h10 ;
			data[66226] <= 8'h10 ;
			data[66227] <= 8'h10 ;
			data[66228] <= 8'h10 ;
			data[66229] <= 8'h10 ;
			data[66230] <= 8'h10 ;
			data[66231] <= 8'h10 ;
			data[66232] <= 8'h10 ;
			data[66233] <= 8'h10 ;
			data[66234] <= 8'h10 ;
			data[66235] <= 8'h10 ;
			data[66236] <= 8'h10 ;
			data[66237] <= 8'h10 ;
			data[66238] <= 8'h10 ;
			data[66239] <= 8'h10 ;
			data[66240] <= 8'h10 ;
			data[66241] <= 8'h10 ;
			data[66242] <= 8'h10 ;
			data[66243] <= 8'h10 ;
			data[66244] <= 8'h10 ;
			data[66245] <= 8'h10 ;
			data[66246] <= 8'h10 ;
			data[66247] <= 8'h10 ;
			data[66248] <= 8'h10 ;
			data[66249] <= 8'h10 ;
			data[66250] <= 8'h10 ;
			data[66251] <= 8'h10 ;
			data[66252] <= 8'h10 ;
			data[66253] <= 8'h10 ;
			data[66254] <= 8'h10 ;
			data[66255] <= 8'h10 ;
			data[66256] <= 8'h10 ;
			data[66257] <= 8'h10 ;
			data[66258] <= 8'h10 ;
			data[66259] <= 8'h10 ;
			data[66260] <= 8'h10 ;
			data[66261] <= 8'h10 ;
			data[66262] <= 8'h10 ;
			data[66263] <= 8'h10 ;
			data[66264] <= 8'h10 ;
			data[66265] <= 8'h10 ;
			data[66266] <= 8'h10 ;
			data[66267] <= 8'h10 ;
			data[66268] <= 8'h10 ;
			data[66269] <= 8'h10 ;
			data[66270] <= 8'h10 ;
			data[66271] <= 8'h10 ;
			data[66272] <= 8'h10 ;
			data[66273] <= 8'h10 ;
			data[66274] <= 8'h10 ;
			data[66275] <= 8'h10 ;
			data[66276] <= 8'h10 ;
			data[66277] <= 8'h10 ;
			data[66278] <= 8'h10 ;
			data[66279] <= 8'h10 ;
			data[66280] <= 8'h10 ;
			data[66281] <= 8'h10 ;
			data[66282] <= 8'h10 ;
			data[66283] <= 8'h10 ;
			data[66284] <= 8'h10 ;
			data[66285] <= 8'h10 ;
			data[66286] <= 8'h10 ;
			data[66287] <= 8'h10 ;
			data[66288] <= 8'h10 ;
			data[66289] <= 8'h10 ;
			data[66290] <= 8'h10 ;
			data[66291] <= 8'h10 ;
			data[66292] <= 8'h10 ;
			data[66293] <= 8'h10 ;
			data[66294] <= 8'h10 ;
			data[66295] <= 8'h10 ;
			data[66296] <= 8'h10 ;
			data[66297] <= 8'h10 ;
			data[66298] <= 8'h10 ;
			data[66299] <= 8'h10 ;
			data[66300] <= 8'h10 ;
			data[66301] <= 8'h10 ;
			data[66302] <= 8'h10 ;
			data[66303] <= 8'h10 ;
			data[66304] <= 8'h10 ;
			data[66305] <= 8'h10 ;
			data[66306] <= 8'h10 ;
			data[66307] <= 8'h10 ;
			data[66308] <= 8'h10 ;
			data[66309] <= 8'h10 ;
			data[66310] <= 8'h10 ;
			data[66311] <= 8'h10 ;
			data[66312] <= 8'h10 ;
			data[66313] <= 8'h10 ;
			data[66314] <= 8'h10 ;
			data[66315] <= 8'h10 ;
			data[66316] <= 8'h10 ;
			data[66317] <= 8'h10 ;
			data[66318] <= 8'h10 ;
			data[66319] <= 8'h10 ;
			data[66320] <= 8'h10 ;
			data[66321] <= 8'h10 ;
			data[66322] <= 8'h10 ;
			data[66323] <= 8'h10 ;
			data[66324] <= 8'h10 ;
			data[66325] <= 8'h10 ;
			data[66326] <= 8'h10 ;
			data[66327] <= 8'h10 ;
			data[66328] <= 8'h10 ;
			data[66329] <= 8'h10 ;
			data[66330] <= 8'h10 ;
			data[66331] <= 8'h10 ;
			data[66332] <= 8'h10 ;
			data[66333] <= 8'h10 ;
			data[66334] <= 8'h10 ;
			data[66335] <= 8'h10 ;
			data[66336] <= 8'h10 ;
			data[66337] <= 8'h10 ;
			data[66338] <= 8'h10 ;
			data[66339] <= 8'h10 ;
			data[66340] <= 8'h10 ;
			data[66341] <= 8'h10 ;
			data[66342] <= 8'h10 ;
			data[66343] <= 8'h10 ;
			data[66344] <= 8'h10 ;
			data[66345] <= 8'h10 ;
			data[66346] <= 8'h10 ;
			data[66347] <= 8'h10 ;
			data[66348] <= 8'h10 ;
			data[66349] <= 8'h10 ;
			data[66350] <= 8'h10 ;
			data[66351] <= 8'h10 ;
			data[66352] <= 8'h10 ;
			data[66353] <= 8'h10 ;
			data[66354] <= 8'h10 ;
			data[66355] <= 8'h10 ;
			data[66356] <= 8'h10 ;
			data[66357] <= 8'h10 ;
			data[66358] <= 8'h10 ;
			data[66359] <= 8'h10 ;
			data[66360] <= 8'h10 ;
			data[66361] <= 8'h10 ;
			data[66362] <= 8'h10 ;
			data[66363] <= 8'h10 ;
			data[66364] <= 8'h10 ;
			data[66365] <= 8'h10 ;
			data[66366] <= 8'h10 ;
			data[66367] <= 8'h10 ;
			data[66368] <= 8'h10 ;
			data[66369] <= 8'h10 ;
			data[66370] <= 8'h10 ;
			data[66371] <= 8'h10 ;
			data[66372] <= 8'h10 ;
			data[66373] <= 8'h10 ;
			data[66374] <= 8'h10 ;
			data[66375] <= 8'h10 ;
			data[66376] <= 8'h10 ;
			data[66377] <= 8'h10 ;
			data[66378] <= 8'h10 ;
			data[66379] <= 8'h10 ;
			data[66380] <= 8'h10 ;
			data[66381] <= 8'h10 ;
			data[66382] <= 8'h10 ;
			data[66383] <= 8'h10 ;
			data[66384] <= 8'h10 ;
			data[66385] <= 8'h10 ;
			data[66386] <= 8'h10 ;
			data[66387] <= 8'h10 ;
			data[66388] <= 8'h10 ;
			data[66389] <= 8'h10 ;
			data[66390] <= 8'h10 ;
			data[66391] <= 8'h10 ;
			data[66392] <= 8'h10 ;
			data[66393] <= 8'h10 ;
			data[66394] <= 8'h10 ;
			data[66395] <= 8'h10 ;
			data[66396] <= 8'h10 ;
			data[66397] <= 8'h10 ;
			data[66398] <= 8'h10 ;
			data[66399] <= 8'h10 ;
			data[66400] <= 8'h10 ;
			data[66401] <= 8'h10 ;
			data[66402] <= 8'h10 ;
			data[66403] <= 8'h10 ;
			data[66404] <= 8'h10 ;
			data[66405] <= 8'h10 ;
			data[66406] <= 8'h10 ;
			data[66407] <= 8'h10 ;
			data[66408] <= 8'h10 ;
			data[66409] <= 8'h10 ;
			data[66410] <= 8'h10 ;
			data[66411] <= 8'h10 ;
			data[66412] <= 8'h10 ;
			data[66413] <= 8'h10 ;
			data[66414] <= 8'h10 ;
			data[66415] <= 8'h10 ;
			data[66416] <= 8'h10 ;
			data[66417] <= 8'h10 ;
			data[66418] <= 8'h10 ;
			data[66419] <= 8'h10 ;
			data[66420] <= 8'h10 ;
			data[66421] <= 8'h10 ;
			data[66422] <= 8'h10 ;
			data[66423] <= 8'h10 ;
			data[66424] <= 8'h10 ;
			data[66425] <= 8'h10 ;
			data[66426] <= 8'h10 ;
			data[66427] <= 8'h10 ;
			data[66428] <= 8'h10 ;
			data[66429] <= 8'h10 ;
			data[66430] <= 8'h10 ;
			data[66431] <= 8'h10 ;
			data[66432] <= 8'h10 ;
			data[66433] <= 8'h10 ;
			data[66434] <= 8'h10 ;
			data[66435] <= 8'h10 ;
			data[66436] <= 8'h10 ;
			data[66437] <= 8'h10 ;
			data[66438] <= 8'h10 ;
			data[66439] <= 8'h10 ;
			data[66440] <= 8'h10 ;
			data[66441] <= 8'h10 ;
			data[66442] <= 8'h10 ;
			data[66443] <= 8'h10 ;
			data[66444] <= 8'h10 ;
			data[66445] <= 8'h10 ;
			data[66446] <= 8'h10 ;
			data[66447] <= 8'h10 ;
			data[66448] <= 8'h10 ;
			data[66449] <= 8'h10 ;
			data[66450] <= 8'h10 ;
			data[66451] <= 8'h10 ;
			data[66452] <= 8'h10 ;
			data[66453] <= 8'h10 ;
			data[66454] <= 8'h10 ;
			data[66455] <= 8'h10 ;
			data[66456] <= 8'h10 ;
			data[66457] <= 8'h10 ;
			data[66458] <= 8'h10 ;
			data[66459] <= 8'h10 ;
			data[66460] <= 8'h10 ;
			data[66461] <= 8'h10 ;
			data[66462] <= 8'h10 ;
			data[66463] <= 8'h10 ;
			data[66464] <= 8'h10 ;
			data[66465] <= 8'h10 ;
			data[66466] <= 8'h10 ;
			data[66467] <= 8'h10 ;
			data[66468] <= 8'h10 ;
			data[66469] <= 8'h10 ;
			data[66470] <= 8'h10 ;
			data[66471] <= 8'h10 ;
			data[66472] <= 8'h10 ;
			data[66473] <= 8'h10 ;
			data[66474] <= 8'h10 ;
			data[66475] <= 8'h10 ;
			data[66476] <= 8'h10 ;
			data[66477] <= 8'h10 ;
			data[66478] <= 8'h10 ;
			data[66479] <= 8'h10 ;
			data[66480] <= 8'h10 ;
			data[66481] <= 8'h10 ;
			data[66482] <= 8'h10 ;
			data[66483] <= 8'h10 ;
			data[66484] <= 8'h10 ;
			data[66485] <= 8'h10 ;
			data[66486] <= 8'h10 ;
			data[66487] <= 8'h10 ;
			data[66488] <= 8'h10 ;
			data[66489] <= 8'h10 ;
			data[66490] <= 8'h10 ;
			data[66491] <= 8'h10 ;
			data[66492] <= 8'h10 ;
			data[66493] <= 8'h10 ;
			data[66494] <= 8'h10 ;
			data[66495] <= 8'h10 ;
			data[66496] <= 8'h10 ;
			data[66497] <= 8'h10 ;
			data[66498] <= 8'h10 ;
			data[66499] <= 8'h10 ;
			data[66500] <= 8'h10 ;
			data[66501] <= 8'h10 ;
			data[66502] <= 8'h10 ;
			data[66503] <= 8'h10 ;
			data[66504] <= 8'h10 ;
			data[66505] <= 8'h10 ;
			data[66506] <= 8'h10 ;
			data[66507] <= 8'h10 ;
			data[66508] <= 8'h10 ;
			data[66509] <= 8'h10 ;
			data[66510] <= 8'h10 ;
			data[66511] <= 8'h10 ;
			data[66512] <= 8'h10 ;
			data[66513] <= 8'h10 ;
			data[66514] <= 8'h10 ;
			data[66515] <= 8'h10 ;
			data[66516] <= 8'h10 ;
			data[66517] <= 8'h10 ;
			data[66518] <= 8'h10 ;
			data[66519] <= 8'h10 ;
			data[66520] <= 8'h10 ;
			data[66521] <= 8'h10 ;
			data[66522] <= 8'h10 ;
			data[66523] <= 8'h10 ;
			data[66524] <= 8'h10 ;
			data[66525] <= 8'h10 ;
			data[66526] <= 8'h10 ;
			data[66527] <= 8'h10 ;
			data[66528] <= 8'h10 ;
			data[66529] <= 8'h10 ;
			data[66530] <= 8'h10 ;
			data[66531] <= 8'h10 ;
			data[66532] <= 8'h10 ;
			data[66533] <= 8'h10 ;
			data[66534] <= 8'h10 ;
			data[66535] <= 8'h10 ;
			data[66536] <= 8'h10 ;
			data[66537] <= 8'h10 ;
			data[66538] <= 8'h10 ;
			data[66539] <= 8'h10 ;
			data[66540] <= 8'h10 ;
			data[66541] <= 8'h10 ;
			data[66542] <= 8'h10 ;
			data[66543] <= 8'h10 ;
			data[66544] <= 8'h10 ;
			data[66545] <= 8'h10 ;
			data[66546] <= 8'h10 ;
			data[66547] <= 8'h10 ;
			data[66548] <= 8'h10 ;
			data[66549] <= 8'h10 ;
			data[66550] <= 8'h10 ;
			data[66551] <= 8'h10 ;
			data[66552] <= 8'h10 ;
			data[66553] <= 8'h10 ;
			data[66554] <= 8'h10 ;
			data[66555] <= 8'h10 ;
			data[66556] <= 8'h10 ;
			data[66557] <= 8'h10 ;
			data[66558] <= 8'h10 ;
			data[66559] <= 8'h10 ;
			data[66560] <= 8'h10 ;
			data[66561] <= 8'h10 ;
			data[66562] <= 8'h10 ;
			data[66563] <= 8'h10 ;
			data[66564] <= 8'h10 ;
			data[66565] <= 8'h10 ;
			data[66566] <= 8'h10 ;
			data[66567] <= 8'h10 ;
			data[66568] <= 8'h10 ;
			data[66569] <= 8'h10 ;
			data[66570] <= 8'h10 ;
			data[66571] <= 8'h10 ;
			data[66572] <= 8'h10 ;
			data[66573] <= 8'h10 ;
			data[66574] <= 8'h10 ;
			data[66575] <= 8'h10 ;
			data[66576] <= 8'h10 ;
			data[66577] <= 8'h10 ;
			data[66578] <= 8'h10 ;
			data[66579] <= 8'h10 ;
			data[66580] <= 8'h10 ;
			data[66581] <= 8'h10 ;
			data[66582] <= 8'h10 ;
			data[66583] <= 8'h10 ;
			data[66584] <= 8'h10 ;
			data[66585] <= 8'h10 ;
			data[66586] <= 8'h10 ;
			data[66587] <= 8'h10 ;
			data[66588] <= 8'h10 ;
			data[66589] <= 8'h10 ;
			data[66590] <= 8'h10 ;
			data[66591] <= 8'h10 ;
			data[66592] <= 8'h10 ;
			data[66593] <= 8'h10 ;
			data[66594] <= 8'h10 ;
			data[66595] <= 8'h10 ;
			data[66596] <= 8'h10 ;
			data[66597] <= 8'h10 ;
			data[66598] <= 8'h10 ;
			data[66599] <= 8'h10 ;
			data[66600] <= 8'h10 ;
			data[66601] <= 8'h10 ;
			data[66602] <= 8'h10 ;
			data[66603] <= 8'h10 ;
			data[66604] <= 8'h10 ;
			data[66605] <= 8'h10 ;
			data[66606] <= 8'h10 ;
			data[66607] <= 8'h10 ;
			data[66608] <= 8'h10 ;
			data[66609] <= 8'h10 ;
			data[66610] <= 8'h10 ;
			data[66611] <= 8'h10 ;
			data[66612] <= 8'h10 ;
			data[66613] <= 8'h10 ;
			data[66614] <= 8'h10 ;
			data[66615] <= 8'h10 ;
			data[66616] <= 8'h10 ;
			data[66617] <= 8'h10 ;
			data[66618] <= 8'h10 ;
			data[66619] <= 8'h10 ;
			data[66620] <= 8'h10 ;
			data[66621] <= 8'h10 ;
			data[66622] <= 8'h10 ;
			data[66623] <= 8'h10 ;
			data[66624] <= 8'h10 ;
			data[66625] <= 8'h10 ;
			data[66626] <= 8'h10 ;
			data[66627] <= 8'h10 ;
			data[66628] <= 8'h10 ;
			data[66629] <= 8'h10 ;
			data[66630] <= 8'h10 ;
			data[66631] <= 8'h10 ;
			data[66632] <= 8'h10 ;
			data[66633] <= 8'h10 ;
			data[66634] <= 8'h10 ;
			data[66635] <= 8'h10 ;
			data[66636] <= 8'h10 ;
			data[66637] <= 8'h10 ;
			data[66638] <= 8'h10 ;
			data[66639] <= 8'h10 ;
			data[66640] <= 8'h10 ;
			data[66641] <= 8'h10 ;
			data[66642] <= 8'h10 ;
			data[66643] <= 8'h10 ;
			data[66644] <= 8'h10 ;
			data[66645] <= 8'h10 ;
			data[66646] <= 8'h10 ;
			data[66647] <= 8'h10 ;
			data[66648] <= 8'h10 ;
			data[66649] <= 8'h10 ;
			data[66650] <= 8'h10 ;
			data[66651] <= 8'h10 ;
			data[66652] <= 8'h10 ;
			data[66653] <= 8'h10 ;
			data[66654] <= 8'h10 ;
			data[66655] <= 8'h10 ;
			data[66656] <= 8'h10 ;
			data[66657] <= 8'h10 ;
			data[66658] <= 8'h10 ;
			data[66659] <= 8'h10 ;
			data[66660] <= 8'h10 ;
			data[66661] <= 8'h10 ;
			data[66662] <= 8'h10 ;
			data[66663] <= 8'h10 ;
			data[66664] <= 8'h10 ;
			data[66665] <= 8'h10 ;
			data[66666] <= 8'h10 ;
			data[66667] <= 8'h10 ;
			data[66668] <= 8'h10 ;
			data[66669] <= 8'h10 ;
			data[66670] <= 8'h10 ;
			data[66671] <= 8'h10 ;
			data[66672] <= 8'h10 ;
			data[66673] <= 8'h10 ;
			data[66674] <= 8'h10 ;
			data[66675] <= 8'h10 ;
			data[66676] <= 8'h10 ;
			data[66677] <= 8'h10 ;
			data[66678] <= 8'h10 ;
			data[66679] <= 8'h10 ;
			data[66680] <= 8'h10 ;
			data[66681] <= 8'h10 ;
			data[66682] <= 8'h10 ;
			data[66683] <= 8'h10 ;
			data[66684] <= 8'h10 ;
			data[66685] <= 8'h10 ;
			data[66686] <= 8'h10 ;
			data[66687] <= 8'h10 ;
			data[66688] <= 8'h10 ;
			data[66689] <= 8'h10 ;
			data[66690] <= 8'h10 ;
			data[66691] <= 8'h10 ;
			data[66692] <= 8'h10 ;
			data[66693] <= 8'h10 ;
			data[66694] <= 8'h10 ;
			data[66695] <= 8'h10 ;
			data[66696] <= 8'h10 ;
			data[66697] <= 8'h10 ;
			data[66698] <= 8'h10 ;
			data[66699] <= 8'h10 ;
			data[66700] <= 8'h10 ;
			data[66701] <= 8'h10 ;
			data[66702] <= 8'h10 ;
			data[66703] <= 8'h10 ;
			data[66704] <= 8'h10 ;
			data[66705] <= 8'h10 ;
			data[66706] <= 8'h10 ;
			data[66707] <= 8'h10 ;
			data[66708] <= 8'h10 ;
			data[66709] <= 8'h10 ;
			data[66710] <= 8'h10 ;
			data[66711] <= 8'h10 ;
			data[66712] <= 8'h10 ;
			data[66713] <= 8'h10 ;
			data[66714] <= 8'h10 ;
			data[66715] <= 8'h10 ;
			data[66716] <= 8'h10 ;
			data[66717] <= 8'h10 ;
			data[66718] <= 8'h10 ;
			data[66719] <= 8'h10 ;
			data[66720] <= 8'h10 ;
			data[66721] <= 8'h10 ;
			data[66722] <= 8'h10 ;
			data[66723] <= 8'h10 ;
			data[66724] <= 8'h10 ;
			data[66725] <= 8'h10 ;
			data[66726] <= 8'h10 ;
			data[66727] <= 8'h10 ;
			data[66728] <= 8'h10 ;
			data[66729] <= 8'h10 ;
			data[66730] <= 8'h10 ;
			data[66731] <= 8'h10 ;
			data[66732] <= 8'h10 ;
			data[66733] <= 8'h10 ;
			data[66734] <= 8'h10 ;
			data[66735] <= 8'h10 ;
			data[66736] <= 8'h10 ;
			data[66737] <= 8'h10 ;
			data[66738] <= 8'h10 ;
			data[66739] <= 8'h10 ;
			data[66740] <= 8'h10 ;
			data[66741] <= 8'h10 ;
			data[66742] <= 8'h10 ;
			data[66743] <= 8'h10 ;
			data[66744] <= 8'h10 ;
			data[66745] <= 8'h10 ;
			data[66746] <= 8'h10 ;
			data[66747] <= 8'h10 ;
			data[66748] <= 8'h10 ;
			data[66749] <= 8'h10 ;
			data[66750] <= 8'h10 ;
			data[66751] <= 8'h10 ;
			data[66752] <= 8'h10 ;
			data[66753] <= 8'h10 ;
			data[66754] <= 8'h10 ;
			data[66755] <= 8'h10 ;
			data[66756] <= 8'h10 ;
			data[66757] <= 8'h10 ;
			data[66758] <= 8'h10 ;
			data[66759] <= 8'h10 ;
			data[66760] <= 8'h10 ;
			data[66761] <= 8'h10 ;
			data[66762] <= 8'h10 ;
			data[66763] <= 8'h10 ;
			data[66764] <= 8'h10 ;
			data[66765] <= 8'h10 ;
			data[66766] <= 8'h10 ;
			data[66767] <= 8'h10 ;
			data[66768] <= 8'h10 ;
			data[66769] <= 8'h10 ;
			data[66770] <= 8'h10 ;
			data[66771] <= 8'h10 ;
			data[66772] <= 8'h10 ;
			data[66773] <= 8'h10 ;
			data[66774] <= 8'h10 ;
			data[66775] <= 8'h10 ;
			data[66776] <= 8'h10 ;
			data[66777] <= 8'h10 ;
			data[66778] <= 8'h10 ;
			data[66779] <= 8'h10 ;
			data[66780] <= 8'h10 ;
			data[66781] <= 8'h10 ;
			data[66782] <= 8'h10 ;
			data[66783] <= 8'h10 ;
			data[66784] <= 8'h10 ;
			data[66785] <= 8'h10 ;
			data[66786] <= 8'h10 ;
			data[66787] <= 8'h10 ;
			data[66788] <= 8'h10 ;
			data[66789] <= 8'h10 ;
			data[66790] <= 8'h10 ;
			data[66791] <= 8'h10 ;
			data[66792] <= 8'h10 ;
			data[66793] <= 8'h10 ;
			data[66794] <= 8'h10 ;
			data[66795] <= 8'h10 ;
			data[66796] <= 8'h10 ;
			data[66797] <= 8'h10 ;
			data[66798] <= 8'h10 ;
			data[66799] <= 8'h10 ;
			data[66800] <= 8'h10 ;
			data[66801] <= 8'h10 ;
			data[66802] <= 8'h10 ;
			data[66803] <= 8'h10 ;
			data[66804] <= 8'h10 ;
			data[66805] <= 8'h10 ;
			data[66806] <= 8'h10 ;
			data[66807] <= 8'h10 ;
			data[66808] <= 8'h10 ;
			data[66809] <= 8'h10 ;
			data[66810] <= 8'h10 ;
			data[66811] <= 8'h10 ;
			data[66812] <= 8'h10 ;
			data[66813] <= 8'h10 ;
			data[66814] <= 8'h10 ;
			data[66815] <= 8'h10 ;
			data[66816] <= 8'h10 ;
			data[66817] <= 8'h10 ;
			data[66818] <= 8'h10 ;
			data[66819] <= 8'h10 ;
			data[66820] <= 8'h10 ;
			data[66821] <= 8'h10 ;
			data[66822] <= 8'h10 ;
			data[66823] <= 8'h10 ;
			data[66824] <= 8'h10 ;
			data[66825] <= 8'h10 ;
			data[66826] <= 8'h10 ;
			data[66827] <= 8'h10 ;
			data[66828] <= 8'h10 ;
			data[66829] <= 8'h10 ;
			data[66830] <= 8'h10 ;
			data[66831] <= 8'h10 ;
			data[66832] <= 8'h10 ;
			data[66833] <= 8'h10 ;
			data[66834] <= 8'h10 ;
			data[66835] <= 8'h10 ;
			data[66836] <= 8'h10 ;
			data[66837] <= 8'h10 ;
			data[66838] <= 8'h10 ;
			data[66839] <= 8'h10 ;
			data[66840] <= 8'h10 ;
			data[66841] <= 8'h10 ;
			data[66842] <= 8'h10 ;
			data[66843] <= 8'h10 ;
			data[66844] <= 8'h10 ;
			data[66845] <= 8'h10 ;
			data[66846] <= 8'h10 ;
			data[66847] <= 8'h10 ;
			data[66848] <= 8'h10 ;
			data[66849] <= 8'h10 ;
			data[66850] <= 8'h10 ;
			data[66851] <= 8'h10 ;
			data[66852] <= 8'h10 ;
			data[66853] <= 8'h10 ;
			data[66854] <= 8'h10 ;
			data[66855] <= 8'h10 ;
			data[66856] <= 8'h10 ;
			data[66857] <= 8'h10 ;
			data[66858] <= 8'h10 ;
			data[66859] <= 8'h10 ;
			data[66860] <= 8'h10 ;
			data[66861] <= 8'h10 ;
			data[66862] <= 8'h10 ;
			data[66863] <= 8'h10 ;
			data[66864] <= 8'h10 ;
			data[66865] <= 8'h10 ;
			data[66866] <= 8'h10 ;
			data[66867] <= 8'h10 ;
			data[66868] <= 8'h10 ;
			data[66869] <= 8'h10 ;
			data[66870] <= 8'h10 ;
			data[66871] <= 8'h10 ;
			data[66872] <= 8'h10 ;
			data[66873] <= 8'h10 ;
			data[66874] <= 8'h10 ;
			data[66875] <= 8'h10 ;
			data[66876] <= 8'h10 ;
			data[66877] <= 8'h10 ;
			data[66878] <= 8'h10 ;
			data[66879] <= 8'h10 ;
			data[66880] <= 8'h10 ;
			data[66881] <= 8'h10 ;
			data[66882] <= 8'h10 ;
			data[66883] <= 8'h10 ;
			data[66884] <= 8'h10 ;
			data[66885] <= 8'h10 ;
			data[66886] <= 8'h10 ;
			data[66887] <= 8'h10 ;
			data[66888] <= 8'h10 ;
			data[66889] <= 8'h10 ;
			data[66890] <= 8'h10 ;
			data[66891] <= 8'h10 ;
			data[66892] <= 8'h10 ;
			data[66893] <= 8'h10 ;
			data[66894] <= 8'h10 ;
			data[66895] <= 8'h10 ;
			data[66896] <= 8'h10 ;
			data[66897] <= 8'h10 ;
			data[66898] <= 8'h10 ;
			data[66899] <= 8'h10 ;
			data[66900] <= 8'h10 ;
			data[66901] <= 8'h10 ;
			data[66902] <= 8'h10 ;
			data[66903] <= 8'h10 ;
			data[66904] <= 8'h10 ;
			data[66905] <= 8'h10 ;
			data[66906] <= 8'h10 ;
			data[66907] <= 8'h10 ;
			data[66908] <= 8'h10 ;
			data[66909] <= 8'h10 ;
			data[66910] <= 8'h10 ;
			data[66911] <= 8'h10 ;
			data[66912] <= 8'h10 ;
			data[66913] <= 8'h10 ;
			data[66914] <= 8'h10 ;
			data[66915] <= 8'h10 ;
			data[66916] <= 8'h10 ;
			data[66917] <= 8'h10 ;
			data[66918] <= 8'h10 ;
			data[66919] <= 8'h10 ;
			data[66920] <= 8'h10 ;
			data[66921] <= 8'h10 ;
			data[66922] <= 8'h10 ;
			data[66923] <= 8'h10 ;
			data[66924] <= 8'h10 ;
			data[66925] <= 8'h10 ;
			data[66926] <= 8'h10 ;
			data[66927] <= 8'h10 ;
			data[66928] <= 8'h10 ;
			data[66929] <= 8'h10 ;
			data[66930] <= 8'h10 ;
			data[66931] <= 8'h10 ;
			data[66932] <= 8'h10 ;
			data[66933] <= 8'h10 ;
			data[66934] <= 8'h10 ;
			data[66935] <= 8'h10 ;
			data[66936] <= 8'h10 ;
			data[66937] <= 8'h10 ;
			data[66938] <= 8'h10 ;
			data[66939] <= 8'h10 ;
			data[66940] <= 8'h10 ;
			data[66941] <= 8'h10 ;
			data[66942] <= 8'h10 ;
			data[66943] <= 8'h10 ;
			data[66944] <= 8'h10 ;
			data[66945] <= 8'h10 ;
			data[66946] <= 8'h10 ;
			data[66947] <= 8'h10 ;
			data[66948] <= 8'h10 ;
			data[66949] <= 8'h10 ;
			data[66950] <= 8'h10 ;
			data[66951] <= 8'h10 ;
			data[66952] <= 8'h10 ;
			data[66953] <= 8'h10 ;
			data[66954] <= 8'h10 ;
			data[66955] <= 8'h10 ;
			data[66956] <= 8'h10 ;
			data[66957] <= 8'h10 ;
			data[66958] <= 8'h10 ;
			data[66959] <= 8'h10 ;
			data[66960] <= 8'h10 ;
			data[66961] <= 8'h10 ;
			data[66962] <= 8'h10 ;
			data[66963] <= 8'h10 ;
			data[66964] <= 8'h10 ;
			data[66965] <= 8'h10 ;
			data[66966] <= 8'h10 ;
			data[66967] <= 8'h10 ;
			data[66968] <= 8'h10 ;
			data[66969] <= 8'h10 ;
			data[66970] <= 8'h10 ;
			data[66971] <= 8'h10 ;
			data[66972] <= 8'h10 ;
			data[66973] <= 8'h10 ;
			data[66974] <= 8'h10 ;
			data[66975] <= 8'h10 ;
			data[66976] <= 8'h10 ;
			data[66977] <= 8'h10 ;
			data[66978] <= 8'h10 ;
			data[66979] <= 8'h10 ;
			data[66980] <= 8'h10 ;
			data[66981] <= 8'h10 ;
			data[66982] <= 8'h10 ;
			data[66983] <= 8'h10 ;
			data[66984] <= 8'h10 ;
			data[66985] <= 8'h10 ;
			data[66986] <= 8'h10 ;
			data[66987] <= 8'h10 ;
			data[66988] <= 8'h10 ;
			data[66989] <= 8'h10 ;
			data[66990] <= 8'h10 ;
			data[66991] <= 8'h10 ;
			data[66992] <= 8'h10 ;
			data[66993] <= 8'h10 ;
			data[66994] <= 8'h10 ;
			data[66995] <= 8'h10 ;
			data[66996] <= 8'h10 ;
			data[66997] <= 8'h10 ;
			data[66998] <= 8'h10 ;
			data[66999] <= 8'h10 ;
			data[67000] <= 8'h10 ;
			data[67001] <= 8'h10 ;
			data[67002] <= 8'h10 ;
			data[67003] <= 8'h10 ;
			data[67004] <= 8'h10 ;
			data[67005] <= 8'h10 ;
			data[67006] <= 8'h10 ;
			data[67007] <= 8'h10 ;
			data[67008] <= 8'h10 ;
			data[67009] <= 8'h10 ;
			data[67010] <= 8'h10 ;
			data[67011] <= 8'h10 ;
			data[67012] <= 8'h10 ;
			data[67013] <= 8'h10 ;
			data[67014] <= 8'h10 ;
			data[67015] <= 8'h10 ;
			data[67016] <= 8'h10 ;
			data[67017] <= 8'h10 ;
			data[67018] <= 8'h10 ;
			data[67019] <= 8'h10 ;
			data[67020] <= 8'h10 ;
			data[67021] <= 8'h10 ;
			data[67022] <= 8'h10 ;
			data[67023] <= 8'h10 ;
			data[67024] <= 8'h10 ;
			data[67025] <= 8'h10 ;
			data[67026] <= 8'h10 ;
			data[67027] <= 8'h10 ;
			data[67028] <= 8'h10 ;
			data[67029] <= 8'h10 ;
			data[67030] <= 8'h10 ;
			data[67031] <= 8'h10 ;
			data[67032] <= 8'h10 ;
			data[67033] <= 8'h10 ;
			data[67034] <= 8'h10 ;
			data[67035] <= 8'h10 ;
			data[67036] <= 8'h10 ;
			data[67037] <= 8'h10 ;
			data[67038] <= 8'h10 ;
			data[67039] <= 8'h10 ;
			data[67040] <= 8'h10 ;
			data[67041] <= 8'h10 ;
			data[67042] <= 8'h10 ;
			data[67043] <= 8'h10 ;
			data[67044] <= 8'h10 ;
			data[67045] <= 8'h10 ;
			data[67046] <= 8'h10 ;
			data[67047] <= 8'h10 ;
			data[67048] <= 8'h10 ;
			data[67049] <= 8'h10 ;
			data[67050] <= 8'h10 ;
			data[67051] <= 8'h10 ;
			data[67052] <= 8'h10 ;
			data[67053] <= 8'h10 ;
			data[67054] <= 8'h10 ;
			data[67055] <= 8'h10 ;
			data[67056] <= 8'h10 ;
			data[67057] <= 8'h10 ;
			data[67058] <= 8'h10 ;
			data[67059] <= 8'h10 ;
			data[67060] <= 8'h10 ;
			data[67061] <= 8'h10 ;
			data[67062] <= 8'h10 ;
			data[67063] <= 8'h10 ;
			data[67064] <= 8'h10 ;
			data[67065] <= 8'h10 ;
			data[67066] <= 8'h10 ;
			data[67067] <= 8'h10 ;
			data[67068] <= 8'h10 ;
			data[67069] <= 8'h10 ;
			data[67070] <= 8'h10 ;
			data[67071] <= 8'h10 ;
			data[67072] <= 8'h10 ;
			data[67073] <= 8'h10 ;
			data[67074] <= 8'h10 ;
			data[67075] <= 8'h10 ;
			data[67076] <= 8'h10 ;
			data[67077] <= 8'h10 ;
			data[67078] <= 8'h10 ;
			data[67079] <= 8'h10 ;
			data[67080] <= 8'h10 ;
			data[67081] <= 8'h10 ;
			data[67082] <= 8'h10 ;
			data[67083] <= 8'h10 ;
			data[67084] <= 8'h10 ;
			data[67085] <= 8'h10 ;
			data[67086] <= 8'h10 ;
			data[67087] <= 8'h10 ;
			data[67088] <= 8'h10 ;
			data[67089] <= 8'h10 ;
			data[67090] <= 8'h10 ;
			data[67091] <= 8'h10 ;
			data[67092] <= 8'h10 ;
			data[67093] <= 8'h10 ;
			data[67094] <= 8'h10 ;
			data[67095] <= 8'h10 ;
			data[67096] <= 8'h10 ;
			data[67097] <= 8'h10 ;
			data[67098] <= 8'h10 ;
			data[67099] <= 8'h10 ;
			data[67100] <= 8'h10 ;
			data[67101] <= 8'h10 ;
			data[67102] <= 8'h10 ;
			data[67103] <= 8'h10 ;
			data[67104] <= 8'h10 ;
			data[67105] <= 8'h10 ;
			data[67106] <= 8'h10 ;
			data[67107] <= 8'h10 ;
			data[67108] <= 8'h10 ;
			data[67109] <= 8'h10 ;
			data[67110] <= 8'h10 ;
			data[67111] <= 8'h10 ;
			data[67112] <= 8'h10 ;
			data[67113] <= 8'h10 ;
			data[67114] <= 8'h10 ;
			data[67115] <= 8'h10 ;
			data[67116] <= 8'h10 ;
			data[67117] <= 8'h10 ;
			data[67118] <= 8'h10 ;
			data[67119] <= 8'h10 ;
			data[67120] <= 8'h10 ;
			data[67121] <= 8'h10 ;
			data[67122] <= 8'h10 ;
			data[67123] <= 8'h10 ;
			data[67124] <= 8'h10 ;
			data[67125] <= 8'h10 ;
			data[67126] <= 8'h10 ;
			data[67127] <= 8'h10 ;
			data[67128] <= 8'h10 ;
			data[67129] <= 8'h10 ;
			data[67130] <= 8'h10 ;
			data[67131] <= 8'h10 ;
			data[67132] <= 8'h10 ;
			data[67133] <= 8'h10 ;
			data[67134] <= 8'h10 ;
			data[67135] <= 8'h10 ;
			data[67136] <= 8'h10 ;
			data[67137] <= 8'h10 ;
			data[67138] <= 8'h10 ;
			data[67139] <= 8'h10 ;
			data[67140] <= 8'h10 ;
			data[67141] <= 8'h10 ;
			data[67142] <= 8'h10 ;
			data[67143] <= 8'h10 ;
			data[67144] <= 8'h10 ;
			data[67145] <= 8'h10 ;
			data[67146] <= 8'h10 ;
			data[67147] <= 8'h10 ;
			data[67148] <= 8'h10 ;
			data[67149] <= 8'h10 ;
			data[67150] <= 8'h10 ;
			data[67151] <= 8'h10 ;
			data[67152] <= 8'h10 ;
			data[67153] <= 8'h10 ;
			data[67154] <= 8'h10 ;
			data[67155] <= 8'h10 ;
			data[67156] <= 8'h10 ;
			data[67157] <= 8'h10 ;
			data[67158] <= 8'h10 ;
			data[67159] <= 8'h10 ;
			data[67160] <= 8'h10 ;
			data[67161] <= 8'h10 ;
			data[67162] <= 8'h10 ;
			data[67163] <= 8'h10 ;
			data[67164] <= 8'h10 ;
			data[67165] <= 8'h10 ;
			data[67166] <= 8'h10 ;
			data[67167] <= 8'h10 ;
			data[67168] <= 8'h10 ;
			data[67169] <= 8'h10 ;
			data[67170] <= 8'h10 ;
			data[67171] <= 8'h10 ;
			data[67172] <= 8'h10 ;
			data[67173] <= 8'h10 ;
			data[67174] <= 8'h10 ;
			data[67175] <= 8'h10 ;
			data[67176] <= 8'h10 ;
			data[67177] <= 8'h10 ;
			data[67178] <= 8'h10 ;
			data[67179] <= 8'h10 ;
			data[67180] <= 8'h10 ;
			data[67181] <= 8'h10 ;
			data[67182] <= 8'h10 ;
			data[67183] <= 8'h10 ;
			data[67184] <= 8'h10 ;
			data[67185] <= 8'h10 ;
			data[67186] <= 8'h10 ;
			data[67187] <= 8'h10 ;
			data[67188] <= 8'h10 ;
			data[67189] <= 8'h10 ;
			data[67190] <= 8'h10 ;
			data[67191] <= 8'h10 ;
			data[67192] <= 8'h10 ;
			data[67193] <= 8'h10 ;
			data[67194] <= 8'h10 ;
			data[67195] <= 8'h10 ;
			data[67196] <= 8'h10 ;
			data[67197] <= 8'h10 ;
			data[67198] <= 8'h10 ;
			data[67199] <= 8'h10 ;
			data[67200] <= 8'h10 ;
			data[67201] <= 8'h10 ;
			data[67202] <= 8'h10 ;
			data[67203] <= 8'h10 ;
			data[67204] <= 8'h10 ;
			data[67205] <= 8'h10 ;
			data[67206] <= 8'h10 ;
			data[67207] <= 8'h10 ;
			data[67208] <= 8'h10 ;
			data[67209] <= 8'h10 ;
			data[67210] <= 8'h10 ;
			data[67211] <= 8'h10 ;
			data[67212] <= 8'h10 ;
			data[67213] <= 8'h10 ;
			data[67214] <= 8'h10 ;
			data[67215] <= 8'h10 ;
			data[67216] <= 8'h10 ;
			data[67217] <= 8'h10 ;
			data[67218] <= 8'h10 ;
			data[67219] <= 8'h10 ;
			data[67220] <= 8'h10 ;
			data[67221] <= 8'h10 ;
			data[67222] <= 8'h10 ;
			data[67223] <= 8'h10 ;
			data[67224] <= 8'h10 ;
			data[67225] <= 8'h10 ;
			data[67226] <= 8'h10 ;
			data[67227] <= 8'h10 ;
			data[67228] <= 8'h10 ;
			data[67229] <= 8'h10 ;
			data[67230] <= 8'h10 ;
			data[67231] <= 8'h10 ;
			data[67232] <= 8'h10 ;
			data[67233] <= 8'h10 ;
			data[67234] <= 8'h10 ;
			data[67235] <= 8'h10 ;
			data[67236] <= 8'h10 ;
			data[67237] <= 8'h10 ;
			data[67238] <= 8'h10 ;
			data[67239] <= 8'h10 ;
			data[67240] <= 8'h10 ;
			data[67241] <= 8'h10 ;
			data[67242] <= 8'h10 ;
			data[67243] <= 8'h10 ;
			data[67244] <= 8'h10 ;
			data[67245] <= 8'h10 ;
			data[67246] <= 8'h10 ;
			data[67247] <= 8'h10 ;
			data[67248] <= 8'h10 ;
			data[67249] <= 8'h10 ;
			data[67250] <= 8'h10 ;
			data[67251] <= 8'h10 ;
			data[67252] <= 8'h10 ;
			data[67253] <= 8'h10 ;
			data[67254] <= 8'h10 ;
			data[67255] <= 8'h10 ;
			data[67256] <= 8'h10 ;
			data[67257] <= 8'h10 ;
			data[67258] <= 8'h10 ;
			data[67259] <= 8'h10 ;
			data[67260] <= 8'h10 ;
			data[67261] <= 8'h10 ;
			data[67262] <= 8'h10 ;
			data[67263] <= 8'h10 ;
			data[67264] <= 8'h10 ;
			data[67265] <= 8'h10 ;
			data[67266] <= 8'h10 ;
			data[67267] <= 8'h10 ;
			data[67268] <= 8'h10 ;
			data[67269] <= 8'h10 ;
			data[67270] <= 8'h10 ;
			data[67271] <= 8'h10 ;
			data[67272] <= 8'h10 ;
			data[67273] <= 8'h10 ;
			data[67274] <= 8'h10 ;
			data[67275] <= 8'h10 ;
			data[67276] <= 8'h10 ;
			data[67277] <= 8'h10 ;
			data[67278] <= 8'h10 ;
			data[67279] <= 8'h10 ;
			data[67280] <= 8'h10 ;
			data[67281] <= 8'h10 ;
			data[67282] <= 8'h10 ;
			data[67283] <= 8'h10 ;
			data[67284] <= 8'h10 ;
			data[67285] <= 8'h10 ;
			data[67286] <= 8'h10 ;
			data[67287] <= 8'h10 ;
			data[67288] <= 8'h10 ;
			data[67289] <= 8'h10 ;
			data[67290] <= 8'h10 ;
			data[67291] <= 8'h10 ;
			data[67292] <= 8'h10 ;
			data[67293] <= 8'h10 ;
			data[67294] <= 8'h10 ;
			data[67295] <= 8'h10 ;
			data[67296] <= 8'h10 ;
			data[67297] <= 8'h10 ;
			data[67298] <= 8'h10 ;
			data[67299] <= 8'h10 ;
			data[67300] <= 8'h10 ;
			data[67301] <= 8'h10 ;
			data[67302] <= 8'h10 ;
			data[67303] <= 8'h10 ;
			data[67304] <= 8'h10 ;
			data[67305] <= 8'h10 ;
			data[67306] <= 8'h10 ;
			data[67307] <= 8'h10 ;
			data[67308] <= 8'h10 ;
			data[67309] <= 8'h10 ;
			data[67310] <= 8'h10 ;
			data[67311] <= 8'h10 ;
			data[67312] <= 8'h10 ;
			data[67313] <= 8'h10 ;
			data[67314] <= 8'h10 ;
			data[67315] <= 8'h10 ;
			data[67316] <= 8'h10 ;
			data[67317] <= 8'h10 ;
			data[67318] <= 8'h10 ;
			data[67319] <= 8'h10 ;
			data[67320] <= 8'h10 ;
			data[67321] <= 8'h10 ;
			data[67322] <= 8'h10 ;
			data[67323] <= 8'h10 ;
			data[67324] <= 8'h10 ;
			data[67325] <= 8'h10 ;
			data[67326] <= 8'h10 ;
			data[67327] <= 8'h10 ;
			data[67328] <= 8'h10 ;
			data[67329] <= 8'h10 ;
			data[67330] <= 8'h10 ;
			data[67331] <= 8'h10 ;
			data[67332] <= 8'h10 ;
			data[67333] <= 8'h10 ;
			data[67334] <= 8'h10 ;
			data[67335] <= 8'h10 ;
			data[67336] <= 8'h10 ;
			data[67337] <= 8'h10 ;
			data[67338] <= 8'h10 ;
			data[67339] <= 8'h10 ;
			data[67340] <= 8'h10 ;
			data[67341] <= 8'h10 ;
			data[67342] <= 8'h10 ;
			data[67343] <= 8'h10 ;
			data[67344] <= 8'h10 ;
			data[67345] <= 8'h10 ;
			data[67346] <= 8'h10 ;
			data[67347] <= 8'h10 ;
			data[67348] <= 8'h10 ;
			data[67349] <= 8'h10 ;
			data[67350] <= 8'h10 ;
			data[67351] <= 8'h10 ;
			data[67352] <= 8'h10 ;
			data[67353] <= 8'h10 ;
			data[67354] <= 8'h10 ;
			data[67355] <= 8'h10 ;
			data[67356] <= 8'h10 ;
			data[67357] <= 8'h10 ;
			data[67358] <= 8'h10 ;
			data[67359] <= 8'h10 ;
			data[67360] <= 8'h10 ;
			data[67361] <= 8'h10 ;
			data[67362] <= 8'h10 ;
			data[67363] <= 8'h10 ;
			data[67364] <= 8'h10 ;
			data[67365] <= 8'h10 ;
			data[67366] <= 8'h10 ;
			data[67367] <= 8'h10 ;
			data[67368] <= 8'h10 ;
			data[67369] <= 8'h10 ;
			data[67370] <= 8'h10 ;
			data[67371] <= 8'h10 ;
			data[67372] <= 8'h10 ;
			data[67373] <= 8'h10 ;
			data[67374] <= 8'h10 ;
			data[67375] <= 8'h10 ;
			data[67376] <= 8'h10 ;
			data[67377] <= 8'h10 ;
			data[67378] <= 8'h10 ;
			data[67379] <= 8'h10 ;
			data[67380] <= 8'h10 ;
			data[67381] <= 8'h10 ;
			data[67382] <= 8'h10 ;
			data[67383] <= 8'h10 ;
			data[67384] <= 8'h10 ;
			data[67385] <= 8'h10 ;
			data[67386] <= 8'h10 ;
			data[67387] <= 8'h10 ;
			data[67388] <= 8'h10 ;
			data[67389] <= 8'h10 ;
			data[67390] <= 8'h10 ;
			data[67391] <= 8'h10 ;
			data[67392] <= 8'h10 ;
			data[67393] <= 8'h10 ;
			data[67394] <= 8'h10 ;
			data[67395] <= 8'h10 ;
			data[67396] <= 8'h10 ;
			data[67397] <= 8'h10 ;
			data[67398] <= 8'h10 ;
			data[67399] <= 8'h10 ;
			data[67400] <= 8'h10 ;
			data[67401] <= 8'h10 ;
			data[67402] <= 8'h10 ;
			data[67403] <= 8'h10 ;
			data[67404] <= 8'h10 ;
			data[67405] <= 8'h10 ;
			data[67406] <= 8'h10 ;
			data[67407] <= 8'h10 ;
			data[67408] <= 8'h10 ;
			data[67409] <= 8'h10 ;
			data[67410] <= 8'h10 ;
			data[67411] <= 8'h10 ;
			data[67412] <= 8'h10 ;
			data[67413] <= 8'h10 ;
			data[67414] <= 8'h10 ;
			data[67415] <= 8'h10 ;
			data[67416] <= 8'h10 ;
			data[67417] <= 8'h10 ;
			data[67418] <= 8'h10 ;
			data[67419] <= 8'h10 ;
			data[67420] <= 8'h10 ;
			data[67421] <= 8'h10 ;
			data[67422] <= 8'h10 ;
			data[67423] <= 8'h10 ;
			data[67424] <= 8'h10 ;
			data[67425] <= 8'h10 ;
			data[67426] <= 8'h10 ;
			data[67427] <= 8'h10 ;
			data[67428] <= 8'h10 ;
			data[67429] <= 8'h10 ;
			data[67430] <= 8'h10 ;
			data[67431] <= 8'h10 ;
			data[67432] <= 8'h10 ;
			data[67433] <= 8'h10 ;
			data[67434] <= 8'h10 ;
			data[67435] <= 8'h10 ;
			data[67436] <= 8'h10 ;
			data[67437] <= 8'h10 ;
			data[67438] <= 8'h10 ;
			data[67439] <= 8'h10 ;
			data[67440] <= 8'h10 ;
			data[67441] <= 8'h10 ;
			data[67442] <= 8'h10 ;
			data[67443] <= 8'h10 ;
			data[67444] <= 8'h10 ;
			data[67445] <= 8'h10 ;
			data[67446] <= 8'h10 ;
			data[67447] <= 8'h10 ;
			data[67448] <= 8'h10 ;
			data[67449] <= 8'h10 ;
			data[67450] <= 8'h10 ;
			data[67451] <= 8'h10 ;
			data[67452] <= 8'h10 ;
			data[67453] <= 8'h10 ;
			data[67454] <= 8'h10 ;
			data[67455] <= 8'h10 ;
			data[67456] <= 8'h10 ;
			data[67457] <= 8'h10 ;
			data[67458] <= 8'h10 ;
			data[67459] <= 8'h10 ;
			data[67460] <= 8'h10 ;
			data[67461] <= 8'h10 ;
			data[67462] <= 8'h10 ;
			data[67463] <= 8'h10 ;
			data[67464] <= 8'h10 ;
			data[67465] <= 8'h10 ;
			data[67466] <= 8'h10 ;
			data[67467] <= 8'h10 ;
			data[67468] <= 8'h10 ;
			data[67469] <= 8'h10 ;
			data[67470] <= 8'h10 ;
			data[67471] <= 8'h10 ;
			data[67472] <= 8'h10 ;
			data[67473] <= 8'h10 ;
			data[67474] <= 8'h10 ;
			data[67475] <= 8'h10 ;
			data[67476] <= 8'h10 ;
			data[67477] <= 8'h10 ;
			data[67478] <= 8'h10 ;
			data[67479] <= 8'h10 ;
			data[67480] <= 8'h10 ;
			data[67481] <= 8'h10 ;
			data[67482] <= 8'h10 ;
			data[67483] <= 8'h10 ;
			data[67484] <= 8'h10 ;
			data[67485] <= 8'h10 ;
			data[67486] <= 8'h10 ;
			data[67487] <= 8'h10 ;
			data[67488] <= 8'h10 ;
			data[67489] <= 8'h10 ;
			data[67490] <= 8'h10 ;
			data[67491] <= 8'h10 ;
			data[67492] <= 8'h10 ;
			data[67493] <= 8'h10 ;
			data[67494] <= 8'h10 ;
			data[67495] <= 8'h10 ;
			data[67496] <= 8'h10 ;
			data[67497] <= 8'h10 ;
			data[67498] <= 8'h10 ;
			data[67499] <= 8'h10 ;
			data[67500] <= 8'h10 ;
			data[67501] <= 8'h10 ;
			data[67502] <= 8'h10 ;
			data[67503] <= 8'h10 ;
			data[67504] <= 8'h10 ;
			data[67505] <= 8'h10 ;
			data[67506] <= 8'h10 ;
			data[67507] <= 8'h10 ;
			data[67508] <= 8'h10 ;
			data[67509] <= 8'h10 ;
			data[67510] <= 8'h10 ;
			data[67511] <= 8'h10 ;
			data[67512] <= 8'h10 ;
			data[67513] <= 8'h10 ;
			data[67514] <= 8'h10 ;
			data[67515] <= 8'h10 ;
			data[67516] <= 8'h10 ;
			data[67517] <= 8'h10 ;
			data[67518] <= 8'h10 ;
			data[67519] <= 8'h10 ;
			data[67520] <= 8'h10 ;
			data[67521] <= 8'h10 ;
			data[67522] <= 8'h10 ;
			data[67523] <= 8'h10 ;
			data[67524] <= 8'h10 ;
			data[67525] <= 8'h10 ;
			data[67526] <= 8'h10 ;
			data[67527] <= 8'h10 ;
			data[67528] <= 8'h10 ;
			data[67529] <= 8'h10 ;
			data[67530] <= 8'h10 ;
			data[67531] <= 8'h10 ;
			data[67532] <= 8'h10 ;
			data[67533] <= 8'h10 ;
			data[67534] <= 8'h10 ;
			data[67535] <= 8'h10 ;
			data[67536] <= 8'h10 ;
			data[67537] <= 8'h10 ;
			data[67538] <= 8'h10 ;
			data[67539] <= 8'h10 ;
			data[67540] <= 8'h10 ;
			data[67541] <= 8'h10 ;
			data[67542] <= 8'h10 ;
			data[67543] <= 8'h10 ;
			data[67544] <= 8'h10 ;
			data[67545] <= 8'h10 ;
			data[67546] <= 8'h10 ;
			data[67547] <= 8'h10 ;
			data[67548] <= 8'h10 ;
			data[67549] <= 8'h10 ;
			data[67550] <= 8'h10 ;
			data[67551] <= 8'h10 ;
			data[67552] <= 8'h10 ;
			data[67553] <= 8'h10 ;
			data[67554] <= 8'h10 ;
			data[67555] <= 8'h10 ;
			data[67556] <= 8'h10 ;
			data[67557] <= 8'h10 ;
			data[67558] <= 8'h10 ;
			data[67559] <= 8'h10 ;
			data[67560] <= 8'h10 ;
			data[67561] <= 8'h10 ;
			data[67562] <= 8'h10 ;
			data[67563] <= 8'h10 ;
			data[67564] <= 8'h10 ;
			data[67565] <= 8'h10 ;
			data[67566] <= 8'h10 ;
			data[67567] <= 8'h10 ;
			data[67568] <= 8'h10 ;
			data[67569] <= 8'h10 ;
			data[67570] <= 8'h10 ;
			data[67571] <= 8'h10 ;
			data[67572] <= 8'h10 ;
			data[67573] <= 8'h10 ;
			data[67574] <= 8'h10 ;
			data[67575] <= 8'h10 ;
			data[67576] <= 8'h10 ;
			data[67577] <= 8'h10 ;
			data[67578] <= 8'h10 ;
			data[67579] <= 8'h10 ;
			data[67580] <= 8'h10 ;
			data[67581] <= 8'h10 ;
			data[67582] <= 8'h10 ;
			data[67583] <= 8'h10 ;
			data[67584] <= 8'h10 ;
			data[67585] <= 8'h10 ;
			data[67586] <= 8'h10 ;
			data[67587] <= 8'h10 ;
			data[67588] <= 8'h10 ;
			data[67589] <= 8'h10 ;
			data[67590] <= 8'h10 ;
			data[67591] <= 8'h10 ;
			data[67592] <= 8'h10 ;
			data[67593] <= 8'h10 ;
			data[67594] <= 8'h10 ;
			data[67595] <= 8'h10 ;
			data[67596] <= 8'h10 ;
			data[67597] <= 8'h10 ;
			data[67598] <= 8'h10 ;
			data[67599] <= 8'h10 ;
			data[67600] <= 8'h10 ;
			data[67601] <= 8'h10 ;
			data[67602] <= 8'h10 ;
			data[67603] <= 8'h10 ;
			data[67604] <= 8'h10 ;
			data[67605] <= 8'h10 ;
			data[67606] <= 8'h10 ;
			data[67607] <= 8'h10 ;
			data[67608] <= 8'h10 ;
			data[67609] <= 8'h10 ;
			data[67610] <= 8'h10 ;
			data[67611] <= 8'h10 ;
			data[67612] <= 8'h10 ;
			data[67613] <= 8'h10 ;
			data[67614] <= 8'h10 ;
			data[67615] <= 8'h10 ;
			data[67616] <= 8'h10 ;
			data[67617] <= 8'h10 ;
			data[67618] <= 8'h10 ;
			data[67619] <= 8'h10 ;
			data[67620] <= 8'h10 ;
			data[67621] <= 8'h10 ;
			data[67622] <= 8'h10 ;
			data[67623] <= 8'h10 ;
			data[67624] <= 8'h10 ;
			data[67625] <= 8'h10 ;
			data[67626] <= 8'h10 ;
			data[67627] <= 8'h10 ;
			data[67628] <= 8'h10 ;
			data[67629] <= 8'h10 ;
			data[67630] <= 8'h10 ;
			data[67631] <= 8'h10 ;
			data[67632] <= 8'h10 ;
			data[67633] <= 8'h10 ;
			data[67634] <= 8'h10 ;
			data[67635] <= 8'h10 ;
			data[67636] <= 8'h10 ;
			data[67637] <= 8'h10 ;
			data[67638] <= 8'h10 ;
			data[67639] <= 8'h10 ;
			data[67640] <= 8'h10 ;
			data[67641] <= 8'h10 ;
			data[67642] <= 8'h10 ;
			data[67643] <= 8'h10 ;
			data[67644] <= 8'h10 ;
			data[67645] <= 8'h10 ;
			data[67646] <= 8'h10 ;
			data[67647] <= 8'h10 ;
			data[67648] <= 8'h10 ;
			data[67649] <= 8'h10 ;
			data[67650] <= 8'h10 ;
			data[67651] <= 8'h10 ;
			data[67652] <= 8'h10 ;
			data[67653] <= 8'h10 ;
			data[67654] <= 8'h10 ;
			data[67655] <= 8'h10 ;
			data[67656] <= 8'h10 ;
			data[67657] <= 8'h10 ;
			data[67658] <= 8'h10 ;
			data[67659] <= 8'h10 ;
			data[67660] <= 8'h10 ;
			data[67661] <= 8'h10 ;
			data[67662] <= 8'h10 ;
			data[67663] <= 8'h10 ;
			data[67664] <= 8'h10 ;
			data[67665] <= 8'h10 ;
			data[67666] <= 8'h10 ;
			data[67667] <= 8'h10 ;
			data[67668] <= 8'h10 ;
			data[67669] <= 8'h10 ;
			data[67670] <= 8'h10 ;
			data[67671] <= 8'h10 ;
			data[67672] <= 8'h10 ;
			data[67673] <= 8'h10 ;
			data[67674] <= 8'h10 ;
			data[67675] <= 8'h10 ;
			data[67676] <= 8'h10 ;
			data[67677] <= 8'h10 ;
			data[67678] <= 8'h10 ;
			data[67679] <= 8'h10 ;
			data[67680] <= 8'h10 ;
			data[67681] <= 8'h10 ;
			data[67682] <= 8'h10 ;
			data[67683] <= 8'h10 ;
			data[67684] <= 8'h10 ;
			data[67685] <= 8'h10 ;
			data[67686] <= 8'h10 ;
			data[67687] <= 8'h10 ;
			data[67688] <= 8'h10 ;
			data[67689] <= 8'h10 ;
			data[67690] <= 8'h10 ;
			data[67691] <= 8'h10 ;
			data[67692] <= 8'h10 ;
			data[67693] <= 8'h10 ;
			data[67694] <= 8'h10 ;
			data[67695] <= 8'h10 ;
			data[67696] <= 8'h10 ;
			data[67697] <= 8'h10 ;
			data[67698] <= 8'h10 ;
			data[67699] <= 8'h10 ;
			data[67700] <= 8'h10 ;
			data[67701] <= 8'h10 ;
			data[67702] <= 8'h10 ;
			data[67703] <= 8'h10 ;
			data[67704] <= 8'h10 ;
			data[67705] <= 8'h10 ;
			data[67706] <= 8'h10 ;
			data[67707] <= 8'h10 ;
			data[67708] <= 8'h10 ;
			data[67709] <= 8'h10 ;
			data[67710] <= 8'h10 ;
			data[67711] <= 8'h10 ;
			data[67712] <= 8'h10 ;
			data[67713] <= 8'h10 ;
			data[67714] <= 8'h10 ;
			data[67715] <= 8'h10 ;
			data[67716] <= 8'h10 ;
			data[67717] <= 8'h10 ;
			data[67718] <= 8'h10 ;
			data[67719] <= 8'h10 ;
			data[67720] <= 8'h10 ;
			data[67721] <= 8'h10 ;
			data[67722] <= 8'h10 ;
			data[67723] <= 8'h10 ;
			data[67724] <= 8'h10 ;
			data[67725] <= 8'h10 ;
			data[67726] <= 8'h10 ;
			data[67727] <= 8'h10 ;
			data[67728] <= 8'h10 ;
			data[67729] <= 8'h10 ;
			data[67730] <= 8'h10 ;
			data[67731] <= 8'h10 ;
			data[67732] <= 8'h10 ;
			data[67733] <= 8'h10 ;
			data[67734] <= 8'h10 ;
			data[67735] <= 8'h10 ;
			data[67736] <= 8'h10 ;
			data[67737] <= 8'h10 ;
			data[67738] <= 8'h10 ;
			data[67739] <= 8'h10 ;
			data[67740] <= 8'h10 ;
			data[67741] <= 8'h10 ;
			data[67742] <= 8'h10 ;
			data[67743] <= 8'h10 ;
			data[67744] <= 8'h10 ;
			data[67745] <= 8'h10 ;
			data[67746] <= 8'h10 ;
			data[67747] <= 8'h10 ;
			data[67748] <= 8'h10 ;
			data[67749] <= 8'h10 ;
			data[67750] <= 8'h10 ;
			data[67751] <= 8'h10 ;
			data[67752] <= 8'h10 ;
			data[67753] <= 8'h10 ;
			data[67754] <= 8'h10 ;
			data[67755] <= 8'h10 ;
			data[67756] <= 8'h10 ;
			data[67757] <= 8'h10 ;
			data[67758] <= 8'h10 ;
			data[67759] <= 8'h10 ;
			data[67760] <= 8'h10 ;
			data[67761] <= 8'h10 ;
			data[67762] <= 8'h10 ;
			data[67763] <= 8'h10 ;
			data[67764] <= 8'h10 ;
			data[67765] <= 8'h10 ;
			data[67766] <= 8'h10 ;
			data[67767] <= 8'h10 ;
			data[67768] <= 8'h10 ;
			data[67769] <= 8'h10 ;
			data[67770] <= 8'h10 ;
			data[67771] <= 8'h10 ;
			data[67772] <= 8'h10 ;
			data[67773] <= 8'h10 ;
			data[67774] <= 8'h10 ;
			data[67775] <= 8'h10 ;
			data[67776] <= 8'h10 ;
			data[67777] <= 8'h10 ;
			data[67778] <= 8'h10 ;
			data[67779] <= 8'h10 ;
			data[67780] <= 8'h10 ;
			data[67781] <= 8'h10 ;
			data[67782] <= 8'h10 ;
			data[67783] <= 8'h10 ;
			data[67784] <= 8'h10 ;
			data[67785] <= 8'h10 ;
			data[67786] <= 8'h10 ;
			data[67787] <= 8'h10 ;
			data[67788] <= 8'h10 ;
			data[67789] <= 8'h10 ;
			data[67790] <= 8'h10 ;
			data[67791] <= 8'h10 ;
			data[67792] <= 8'h10 ;
			data[67793] <= 8'h10 ;
			data[67794] <= 8'h10 ;
			data[67795] <= 8'h10 ;
			data[67796] <= 8'h10 ;
			data[67797] <= 8'h10 ;
			data[67798] <= 8'h10 ;
			data[67799] <= 8'h10 ;
			data[67800] <= 8'h10 ;
			data[67801] <= 8'h10 ;
			data[67802] <= 8'h10 ;
			data[67803] <= 8'h10 ;
			data[67804] <= 8'h10 ;
			data[67805] <= 8'h10 ;
			data[67806] <= 8'h10 ;
			data[67807] <= 8'h10 ;
			data[67808] <= 8'h10 ;
			data[67809] <= 8'h10 ;
			data[67810] <= 8'h10 ;
			data[67811] <= 8'h10 ;
			data[67812] <= 8'h10 ;
			data[67813] <= 8'h10 ;
			data[67814] <= 8'h10 ;
			data[67815] <= 8'h10 ;
			data[67816] <= 8'h10 ;
			data[67817] <= 8'h10 ;
			data[67818] <= 8'h10 ;
			data[67819] <= 8'h10 ;
			data[67820] <= 8'h10 ;
			data[67821] <= 8'h10 ;
			data[67822] <= 8'h10 ;
			data[67823] <= 8'h10 ;
			data[67824] <= 8'h10 ;
			data[67825] <= 8'h10 ;
			data[67826] <= 8'h10 ;
			data[67827] <= 8'h10 ;
			data[67828] <= 8'h10 ;
			data[67829] <= 8'h10 ;
			data[67830] <= 8'h10 ;
			data[67831] <= 8'h10 ;
			data[67832] <= 8'h10 ;
			data[67833] <= 8'h10 ;
			data[67834] <= 8'h10 ;
			data[67835] <= 8'h10 ;
			data[67836] <= 8'h10 ;
			data[67837] <= 8'h10 ;
			data[67838] <= 8'h10 ;
			data[67839] <= 8'h10 ;
			data[67840] <= 8'h10 ;
			data[67841] <= 8'h10 ;
			data[67842] <= 8'h10 ;
			data[67843] <= 8'h10 ;
			data[67844] <= 8'h10 ;
			data[67845] <= 8'h10 ;
			data[67846] <= 8'h10 ;
			data[67847] <= 8'h10 ;
			data[67848] <= 8'h10 ;
			data[67849] <= 8'h10 ;
			data[67850] <= 8'h10 ;
			data[67851] <= 8'h10 ;
			data[67852] <= 8'h10 ;
			data[67853] <= 8'h10 ;
			data[67854] <= 8'h10 ;
			data[67855] <= 8'h10 ;
			data[67856] <= 8'h10 ;
			data[67857] <= 8'h10 ;
			data[67858] <= 8'h10 ;
			data[67859] <= 8'h10 ;
			data[67860] <= 8'h10 ;
			data[67861] <= 8'h10 ;
			data[67862] <= 8'h10 ;
			data[67863] <= 8'h10 ;
			data[67864] <= 8'h10 ;
			data[67865] <= 8'h10 ;
			data[67866] <= 8'h10 ;
			data[67867] <= 8'h10 ;
			data[67868] <= 8'h10 ;
			data[67869] <= 8'h10 ;
			data[67870] <= 8'h10 ;
			data[67871] <= 8'h10 ;
			data[67872] <= 8'h10 ;
			data[67873] <= 8'h10 ;
			data[67874] <= 8'h10 ;
			data[67875] <= 8'h10 ;
			data[67876] <= 8'h10 ;
			data[67877] <= 8'h10 ;
			data[67878] <= 8'h10 ;
			data[67879] <= 8'h10 ;
			data[67880] <= 8'h10 ;
			data[67881] <= 8'h10 ;
			data[67882] <= 8'h10 ;
			data[67883] <= 8'h10 ;
			data[67884] <= 8'h10 ;
			data[67885] <= 8'h10 ;
			data[67886] <= 8'h10 ;
			data[67887] <= 8'h10 ;
			data[67888] <= 8'h10 ;
			data[67889] <= 8'h10 ;
			data[67890] <= 8'h10 ;
			data[67891] <= 8'h10 ;
			data[67892] <= 8'h10 ;
			data[67893] <= 8'h10 ;
			data[67894] <= 8'h10 ;
			data[67895] <= 8'h10 ;
			data[67896] <= 8'h10 ;
			data[67897] <= 8'h10 ;
			data[67898] <= 8'h10 ;
			data[67899] <= 8'h10 ;
			data[67900] <= 8'h10 ;
			data[67901] <= 8'h10 ;
			data[67902] <= 8'h10 ;
			data[67903] <= 8'h10 ;
			data[67904] <= 8'h10 ;
			data[67905] <= 8'h10 ;
			data[67906] <= 8'h10 ;
			data[67907] <= 8'h10 ;
			data[67908] <= 8'h10 ;
			data[67909] <= 8'h10 ;
			data[67910] <= 8'h10 ;
			data[67911] <= 8'h10 ;
			data[67912] <= 8'h10 ;
			data[67913] <= 8'h10 ;
			data[67914] <= 8'h10 ;
			data[67915] <= 8'h10 ;
			data[67916] <= 8'h10 ;
			data[67917] <= 8'h10 ;
			data[67918] <= 8'h10 ;
			data[67919] <= 8'h10 ;
			data[67920] <= 8'h10 ;
			data[67921] <= 8'h10 ;
			data[67922] <= 8'h10 ;
			data[67923] <= 8'h10 ;
			data[67924] <= 8'h10 ;
			data[67925] <= 8'h10 ;
			data[67926] <= 8'h10 ;
			data[67927] <= 8'h10 ;
			data[67928] <= 8'h10 ;
			data[67929] <= 8'h10 ;
			data[67930] <= 8'h10 ;
			data[67931] <= 8'h10 ;
			data[67932] <= 8'h10 ;
			data[67933] <= 8'h10 ;
			data[67934] <= 8'h10 ;
			data[67935] <= 8'h10 ;
			data[67936] <= 8'h10 ;
			data[67937] <= 8'h10 ;
			data[67938] <= 8'h10 ;
			data[67939] <= 8'h10 ;
			data[67940] <= 8'h10 ;
			data[67941] <= 8'h10 ;
			data[67942] <= 8'h10 ;
			data[67943] <= 8'h10 ;
			data[67944] <= 8'h10 ;
			data[67945] <= 8'h10 ;
			data[67946] <= 8'h10 ;
			data[67947] <= 8'h10 ;
			data[67948] <= 8'h10 ;
			data[67949] <= 8'h10 ;
			data[67950] <= 8'h10 ;
			data[67951] <= 8'h10 ;
			data[67952] <= 8'h10 ;
			data[67953] <= 8'h10 ;
			data[67954] <= 8'h10 ;
			data[67955] <= 8'h10 ;
			data[67956] <= 8'h10 ;
			data[67957] <= 8'h10 ;
			data[67958] <= 8'h10 ;
			data[67959] <= 8'h10 ;
			data[67960] <= 8'h10 ;
			data[67961] <= 8'h10 ;
			data[67962] <= 8'h10 ;
			data[67963] <= 8'h10 ;
			data[67964] <= 8'h10 ;
			data[67965] <= 8'h10 ;
			data[67966] <= 8'h10 ;
			data[67967] <= 8'h10 ;
			data[67968] <= 8'h10 ;
			data[67969] <= 8'h10 ;
			data[67970] <= 8'h10 ;
			data[67971] <= 8'h10 ;
			data[67972] <= 8'h10 ;
			data[67973] <= 8'h10 ;
			data[67974] <= 8'h10 ;
			data[67975] <= 8'h10 ;
			data[67976] <= 8'h10 ;
			data[67977] <= 8'h10 ;
			data[67978] <= 8'h10 ;
			data[67979] <= 8'h10 ;
			data[67980] <= 8'h10 ;
			data[67981] <= 8'h10 ;
			data[67982] <= 8'h10 ;
			data[67983] <= 8'h10 ;
			data[67984] <= 8'h10 ;
			data[67985] <= 8'h10 ;
			data[67986] <= 8'h10 ;
			data[67987] <= 8'h10 ;
			data[67988] <= 8'h10 ;
			data[67989] <= 8'h10 ;
			data[67990] <= 8'h10 ;
			data[67991] <= 8'h10 ;
			data[67992] <= 8'h10 ;
			data[67993] <= 8'h10 ;
			data[67994] <= 8'h10 ;
			data[67995] <= 8'h10 ;
			data[67996] <= 8'h10 ;
			data[67997] <= 8'h10 ;
			data[67998] <= 8'h10 ;
			data[67999] <= 8'h10 ;
			data[68000] <= 8'h10 ;
			data[68001] <= 8'h10 ;
			data[68002] <= 8'h10 ;
			data[68003] <= 8'h10 ;
			data[68004] <= 8'h10 ;
			data[68005] <= 8'h10 ;
			data[68006] <= 8'h10 ;
			data[68007] <= 8'h10 ;
			data[68008] <= 8'h10 ;
			data[68009] <= 8'h10 ;
			data[68010] <= 8'h10 ;
			data[68011] <= 8'h10 ;
			data[68012] <= 8'h10 ;
			data[68013] <= 8'h10 ;
			data[68014] <= 8'h10 ;
			data[68015] <= 8'h10 ;
			data[68016] <= 8'h10 ;
			data[68017] <= 8'h10 ;
			data[68018] <= 8'h10 ;
			data[68019] <= 8'h10 ;
			data[68020] <= 8'h10 ;
			data[68021] <= 8'h10 ;
			data[68022] <= 8'h10 ;
			data[68023] <= 8'h10 ;
			data[68024] <= 8'h10 ;
			data[68025] <= 8'h10 ;
			data[68026] <= 8'h10 ;
			data[68027] <= 8'h10 ;
			data[68028] <= 8'h10 ;
			data[68029] <= 8'h10 ;
			data[68030] <= 8'h10 ;
			data[68031] <= 8'h10 ;
			data[68032] <= 8'h10 ;
			data[68033] <= 8'h10 ;
			data[68034] <= 8'h10 ;
			data[68035] <= 8'h10 ;
			data[68036] <= 8'h10 ;
			data[68037] <= 8'h10 ;
			data[68038] <= 8'h10 ;
			data[68039] <= 8'h10 ;
			data[68040] <= 8'h10 ;
			data[68041] <= 8'h10 ;
			data[68042] <= 8'h10 ;
			data[68043] <= 8'h10 ;
			data[68044] <= 8'h10 ;
			data[68045] <= 8'h10 ;
			data[68046] <= 8'h10 ;
			data[68047] <= 8'h10 ;
			data[68048] <= 8'h10 ;
			data[68049] <= 8'h10 ;
			data[68050] <= 8'h10 ;
			data[68051] <= 8'h10 ;
			data[68052] <= 8'h10 ;
			data[68053] <= 8'h10 ;
			data[68054] <= 8'h10 ;
			data[68055] <= 8'h10 ;
			data[68056] <= 8'h10 ;
			data[68057] <= 8'h10 ;
			data[68058] <= 8'h10 ;
			data[68059] <= 8'h10 ;
			data[68060] <= 8'h10 ;
			data[68061] <= 8'h10 ;
			data[68062] <= 8'h10 ;
			data[68063] <= 8'h10 ;
			data[68064] <= 8'h10 ;
			data[68065] <= 8'h10 ;
			data[68066] <= 8'h10 ;
			data[68067] <= 8'h10 ;
			data[68068] <= 8'h10 ;
			data[68069] <= 8'h10 ;
			data[68070] <= 8'h10 ;
			data[68071] <= 8'h10 ;
			data[68072] <= 8'h10 ;
			data[68073] <= 8'h10 ;
			data[68074] <= 8'h10 ;
			data[68075] <= 8'h10 ;
			data[68076] <= 8'h10 ;
			data[68077] <= 8'h10 ;
			data[68078] <= 8'h10 ;
			data[68079] <= 8'h10 ;
			data[68080] <= 8'h10 ;
			data[68081] <= 8'h10 ;
			data[68082] <= 8'h10 ;
			data[68083] <= 8'h10 ;
			data[68084] <= 8'h10 ;
			data[68085] <= 8'h10 ;
			data[68086] <= 8'h10 ;
			data[68087] <= 8'h10 ;
			data[68088] <= 8'h10 ;
			data[68089] <= 8'h10 ;
			data[68090] <= 8'h10 ;
			data[68091] <= 8'h10 ;
			data[68092] <= 8'h10 ;
			data[68093] <= 8'h10 ;
			data[68094] <= 8'h10 ;
			data[68095] <= 8'h10 ;
			data[68096] <= 8'h10 ;
			data[68097] <= 8'h10 ;
			data[68098] <= 8'h10 ;
			data[68099] <= 8'h10 ;
			data[68100] <= 8'h10 ;
			data[68101] <= 8'h10 ;
			data[68102] <= 8'h10 ;
			data[68103] <= 8'h10 ;
			data[68104] <= 8'h10 ;
			data[68105] <= 8'h10 ;
			data[68106] <= 8'h10 ;
			data[68107] <= 8'h10 ;
			data[68108] <= 8'h10 ;
			data[68109] <= 8'h10 ;
			data[68110] <= 8'h10 ;
			data[68111] <= 8'h10 ;
			data[68112] <= 8'h10 ;
			data[68113] <= 8'h10 ;
			data[68114] <= 8'h10 ;
			data[68115] <= 8'h10 ;
			data[68116] <= 8'h10 ;
			data[68117] <= 8'h10 ;
			data[68118] <= 8'h10 ;
			data[68119] <= 8'h10 ;
			data[68120] <= 8'h10 ;
			data[68121] <= 8'h10 ;
			data[68122] <= 8'h10 ;
			data[68123] <= 8'h10 ;
			data[68124] <= 8'h10 ;
			data[68125] <= 8'h10 ;
			data[68126] <= 8'h10 ;
			data[68127] <= 8'h10 ;
			data[68128] <= 8'h10 ;
			data[68129] <= 8'h10 ;
			data[68130] <= 8'h10 ;
			data[68131] <= 8'h10 ;
			data[68132] <= 8'h10 ;
			data[68133] <= 8'h10 ;
			data[68134] <= 8'h10 ;
			data[68135] <= 8'h10 ;
			data[68136] <= 8'h10 ;
			data[68137] <= 8'h10 ;
			data[68138] <= 8'h10 ;
			data[68139] <= 8'h10 ;
			data[68140] <= 8'h10 ;
			data[68141] <= 8'h10 ;
			data[68142] <= 8'h10 ;
			data[68143] <= 8'h10 ;
			data[68144] <= 8'h10 ;
			data[68145] <= 8'h10 ;
			data[68146] <= 8'h10 ;
			data[68147] <= 8'h10 ;
			data[68148] <= 8'h10 ;
			data[68149] <= 8'h10 ;
			data[68150] <= 8'h10 ;
			data[68151] <= 8'h10 ;
			data[68152] <= 8'h10 ;
			data[68153] <= 8'h10 ;
			data[68154] <= 8'h10 ;
			data[68155] <= 8'h10 ;
			data[68156] <= 8'h10 ;
			data[68157] <= 8'h10 ;
			data[68158] <= 8'h10 ;
			data[68159] <= 8'h10 ;
			data[68160] <= 8'h10 ;
			data[68161] <= 8'h10 ;
			data[68162] <= 8'h10 ;
			data[68163] <= 8'h10 ;
			data[68164] <= 8'h10 ;
			data[68165] <= 8'h10 ;
			data[68166] <= 8'h10 ;
			data[68167] <= 8'h10 ;
			data[68168] <= 8'h10 ;
			data[68169] <= 8'h10 ;
			data[68170] <= 8'h10 ;
			data[68171] <= 8'h10 ;
			data[68172] <= 8'h10 ;
			data[68173] <= 8'h10 ;
			data[68174] <= 8'h10 ;
			data[68175] <= 8'h10 ;
			data[68176] <= 8'h10 ;
			data[68177] <= 8'h10 ;
			data[68178] <= 8'h10 ;
			data[68179] <= 8'h10 ;
			data[68180] <= 8'h10 ;
			data[68181] <= 8'h10 ;
			data[68182] <= 8'h10 ;
			data[68183] <= 8'h10 ;
			data[68184] <= 8'h10 ;
			data[68185] <= 8'h10 ;
			data[68186] <= 8'h10 ;
			data[68187] <= 8'h10 ;
			data[68188] <= 8'h10 ;
			data[68189] <= 8'h10 ;
			data[68190] <= 8'h10 ;
			data[68191] <= 8'h10 ;
			data[68192] <= 8'h10 ;
			data[68193] <= 8'h10 ;
			data[68194] <= 8'h10 ;
			data[68195] <= 8'h10 ;
			data[68196] <= 8'h10 ;
			data[68197] <= 8'h10 ;
			data[68198] <= 8'h10 ;
			data[68199] <= 8'h10 ;
			data[68200] <= 8'h10 ;
			data[68201] <= 8'h10 ;
			data[68202] <= 8'h10 ;
			data[68203] <= 8'h10 ;
			data[68204] <= 8'h10 ;
			data[68205] <= 8'h10 ;
			data[68206] <= 8'h10 ;
			data[68207] <= 8'h10 ;
			data[68208] <= 8'h10 ;
			data[68209] <= 8'h10 ;
			data[68210] <= 8'h10 ;
			data[68211] <= 8'h10 ;
			data[68212] <= 8'h10 ;
			data[68213] <= 8'h10 ;
			data[68214] <= 8'h10 ;
			data[68215] <= 8'h10 ;
			data[68216] <= 8'h10 ;
			data[68217] <= 8'h10 ;
			data[68218] <= 8'h10 ;
			data[68219] <= 8'h10 ;
			data[68220] <= 8'h10 ;
			data[68221] <= 8'h10 ;
			data[68222] <= 8'h10 ;
			data[68223] <= 8'h10 ;
			data[68224] <= 8'h10 ;
			data[68225] <= 8'h10 ;
			data[68226] <= 8'h10 ;
			data[68227] <= 8'h10 ;
			data[68228] <= 8'h10 ;
			data[68229] <= 8'h10 ;
			data[68230] <= 8'h10 ;
			data[68231] <= 8'h10 ;
			data[68232] <= 8'h10 ;
			data[68233] <= 8'h10 ;
			data[68234] <= 8'h10 ;
			data[68235] <= 8'h10 ;
			data[68236] <= 8'h10 ;
			data[68237] <= 8'h10 ;
			data[68238] <= 8'h10 ;
			data[68239] <= 8'h10 ;
			data[68240] <= 8'h10 ;
			data[68241] <= 8'h10 ;
			data[68242] <= 8'h10 ;
			data[68243] <= 8'h10 ;
			data[68244] <= 8'h10 ;
			data[68245] <= 8'h10 ;
			data[68246] <= 8'h10 ;
			data[68247] <= 8'h10 ;
			data[68248] <= 8'h10 ;
			data[68249] <= 8'h10 ;
			data[68250] <= 8'h10 ;
			data[68251] <= 8'h10 ;
			data[68252] <= 8'h10 ;
			data[68253] <= 8'h10 ;
			data[68254] <= 8'h10 ;
			data[68255] <= 8'h10 ;
			data[68256] <= 8'h10 ;
			data[68257] <= 8'h10 ;
			data[68258] <= 8'h10 ;
			data[68259] <= 8'h10 ;
			data[68260] <= 8'h10 ;
			data[68261] <= 8'h10 ;
			data[68262] <= 8'h10 ;
			data[68263] <= 8'h10 ;
			data[68264] <= 8'h10 ;
			data[68265] <= 8'h10 ;
			data[68266] <= 8'h10 ;
			data[68267] <= 8'h10 ;
			data[68268] <= 8'h10 ;
			data[68269] <= 8'h10 ;
			data[68270] <= 8'h10 ;
			data[68271] <= 8'h10 ;
			data[68272] <= 8'h10 ;
			data[68273] <= 8'h10 ;
			data[68274] <= 8'h10 ;
			data[68275] <= 8'h10 ;
			data[68276] <= 8'h10 ;
			data[68277] <= 8'h10 ;
			data[68278] <= 8'h10 ;
			data[68279] <= 8'h10 ;
			data[68280] <= 8'h10 ;
			data[68281] <= 8'h10 ;
			data[68282] <= 8'h10 ;
			data[68283] <= 8'h10 ;
			data[68284] <= 8'h10 ;
			data[68285] <= 8'h10 ;
			data[68286] <= 8'h10 ;
			data[68287] <= 8'h10 ;
			data[68288] <= 8'h10 ;
			data[68289] <= 8'h10 ;
			data[68290] <= 8'h10 ;
			data[68291] <= 8'h10 ;
			data[68292] <= 8'h10 ;
			data[68293] <= 8'h10 ;
			data[68294] <= 8'h10 ;
			data[68295] <= 8'h10 ;
			data[68296] <= 8'h10 ;
			data[68297] <= 8'h10 ;
			data[68298] <= 8'h10 ;
			data[68299] <= 8'h10 ;
			data[68300] <= 8'h10 ;
			data[68301] <= 8'h10 ;
			data[68302] <= 8'h10 ;
			data[68303] <= 8'h10 ;
			data[68304] <= 8'h10 ;
			data[68305] <= 8'h10 ;
			data[68306] <= 8'h10 ;
			data[68307] <= 8'h10 ;
			data[68308] <= 8'h10 ;
			data[68309] <= 8'h10 ;
			data[68310] <= 8'h10 ;
			data[68311] <= 8'h10 ;
			data[68312] <= 8'h10 ;
			data[68313] <= 8'h10 ;
			data[68314] <= 8'h10 ;
			data[68315] <= 8'h10 ;
			data[68316] <= 8'h10 ;
			data[68317] <= 8'h10 ;
			data[68318] <= 8'h10 ;
			data[68319] <= 8'h10 ;
			data[68320] <= 8'h10 ;
			data[68321] <= 8'h10 ;
			data[68322] <= 8'h10 ;
			data[68323] <= 8'h10 ;
			data[68324] <= 8'h10 ;
			data[68325] <= 8'h10 ;
			data[68326] <= 8'h10 ;
			data[68327] <= 8'h10 ;
			data[68328] <= 8'h10 ;
			data[68329] <= 8'h10 ;
			data[68330] <= 8'h10 ;
			data[68331] <= 8'h10 ;
			data[68332] <= 8'h10 ;
			data[68333] <= 8'h10 ;
			data[68334] <= 8'h10 ;
			data[68335] <= 8'h10 ;
			data[68336] <= 8'h10 ;
			data[68337] <= 8'h10 ;
			data[68338] <= 8'h10 ;
			data[68339] <= 8'h10 ;
			data[68340] <= 8'h10 ;
			data[68341] <= 8'h10 ;
			data[68342] <= 8'h10 ;
			data[68343] <= 8'h10 ;
			data[68344] <= 8'h10 ;
			data[68345] <= 8'h10 ;
			data[68346] <= 8'h10 ;
			data[68347] <= 8'h10 ;
			data[68348] <= 8'h10 ;
			data[68349] <= 8'h10 ;
			data[68350] <= 8'h10 ;
			data[68351] <= 8'h10 ;
			data[68352] <= 8'h10 ;
			data[68353] <= 8'h10 ;
			data[68354] <= 8'h10 ;
			data[68355] <= 8'h10 ;
			data[68356] <= 8'h10 ;
			data[68357] <= 8'h10 ;
			data[68358] <= 8'h10 ;
			data[68359] <= 8'h10 ;
			data[68360] <= 8'h10 ;
			data[68361] <= 8'h10 ;
			data[68362] <= 8'h10 ;
			data[68363] <= 8'h10 ;
			data[68364] <= 8'h10 ;
			data[68365] <= 8'h10 ;
			data[68366] <= 8'h10 ;
			data[68367] <= 8'h10 ;
			data[68368] <= 8'h10 ;
			data[68369] <= 8'h10 ;
			data[68370] <= 8'h10 ;
			data[68371] <= 8'h10 ;
			data[68372] <= 8'h10 ;
			data[68373] <= 8'h10 ;
			data[68374] <= 8'h10 ;
			data[68375] <= 8'h10 ;
			data[68376] <= 8'h10 ;
			data[68377] <= 8'h10 ;
			data[68378] <= 8'h10 ;
			data[68379] <= 8'h10 ;
			data[68380] <= 8'h10 ;
			data[68381] <= 8'h10 ;
			data[68382] <= 8'h10 ;
			data[68383] <= 8'h10 ;
			data[68384] <= 8'h10 ;
			data[68385] <= 8'h10 ;
			data[68386] <= 8'h10 ;
			data[68387] <= 8'h10 ;
			data[68388] <= 8'h10 ;
			data[68389] <= 8'h10 ;
			data[68390] <= 8'h10 ;
			data[68391] <= 8'h10 ;
			data[68392] <= 8'h10 ;
			data[68393] <= 8'h10 ;
			data[68394] <= 8'h10 ;
			data[68395] <= 8'h10 ;
			data[68396] <= 8'h10 ;
			data[68397] <= 8'h10 ;
			data[68398] <= 8'h10 ;
			data[68399] <= 8'h10 ;
			data[68400] <= 8'h10 ;
			data[68401] <= 8'h10 ;
			data[68402] <= 8'h10 ;
			data[68403] <= 8'h10 ;
			data[68404] <= 8'h10 ;
			data[68405] <= 8'h10 ;
			data[68406] <= 8'h10 ;
			data[68407] <= 8'h10 ;
			data[68408] <= 8'h10 ;
			data[68409] <= 8'h10 ;
			data[68410] <= 8'h10 ;
			data[68411] <= 8'h10 ;
			data[68412] <= 8'h10 ;
			data[68413] <= 8'h10 ;
			data[68414] <= 8'h10 ;
			data[68415] <= 8'h10 ;
			data[68416] <= 8'h10 ;
			data[68417] <= 8'h10 ;
			data[68418] <= 8'h10 ;
			data[68419] <= 8'h10 ;
			data[68420] <= 8'h10 ;
			data[68421] <= 8'h10 ;
			data[68422] <= 8'h10 ;
			data[68423] <= 8'h10 ;
			data[68424] <= 8'h10 ;
			data[68425] <= 8'h10 ;
			data[68426] <= 8'h10 ;
			data[68427] <= 8'h10 ;
			data[68428] <= 8'h10 ;
			data[68429] <= 8'h10 ;
			data[68430] <= 8'h10 ;
			data[68431] <= 8'h10 ;
			data[68432] <= 8'h10 ;
			data[68433] <= 8'h10 ;
			data[68434] <= 8'h10 ;
			data[68435] <= 8'h10 ;
			data[68436] <= 8'h10 ;
			data[68437] <= 8'h10 ;
			data[68438] <= 8'h10 ;
			data[68439] <= 8'h10 ;
			data[68440] <= 8'h10 ;
			data[68441] <= 8'h10 ;
			data[68442] <= 8'h10 ;
			data[68443] <= 8'h10 ;
			data[68444] <= 8'h10 ;
			data[68445] <= 8'h10 ;
			data[68446] <= 8'h10 ;
			data[68447] <= 8'h10 ;
			data[68448] <= 8'h10 ;
			data[68449] <= 8'h10 ;
			data[68450] <= 8'h10 ;
			data[68451] <= 8'h10 ;
			data[68452] <= 8'h10 ;
			data[68453] <= 8'h10 ;
			data[68454] <= 8'h10 ;
			data[68455] <= 8'h10 ;
			data[68456] <= 8'h10 ;
			data[68457] <= 8'h10 ;
			data[68458] <= 8'h10 ;
			data[68459] <= 8'h10 ;
			data[68460] <= 8'h10 ;
			data[68461] <= 8'h10 ;
			data[68462] <= 8'h10 ;
			data[68463] <= 8'h10 ;
			data[68464] <= 8'h10 ;
			data[68465] <= 8'h10 ;
			data[68466] <= 8'h10 ;
			data[68467] <= 8'h10 ;
			data[68468] <= 8'h10 ;
			data[68469] <= 8'h10 ;
			data[68470] <= 8'h10 ;
			data[68471] <= 8'h10 ;
			data[68472] <= 8'h10 ;
			data[68473] <= 8'h10 ;
			data[68474] <= 8'h10 ;
			data[68475] <= 8'h10 ;
			data[68476] <= 8'h10 ;
			data[68477] <= 8'h10 ;
			data[68478] <= 8'h10 ;
			data[68479] <= 8'h10 ;
			data[68480] <= 8'h10 ;
			data[68481] <= 8'h10 ;
			data[68482] <= 8'h10 ;
			data[68483] <= 8'h10 ;
			data[68484] <= 8'h10 ;
			data[68485] <= 8'h10 ;
			data[68486] <= 8'h10 ;
			data[68487] <= 8'h10 ;
			data[68488] <= 8'h10 ;
			data[68489] <= 8'h10 ;
			data[68490] <= 8'h10 ;
			data[68491] <= 8'h10 ;
			data[68492] <= 8'h10 ;
			data[68493] <= 8'h10 ;
			data[68494] <= 8'h10 ;
			data[68495] <= 8'h10 ;
			data[68496] <= 8'h10 ;
			data[68497] <= 8'h10 ;
			data[68498] <= 8'h10 ;
			data[68499] <= 8'h10 ;
			data[68500] <= 8'h10 ;
			data[68501] <= 8'h10 ;
			data[68502] <= 8'h10 ;
			data[68503] <= 8'h10 ;
			data[68504] <= 8'h10 ;
			data[68505] <= 8'h10 ;
			data[68506] <= 8'h10 ;
			data[68507] <= 8'h10 ;
			data[68508] <= 8'h10 ;
			data[68509] <= 8'h10 ;
			data[68510] <= 8'h10 ;
			data[68511] <= 8'h10 ;
			data[68512] <= 8'h10 ;
			data[68513] <= 8'h10 ;
			data[68514] <= 8'h10 ;
			data[68515] <= 8'h10 ;
			data[68516] <= 8'h10 ;
			data[68517] <= 8'h10 ;
			data[68518] <= 8'h10 ;
			data[68519] <= 8'h10 ;
			data[68520] <= 8'h10 ;
			data[68521] <= 8'h10 ;
			data[68522] <= 8'h10 ;
			data[68523] <= 8'h10 ;
			data[68524] <= 8'h10 ;
			data[68525] <= 8'h10 ;
			data[68526] <= 8'h10 ;
			data[68527] <= 8'h10 ;
			data[68528] <= 8'h10 ;
			data[68529] <= 8'h10 ;
			data[68530] <= 8'h10 ;
			data[68531] <= 8'h10 ;
			data[68532] <= 8'h10 ;
			data[68533] <= 8'h10 ;
			data[68534] <= 8'h10 ;
			data[68535] <= 8'h10 ;
			data[68536] <= 8'h10 ;
			data[68537] <= 8'h10 ;
			data[68538] <= 8'h10 ;
			data[68539] <= 8'h10 ;
			data[68540] <= 8'h10 ;
			data[68541] <= 8'h10 ;
			data[68542] <= 8'h10 ;
			data[68543] <= 8'h10 ;
			data[68544] <= 8'h10 ;
			data[68545] <= 8'h10 ;
			data[68546] <= 8'h10 ;
			data[68547] <= 8'h10 ;
			data[68548] <= 8'h10 ;
			data[68549] <= 8'h10 ;
			data[68550] <= 8'h10 ;
			data[68551] <= 8'h10 ;
			data[68552] <= 8'h10 ;
			data[68553] <= 8'h10 ;
			data[68554] <= 8'h10 ;
			data[68555] <= 8'h10 ;
			data[68556] <= 8'h10 ;
			data[68557] <= 8'h10 ;
			data[68558] <= 8'h10 ;
			data[68559] <= 8'h10 ;
			data[68560] <= 8'h10 ;
			data[68561] <= 8'h10 ;
			data[68562] <= 8'h10 ;
			data[68563] <= 8'h10 ;
			data[68564] <= 8'h10 ;
			data[68565] <= 8'h10 ;
			data[68566] <= 8'h10 ;
			data[68567] <= 8'h10 ;
			data[68568] <= 8'h10 ;
			data[68569] <= 8'h10 ;
			data[68570] <= 8'h10 ;
			data[68571] <= 8'h10 ;
			data[68572] <= 8'h10 ;
			data[68573] <= 8'h10 ;
			data[68574] <= 8'h10 ;
			data[68575] <= 8'h10 ;
			data[68576] <= 8'h10 ;
			data[68577] <= 8'h10 ;
			data[68578] <= 8'h10 ;
			data[68579] <= 8'h10 ;
			data[68580] <= 8'h10 ;
			data[68581] <= 8'h10 ;
			data[68582] <= 8'h10 ;
			data[68583] <= 8'h10 ;
			data[68584] <= 8'h10 ;
			data[68585] <= 8'h10 ;
			data[68586] <= 8'h10 ;
			data[68587] <= 8'h10 ;
			data[68588] <= 8'h10 ;
			data[68589] <= 8'h10 ;
			data[68590] <= 8'h10 ;
			data[68591] <= 8'h10 ;
			data[68592] <= 8'h10 ;
			data[68593] <= 8'h10 ;
			data[68594] <= 8'h10 ;
			data[68595] <= 8'h10 ;
			data[68596] <= 8'h10 ;
			data[68597] <= 8'h10 ;
			data[68598] <= 8'h10 ;
			data[68599] <= 8'h10 ;
			data[68600] <= 8'h10 ;
			data[68601] <= 8'h10 ;
			data[68602] <= 8'h10 ;
			data[68603] <= 8'h10 ;
			data[68604] <= 8'h10 ;
			data[68605] <= 8'h10 ;
			data[68606] <= 8'h10 ;
			data[68607] <= 8'h10 ;
			data[68608] <= 8'h10 ;
			data[68609] <= 8'h10 ;
			data[68610] <= 8'h10 ;
			data[68611] <= 8'h10 ;
			data[68612] <= 8'h10 ;
			data[68613] <= 8'h10 ;
			data[68614] <= 8'h10 ;
			data[68615] <= 8'h10 ;
			data[68616] <= 8'h10 ;
			data[68617] <= 8'h10 ;
			data[68618] <= 8'h10 ;
			data[68619] <= 8'h10 ;
			data[68620] <= 8'h10 ;
			data[68621] <= 8'h10 ;
			data[68622] <= 8'h10 ;
			data[68623] <= 8'h10 ;
			data[68624] <= 8'h10 ;
			data[68625] <= 8'h10 ;
			data[68626] <= 8'h10 ;
			data[68627] <= 8'h10 ;
			data[68628] <= 8'h10 ;
			data[68629] <= 8'h10 ;
			data[68630] <= 8'h10 ;
			data[68631] <= 8'h10 ;
			data[68632] <= 8'h10 ;
			data[68633] <= 8'h10 ;
			data[68634] <= 8'h10 ;
			data[68635] <= 8'h10 ;
			data[68636] <= 8'h10 ;
			data[68637] <= 8'h10 ;
			data[68638] <= 8'h10 ;
			data[68639] <= 8'h10 ;
			data[68640] <= 8'h10 ;
			data[68641] <= 8'h10 ;
			data[68642] <= 8'h10 ;
			data[68643] <= 8'h10 ;
			data[68644] <= 8'h10 ;
			data[68645] <= 8'h10 ;
			data[68646] <= 8'h10 ;
			data[68647] <= 8'h10 ;
			data[68648] <= 8'h10 ;
			data[68649] <= 8'h10 ;
			data[68650] <= 8'h10 ;
			data[68651] <= 8'h10 ;
			data[68652] <= 8'h10 ;
			data[68653] <= 8'h10 ;
			data[68654] <= 8'h10 ;
			data[68655] <= 8'h10 ;
			data[68656] <= 8'h10 ;
			data[68657] <= 8'h10 ;
			data[68658] <= 8'h10 ;
			data[68659] <= 8'h10 ;
			data[68660] <= 8'h10 ;
			data[68661] <= 8'h10 ;
			data[68662] <= 8'h10 ;
			data[68663] <= 8'h10 ;
			data[68664] <= 8'h10 ;
			data[68665] <= 8'h10 ;
			data[68666] <= 8'h10 ;
			data[68667] <= 8'h10 ;
			data[68668] <= 8'h10 ;
			data[68669] <= 8'h10 ;
			data[68670] <= 8'h10 ;
			data[68671] <= 8'h10 ;
			data[68672] <= 8'h10 ;
			data[68673] <= 8'h10 ;
			data[68674] <= 8'h10 ;
			data[68675] <= 8'h10 ;
			data[68676] <= 8'h10 ;
			data[68677] <= 8'h10 ;
			data[68678] <= 8'h10 ;
			data[68679] <= 8'h10 ;
			data[68680] <= 8'h10 ;
			data[68681] <= 8'h10 ;
			data[68682] <= 8'h10 ;
			data[68683] <= 8'h10 ;
			data[68684] <= 8'h10 ;
			data[68685] <= 8'h10 ;
			data[68686] <= 8'h10 ;
			data[68687] <= 8'h10 ;
			data[68688] <= 8'h10 ;
			data[68689] <= 8'h10 ;
			data[68690] <= 8'h10 ;
			data[68691] <= 8'h10 ;
			data[68692] <= 8'h10 ;
			data[68693] <= 8'h10 ;
			data[68694] <= 8'h10 ;
			data[68695] <= 8'h10 ;
			data[68696] <= 8'h10 ;
			data[68697] <= 8'h10 ;
			data[68698] <= 8'h10 ;
			data[68699] <= 8'h10 ;
			data[68700] <= 8'h10 ;
			data[68701] <= 8'h10 ;
			data[68702] <= 8'h10 ;
			data[68703] <= 8'h10 ;
			data[68704] <= 8'h10 ;
			data[68705] <= 8'h10 ;
			data[68706] <= 8'h10 ;
			data[68707] <= 8'h10 ;
			data[68708] <= 8'h10 ;
			data[68709] <= 8'h10 ;
			data[68710] <= 8'h10 ;
			data[68711] <= 8'h10 ;
			data[68712] <= 8'h10 ;
			data[68713] <= 8'h10 ;
			data[68714] <= 8'h10 ;
			data[68715] <= 8'h10 ;
			data[68716] <= 8'h10 ;
			data[68717] <= 8'h10 ;
			data[68718] <= 8'h10 ;
			data[68719] <= 8'h10 ;
			data[68720] <= 8'h10 ;
			data[68721] <= 8'h10 ;
			data[68722] <= 8'h10 ;
			data[68723] <= 8'h10 ;
			data[68724] <= 8'h10 ;
			data[68725] <= 8'h10 ;
			data[68726] <= 8'h10 ;
			data[68727] <= 8'h10 ;
			data[68728] <= 8'h10 ;
			data[68729] <= 8'h10 ;
			data[68730] <= 8'h10 ;
			data[68731] <= 8'h10 ;
			data[68732] <= 8'h10 ;
			data[68733] <= 8'h10 ;
			data[68734] <= 8'h10 ;
			data[68735] <= 8'h10 ;
			data[68736] <= 8'h10 ;
			data[68737] <= 8'h10 ;
			data[68738] <= 8'h10 ;
			data[68739] <= 8'h10 ;
			data[68740] <= 8'h10 ;
			data[68741] <= 8'h10 ;
			data[68742] <= 8'h10 ;
			data[68743] <= 8'h10 ;
			data[68744] <= 8'h10 ;
			data[68745] <= 8'h10 ;
			data[68746] <= 8'h10 ;
			data[68747] <= 8'h10 ;
			data[68748] <= 8'h10 ;
			data[68749] <= 8'h10 ;
			data[68750] <= 8'h10 ;
			data[68751] <= 8'h10 ;
			data[68752] <= 8'h10 ;
			data[68753] <= 8'h10 ;
			data[68754] <= 8'h10 ;
			data[68755] <= 8'h10 ;
			data[68756] <= 8'h10 ;
			data[68757] <= 8'h10 ;
			data[68758] <= 8'h10 ;
			data[68759] <= 8'h10 ;
			data[68760] <= 8'h10 ;
			data[68761] <= 8'h10 ;
			data[68762] <= 8'h10 ;
			data[68763] <= 8'h10 ;
			data[68764] <= 8'h10 ;
			data[68765] <= 8'h10 ;
			data[68766] <= 8'h10 ;
			data[68767] <= 8'h10 ;
			data[68768] <= 8'h10 ;
			data[68769] <= 8'h10 ;
			data[68770] <= 8'h10 ;
			data[68771] <= 8'h10 ;
			data[68772] <= 8'h10 ;
			data[68773] <= 8'h10 ;
			data[68774] <= 8'h10 ;
			data[68775] <= 8'h10 ;
			data[68776] <= 8'h10 ;
			data[68777] <= 8'h10 ;
			data[68778] <= 8'h10 ;
			data[68779] <= 8'h10 ;
			data[68780] <= 8'h10 ;
			data[68781] <= 8'h10 ;
			data[68782] <= 8'h10 ;
			data[68783] <= 8'h10 ;
			data[68784] <= 8'h10 ;
			data[68785] <= 8'h10 ;
			data[68786] <= 8'h10 ;
			data[68787] <= 8'h10 ;
			data[68788] <= 8'h10 ;
			data[68789] <= 8'h10 ;
			data[68790] <= 8'h10 ;
			data[68791] <= 8'h10 ;
			data[68792] <= 8'h10 ;
			data[68793] <= 8'h10 ;
			data[68794] <= 8'h10 ;
			data[68795] <= 8'h10 ;
			data[68796] <= 8'h10 ;
			data[68797] <= 8'h10 ;
			data[68798] <= 8'h10 ;
			data[68799] <= 8'h10 ;
			data[68800] <= 8'h10 ;
			data[68801] <= 8'h10 ;
			data[68802] <= 8'h10 ;
			data[68803] <= 8'h10 ;
			data[68804] <= 8'h10 ;
			data[68805] <= 8'h10 ;
			data[68806] <= 8'h10 ;
			data[68807] <= 8'h10 ;
			data[68808] <= 8'h10 ;
			data[68809] <= 8'h10 ;
			data[68810] <= 8'h10 ;
			data[68811] <= 8'h10 ;
			data[68812] <= 8'h10 ;
			data[68813] <= 8'h10 ;
			data[68814] <= 8'h10 ;
			data[68815] <= 8'h10 ;
			data[68816] <= 8'h10 ;
			data[68817] <= 8'h10 ;
			data[68818] <= 8'h10 ;
			data[68819] <= 8'h10 ;
			data[68820] <= 8'h10 ;
			data[68821] <= 8'h10 ;
			data[68822] <= 8'h10 ;
			data[68823] <= 8'h10 ;
			data[68824] <= 8'h10 ;
			data[68825] <= 8'h10 ;
			data[68826] <= 8'h10 ;
			data[68827] <= 8'h10 ;
			data[68828] <= 8'h10 ;
			data[68829] <= 8'h10 ;
			data[68830] <= 8'h10 ;
			data[68831] <= 8'h10 ;
			data[68832] <= 8'h10 ;
			data[68833] <= 8'h10 ;
			data[68834] <= 8'h10 ;
			data[68835] <= 8'h10 ;
			data[68836] <= 8'h10 ;
			data[68837] <= 8'h10 ;
			data[68838] <= 8'h10 ;
			data[68839] <= 8'h10 ;
			data[68840] <= 8'h10 ;
			data[68841] <= 8'h10 ;
			data[68842] <= 8'h10 ;
			data[68843] <= 8'h10 ;
			data[68844] <= 8'h10 ;
			data[68845] <= 8'h10 ;
			data[68846] <= 8'h10 ;
			data[68847] <= 8'h10 ;
			data[68848] <= 8'h10 ;
			data[68849] <= 8'h10 ;
			data[68850] <= 8'h10 ;
			data[68851] <= 8'h10 ;
			data[68852] <= 8'h10 ;
			data[68853] <= 8'h10 ;
			data[68854] <= 8'h10 ;
			data[68855] <= 8'h10 ;
			data[68856] <= 8'h10 ;
			data[68857] <= 8'h10 ;
			data[68858] <= 8'h10 ;
			data[68859] <= 8'h10 ;
			data[68860] <= 8'h10 ;
			data[68861] <= 8'h10 ;
			data[68862] <= 8'h10 ;
			data[68863] <= 8'h10 ;
			data[68864] <= 8'h10 ;
			data[68865] <= 8'h10 ;
			data[68866] <= 8'h10 ;
			data[68867] <= 8'h10 ;
			data[68868] <= 8'h10 ;
			data[68869] <= 8'h10 ;
			data[68870] <= 8'h10 ;
			data[68871] <= 8'h10 ;
			data[68872] <= 8'h10 ;
			data[68873] <= 8'h10 ;
			data[68874] <= 8'h10 ;
			data[68875] <= 8'h10 ;
			data[68876] <= 8'h10 ;
			data[68877] <= 8'h10 ;
			data[68878] <= 8'h10 ;
			data[68879] <= 8'h10 ;
			data[68880] <= 8'h10 ;
			data[68881] <= 8'h10 ;
			data[68882] <= 8'h10 ;
			data[68883] <= 8'h10 ;
			data[68884] <= 8'h10 ;
			data[68885] <= 8'h10 ;
			data[68886] <= 8'h10 ;
			data[68887] <= 8'h10 ;
			data[68888] <= 8'h10 ;
			data[68889] <= 8'h10 ;
			data[68890] <= 8'h10 ;
			data[68891] <= 8'h10 ;
			data[68892] <= 8'h10 ;
			data[68893] <= 8'h10 ;
			data[68894] <= 8'h10 ;
			data[68895] <= 8'h10 ;
			data[68896] <= 8'h10 ;
			data[68897] <= 8'h10 ;
			data[68898] <= 8'h10 ;
			data[68899] <= 8'h10 ;
			data[68900] <= 8'h10 ;
			data[68901] <= 8'h10 ;
			data[68902] <= 8'h10 ;
			data[68903] <= 8'h10 ;
			data[68904] <= 8'h10 ;
			data[68905] <= 8'h10 ;
			data[68906] <= 8'h10 ;
			data[68907] <= 8'h10 ;
			data[68908] <= 8'h10 ;
			data[68909] <= 8'h10 ;
			data[68910] <= 8'h10 ;
			data[68911] <= 8'h10 ;
			data[68912] <= 8'h10 ;
			data[68913] <= 8'h10 ;
			data[68914] <= 8'h10 ;
			data[68915] <= 8'h10 ;
			data[68916] <= 8'h10 ;
			data[68917] <= 8'h10 ;
			data[68918] <= 8'h10 ;
			data[68919] <= 8'h10 ;
			data[68920] <= 8'h10 ;
			data[68921] <= 8'h10 ;
			data[68922] <= 8'h10 ;
			data[68923] <= 8'h10 ;
			data[68924] <= 8'h10 ;
			data[68925] <= 8'h10 ;
			data[68926] <= 8'h10 ;
			data[68927] <= 8'h10 ;
			data[68928] <= 8'h10 ;
			data[68929] <= 8'h10 ;
			data[68930] <= 8'h10 ;
			data[68931] <= 8'h10 ;
			data[68932] <= 8'h10 ;
			data[68933] <= 8'h10 ;
			data[68934] <= 8'h10 ;
			data[68935] <= 8'h10 ;
			data[68936] <= 8'h10 ;
			data[68937] <= 8'h10 ;
			data[68938] <= 8'h10 ;
			data[68939] <= 8'h10 ;
			data[68940] <= 8'h10 ;
			data[68941] <= 8'h10 ;
			data[68942] <= 8'h10 ;
			data[68943] <= 8'h10 ;
			data[68944] <= 8'h10 ;
			data[68945] <= 8'h10 ;
			data[68946] <= 8'h10 ;
			data[68947] <= 8'h10 ;
			data[68948] <= 8'h10 ;
			data[68949] <= 8'h10 ;
			data[68950] <= 8'h10 ;
			data[68951] <= 8'h10 ;
			data[68952] <= 8'h10 ;
			data[68953] <= 8'h10 ;
			data[68954] <= 8'h10 ;
			data[68955] <= 8'h10 ;
			data[68956] <= 8'h10 ;
			data[68957] <= 8'h10 ;
			data[68958] <= 8'h10 ;
			data[68959] <= 8'h10 ;
			data[68960] <= 8'h10 ;
			data[68961] <= 8'h10 ;
			data[68962] <= 8'h10 ;
			data[68963] <= 8'h10 ;
			data[68964] <= 8'h10 ;
			data[68965] <= 8'h10 ;
			data[68966] <= 8'h10 ;
			data[68967] <= 8'h10 ;
			data[68968] <= 8'h10 ;
			data[68969] <= 8'h10 ;
			data[68970] <= 8'h10 ;
			data[68971] <= 8'h10 ;
			data[68972] <= 8'h10 ;
			data[68973] <= 8'h10 ;
			data[68974] <= 8'h10 ;
			data[68975] <= 8'h10 ;
			data[68976] <= 8'h10 ;
			data[68977] <= 8'h10 ;
			data[68978] <= 8'h10 ;
			data[68979] <= 8'h10 ;
			data[68980] <= 8'h10 ;
			data[68981] <= 8'h10 ;
			data[68982] <= 8'h10 ;
			data[68983] <= 8'h10 ;
			data[68984] <= 8'h10 ;
			data[68985] <= 8'h10 ;
			data[68986] <= 8'h10 ;
			data[68987] <= 8'h10 ;
			data[68988] <= 8'h10 ;
			data[68989] <= 8'h10 ;
			data[68990] <= 8'h10 ;
			data[68991] <= 8'h10 ;
			data[68992] <= 8'h10 ;
			data[68993] <= 8'h10 ;
			data[68994] <= 8'h10 ;
			data[68995] <= 8'h10 ;
			data[68996] <= 8'h10 ;
			data[68997] <= 8'h10 ;
			data[68998] <= 8'h10 ;
			data[68999] <= 8'h10 ;
			data[69000] <= 8'h10 ;
			data[69001] <= 8'h10 ;
			data[69002] <= 8'h10 ;
			data[69003] <= 8'h10 ;
			data[69004] <= 8'h10 ;
			data[69005] <= 8'h10 ;
			data[69006] <= 8'h10 ;
			data[69007] <= 8'h10 ;
			data[69008] <= 8'h10 ;
			data[69009] <= 8'h10 ;
			data[69010] <= 8'h10 ;
			data[69011] <= 8'h10 ;
			data[69012] <= 8'h10 ;
			data[69013] <= 8'h10 ;
			data[69014] <= 8'h10 ;
			data[69015] <= 8'h10 ;
			data[69016] <= 8'h10 ;
			data[69017] <= 8'h10 ;
			data[69018] <= 8'h10 ;
			data[69019] <= 8'h10 ;
			data[69020] <= 8'h10 ;
			data[69021] <= 8'h10 ;
			data[69022] <= 8'h10 ;
			data[69023] <= 8'h10 ;
			data[69024] <= 8'h10 ;
			data[69025] <= 8'h10 ;
			data[69026] <= 8'h10 ;
			data[69027] <= 8'h10 ;
			data[69028] <= 8'h10 ;
			data[69029] <= 8'h10 ;
			data[69030] <= 8'h10 ;
			data[69031] <= 8'h10 ;
			data[69032] <= 8'h10 ;
			data[69033] <= 8'h10 ;
			data[69034] <= 8'h10 ;
			data[69035] <= 8'h10 ;
			data[69036] <= 8'h10 ;
			data[69037] <= 8'h10 ;
			data[69038] <= 8'h10 ;
			data[69039] <= 8'h10 ;
			data[69040] <= 8'h10 ;
			data[69041] <= 8'h10 ;
			data[69042] <= 8'h10 ;
			data[69043] <= 8'h10 ;
			data[69044] <= 8'h10 ;
			data[69045] <= 8'h10 ;
			data[69046] <= 8'h10 ;
			data[69047] <= 8'h10 ;
			data[69048] <= 8'h10 ;
			data[69049] <= 8'h10 ;
			data[69050] <= 8'h10 ;
			data[69051] <= 8'h10 ;
			data[69052] <= 8'h10 ;
			data[69053] <= 8'h10 ;
			data[69054] <= 8'h10 ;
			data[69055] <= 8'h10 ;
			data[69056] <= 8'h10 ;
			data[69057] <= 8'h10 ;
			data[69058] <= 8'h10 ;
			data[69059] <= 8'h10 ;
			data[69060] <= 8'h10 ;
			data[69061] <= 8'h10 ;
			data[69062] <= 8'h10 ;
			data[69063] <= 8'h10 ;
			data[69064] <= 8'h10 ;
			data[69065] <= 8'h10 ;
			data[69066] <= 8'h10 ;
			data[69067] <= 8'h10 ;
			data[69068] <= 8'h10 ;
			data[69069] <= 8'h10 ;
			data[69070] <= 8'h10 ;
			data[69071] <= 8'h10 ;
			data[69072] <= 8'h10 ;
			data[69073] <= 8'h10 ;
			data[69074] <= 8'h10 ;
			data[69075] <= 8'h10 ;
			data[69076] <= 8'h10 ;
			data[69077] <= 8'h10 ;
			data[69078] <= 8'h10 ;
			data[69079] <= 8'h10 ;
			data[69080] <= 8'h10 ;
			data[69081] <= 8'h10 ;
			data[69082] <= 8'h10 ;
			data[69083] <= 8'h10 ;
			data[69084] <= 8'h10 ;
			data[69085] <= 8'h10 ;
			data[69086] <= 8'h10 ;
			data[69087] <= 8'h10 ;
			data[69088] <= 8'h10 ;
			data[69089] <= 8'h10 ;
			data[69090] <= 8'h10 ;
			data[69091] <= 8'h10 ;
			data[69092] <= 8'h10 ;
			data[69093] <= 8'h10 ;
			data[69094] <= 8'h10 ;
			data[69095] <= 8'h10 ;
			data[69096] <= 8'h10 ;
			data[69097] <= 8'h10 ;
			data[69098] <= 8'h10 ;
			data[69099] <= 8'h10 ;
			data[69100] <= 8'h10 ;
			data[69101] <= 8'h10 ;
			data[69102] <= 8'h10 ;
			data[69103] <= 8'h10 ;
			data[69104] <= 8'h10 ;
			data[69105] <= 8'h10 ;
			data[69106] <= 8'h10 ;
			data[69107] <= 8'h10 ;
			data[69108] <= 8'h10 ;
			data[69109] <= 8'h10 ;
			data[69110] <= 8'h10 ;
			data[69111] <= 8'h10 ;
			data[69112] <= 8'h10 ;
			data[69113] <= 8'h10 ;
			data[69114] <= 8'h10 ;
			data[69115] <= 8'h10 ;
			data[69116] <= 8'h10 ;
			data[69117] <= 8'h10 ;
			data[69118] <= 8'h10 ;
			data[69119] <= 8'h10 ;
			data[69120] <= 8'h10 ;
			data[69121] <= 8'h10 ;
			data[69122] <= 8'h10 ;
			data[69123] <= 8'h10 ;
			data[69124] <= 8'h10 ;
			data[69125] <= 8'h10 ;
			data[69126] <= 8'h10 ;
			data[69127] <= 8'h10 ;
			data[69128] <= 8'h10 ;
			data[69129] <= 8'h10 ;
			data[69130] <= 8'h10 ;
			data[69131] <= 8'h10 ;
			data[69132] <= 8'h10 ;
			data[69133] <= 8'h10 ;
			data[69134] <= 8'h10 ;
			data[69135] <= 8'h10 ;
			data[69136] <= 8'h10 ;
			data[69137] <= 8'h10 ;
			data[69138] <= 8'h10 ;
			data[69139] <= 8'h10 ;
			data[69140] <= 8'h10 ;
			data[69141] <= 8'h10 ;
			data[69142] <= 8'h10 ;
			data[69143] <= 8'h10 ;
			data[69144] <= 8'h10 ;
			data[69145] <= 8'h10 ;
			data[69146] <= 8'h10 ;
			data[69147] <= 8'h10 ;
			data[69148] <= 8'h10 ;
			data[69149] <= 8'h10 ;
			data[69150] <= 8'h10 ;
			data[69151] <= 8'h10 ;
			data[69152] <= 8'h10 ;
			data[69153] <= 8'h10 ;
			data[69154] <= 8'h10 ;
			data[69155] <= 8'h10 ;
			data[69156] <= 8'h10 ;
			data[69157] <= 8'h10 ;
			data[69158] <= 8'h10 ;
			data[69159] <= 8'h10 ;
			data[69160] <= 8'h10 ;
			data[69161] <= 8'h10 ;
			data[69162] <= 8'h10 ;
			data[69163] <= 8'h10 ;
			data[69164] <= 8'h10 ;
			data[69165] <= 8'h10 ;
			data[69166] <= 8'h10 ;
			data[69167] <= 8'h10 ;
			data[69168] <= 8'h10 ;
			data[69169] <= 8'h10 ;
			data[69170] <= 8'h10 ;
			data[69171] <= 8'h10 ;
			data[69172] <= 8'h10 ;
			data[69173] <= 8'h10 ;
			data[69174] <= 8'h10 ;
			data[69175] <= 8'h10 ;
			data[69176] <= 8'h10 ;
			data[69177] <= 8'h10 ;
			data[69178] <= 8'h10 ;
			data[69179] <= 8'h10 ;
			data[69180] <= 8'h10 ;
			data[69181] <= 8'h10 ;
			data[69182] <= 8'h10 ;
			data[69183] <= 8'h10 ;
			data[69184] <= 8'h10 ;
			data[69185] <= 8'h10 ;
			data[69186] <= 8'h10 ;
			data[69187] <= 8'h10 ;
			data[69188] <= 8'h10 ;
			data[69189] <= 8'h10 ;
			data[69190] <= 8'h10 ;
			data[69191] <= 8'h10 ;
			data[69192] <= 8'h10 ;
			data[69193] <= 8'h10 ;
			data[69194] <= 8'h10 ;
			data[69195] <= 8'h10 ;
			data[69196] <= 8'h10 ;
			data[69197] <= 8'h10 ;
			data[69198] <= 8'h10 ;
			data[69199] <= 8'h10 ;
			data[69200] <= 8'h10 ;
			data[69201] <= 8'h10 ;
			data[69202] <= 8'h10 ;
			data[69203] <= 8'h10 ;
			data[69204] <= 8'h10 ;
			data[69205] <= 8'h10 ;
			data[69206] <= 8'h10 ;
			data[69207] <= 8'h10 ;
			data[69208] <= 8'h10 ;
			data[69209] <= 8'h10 ;
			data[69210] <= 8'h10 ;
			data[69211] <= 8'h10 ;
			data[69212] <= 8'h10 ;
			data[69213] <= 8'h10 ;
			data[69214] <= 8'h10 ;
			data[69215] <= 8'h10 ;
			data[69216] <= 8'h10 ;
			data[69217] <= 8'h10 ;
			data[69218] <= 8'h10 ;
			data[69219] <= 8'h10 ;
			data[69220] <= 8'h10 ;
			data[69221] <= 8'h10 ;
			data[69222] <= 8'h10 ;
			data[69223] <= 8'h10 ;
			data[69224] <= 8'h10 ;
			data[69225] <= 8'h10 ;
			data[69226] <= 8'h10 ;
			data[69227] <= 8'h10 ;
			data[69228] <= 8'h10 ;
			data[69229] <= 8'h10 ;
			data[69230] <= 8'h10 ;
			data[69231] <= 8'h10 ;
			data[69232] <= 8'h10 ;
			data[69233] <= 8'h10 ;
			data[69234] <= 8'h10 ;
			data[69235] <= 8'h10 ;
			data[69236] <= 8'h10 ;
			data[69237] <= 8'h10 ;
			data[69238] <= 8'h10 ;
			data[69239] <= 8'h10 ;
			data[69240] <= 8'h10 ;
			data[69241] <= 8'h10 ;
			data[69242] <= 8'h10 ;
			data[69243] <= 8'h10 ;
			data[69244] <= 8'h10 ;
			data[69245] <= 8'h10 ;
			data[69246] <= 8'h10 ;
			data[69247] <= 8'h10 ;
			data[69248] <= 8'h10 ;
			data[69249] <= 8'h10 ;
			data[69250] <= 8'h10 ;
			data[69251] <= 8'h10 ;
			data[69252] <= 8'h10 ;
			data[69253] <= 8'h10 ;
			data[69254] <= 8'h10 ;
			data[69255] <= 8'h10 ;
			data[69256] <= 8'h10 ;
			data[69257] <= 8'h10 ;
			data[69258] <= 8'h10 ;
			data[69259] <= 8'h10 ;
			data[69260] <= 8'h10 ;
			data[69261] <= 8'h10 ;
			data[69262] <= 8'h10 ;
			data[69263] <= 8'h10 ;
			data[69264] <= 8'h10 ;
			data[69265] <= 8'h10 ;
			data[69266] <= 8'h10 ;
			data[69267] <= 8'h10 ;
			data[69268] <= 8'h10 ;
			data[69269] <= 8'h10 ;
			data[69270] <= 8'h10 ;
			data[69271] <= 8'h10 ;
			data[69272] <= 8'h10 ;
			data[69273] <= 8'h10 ;
			data[69274] <= 8'h10 ;
			data[69275] <= 8'h10 ;
			data[69276] <= 8'h10 ;
			data[69277] <= 8'h10 ;
			data[69278] <= 8'h10 ;
			data[69279] <= 8'h10 ;
			data[69280] <= 8'h10 ;
			data[69281] <= 8'h10 ;
			data[69282] <= 8'h10 ;
			data[69283] <= 8'h10 ;
			data[69284] <= 8'h10 ;
			data[69285] <= 8'h10 ;
			data[69286] <= 8'h10 ;
			data[69287] <= 8'h10 ;
			data[69288] <= 8'h10 ;
			data[69289] <= 8'h10 ;
			data[69290] <= 8'h10 ;
			data[69291] <= 8'h10 ;
			data[69292] <= 8'h10 ;
			data[69293] <= 8'h10 ;
			data[69294] <= 8'h10 ;
			data[69295] <= 8'h10 ;
			data[69296] <= 8'h10 ;
			data[69297] <= 8'h10 ;
			data[69298] <= 8'h10 ;
			data[69299] <= 8'h10 ;
			data[69300] <= 8'h10 ;
			data[69301] <= 8'h10 ;
			data[69302] <= 8'h10 ;
			data[69303] <= 8'h10 ;
			data[69304] <= 8'h10 ;
			data[69305] <= 8'h10 ;
			data[69306] <= 8'h10 ;
			data[69307] <= 8'h10 ;
			data[69308] <= 8'h10 ;
			data[69309] <= 8'h10 ;
			data[69310] <= 8'h10 ;
			data[69311] <= 8'h10 ;
			data[69312] <= 8'h10 ;
			data[69313] <= 8'h10 ;
			data[69314] <= 8'h10 ;
			data[69315] <= 8'h10 ;
			data[69316] <= 8'h10 ;
			data[69317] <= 8'h10 ;
			data[69318] <= 8'h10 ;
			data[69319] <= 8'h10 ;
			data[69320] <= 8'h10 ;
			data[69321] <= 8'h10 ;
			data[69322] <= 8'h10 ;
			data[69323] <= 8'h10 ;
			data[69324] <= 8'h10 ;
			data[69325] <= 8'h10 ;
			data[69326] <= 8'h10 ;
			data[69327] <= 8'h10 ;
			data[69328] <= 8'h10 ;
			data[69329] <= 8'h10 ;
			data[69330] <= 8'h10 ;
			data[69331] <= 8'h10 ;
			data[69332] <= 8'h10 ;
			data[69333] <= 8'h10 ;
			data[69334] <= 8'h10 ;
			data[69335] <= 8'h10 ;
			data[69336] <= 8'h10 ;
			data[69337] <= 8'h10 ;
			data[69338] <= 8'h10 ;
			data[69339] <= 8'h10 ;
			data[69340] <= 8'h10 ;
			data[69341] <= 8'h10 ;
			data[69342] <= 8'h10 ;
			data[69343] <= 8'h10 ;
			data[69344] <= 8'h10 ;
			data[69345] <= 8'h10 ;
			data[69346] <= 8'h10 ;
			data[69347] <= 8'h10 ;
			data[69348] <= 8'h10 ;
			data[69349] <= 8'h10 ;
			data[69350] <= 8'h10 ;
			data[69351] <= 8'h10 ;
			data[69352] <= 8'h10 ;
			data[69353] <= 8'h10 ;
			data[69354] <= 8'h10 ;
			data[69355] <= 8'h10 ;
			data[69356] <= 8'h10 ;
			data[69357] <= 8'h10 ;
			data[69358] <= 8'h10 ;
			data[69359] <= 8'h10 ;
			data[69360] <= 8'h10 ;
			data[69361] <= 8'h10 ;
			data[69362] <= 8'h10 ;
			data[69363] <= 8'h10 ;
			data[69364] <= 8'h10 ;
			data[69365] <= 8'h10 ;
			data[69366] <= 8'h10 ;
			data[69367] <= 8'h10 ;
			data[69368] <= 8'h10 ;
			data[69369] <= 8'h10 ;
			data[69370] <= 8'h10 ;
			data[69371] <= 8'h10 ;
			data[69372] <= 8'h10 ;
			data[69373] <= 8'h10 ;
			data[69374] <= 8'h10 ;
			data[69375] <= 8'h10 ;
			data[69376] <= 8'h10 ;
			data[69377] <= 8'h10 ;
			data[69378] <= 8'h10 ;
			data[69379] <= 8'h10 ;
			data[69380] <= 8'h10 ;
			data[69381] <= 8'h10 ;
			data[69382] <= 8'h10 ;
			data[69383] <= 8'h10 ;
			data[69384] <= 8'h10 ;
			data[69385] <= 8'h10 ;
			data[69386] <= 8'h10 ;
			data[69387] <= 8'h10 ;
			data[69388] <= 8'h10 ;
			data[69389] <= 8'h10 ;
			data[69390] <= 8'h10 ;
			data[69391] <= 8'h10 ;
			data[69392] <= 8'h10 ;
			data[69393] <= 8'h10 ;
			data[69394] <= 8'h10 ;
			data[69395] <= 8'h10 ;
			data[69396] <= 8'h10 ;
			data[69397] <= 8'h10 ;
			data[69398] <= 8'h10 ;
			data[69399] <= 8'h10 ;
			data[69400] <= 8'h10 ;
			data[69401] <= 8'h10 ;
			data[69402] <= 8'h10 ;
			data[69403] <= 8'h10 ;
			data[69404] <= 8'h10 ;
			data[69405] <= 8'h10 ;
			data[69406] <= 8'h10 ;
			data[69407] <= 8'h10 ;
			data[69408] <= 8'h10 ;
			data[69409] <= 8'h10 ;
			data[69410] <= 8'h10 ;
			data[69411] <= 8'h10 ;
			data[69412] <= 8'h10 ;
			data[69413] <= 8'h10 ;
			data[69414] <= 8'h10 ;
			data[69415] <= 8'h10 ;
			data[69416] <= 8'h10 ;
			data[69417] <= 8'h10 ;
			data[69418] <= 8'h10 ;
			data[69419] <= 8'h10 ;
			data[69420] <= 8'h10 ;
			data[69421] <= 8'h10 ;
			data[69422] <= 8'h10 ;
			data[69423] <= 8'h10 ;
			data[69424] <= 8'h10 ;
			data[69425] <= 8'h10 ;
			data[69426] <= 8'h10 ;
			data[69427] <= 8'h10 ;
			data[69428] <= 8'h10 ;
			data[69429] <= 8'h10 ;
			data[69430] <= 8'h10 ;
			data[69431] <= 8'h10 ;
			data[69432] <= 8'h10 ;
			data[69433] <= 8'h10 ;
			data[69434] <= 8'h10 ;
			data[69435] <= 8'h10 ;
			data[69436] <= 8'h10 ;
			data[69437] <= 8'h10 ;
			data[69438] <= 8'h10 ;
			data[69439] <= 8'h10 ;
			data[69440] <= 8'h10 ;
			data[69441] <= 8'h10 ;
			data[69442] <= 8'h10 ;
			data[69443] <= 8'h10 ;
			data[69444] <= 8'h10 ;
			data[69445] <= 8'h10 ;
			data[69446] <= 8'h10 ;
			data[69447] <= 8'h10 ;
			data[69448] <= 8'h10 ;
			data[69449] <= 8'h10 ;
			data[69450] <= 8'h10 ;
			data[69451] <= 8'h10 ;
			data[69452] <= 8'h10 ;
			data[69453] <= 8'h10 ;
			data[69454] <= 8'h10 ;
			data[69455] <= 8'h10 ;
			data[69456] <= 8'h10 ;
			data[69457] <= 8'h10 ;
			data[69458] <= 8'h10 ;
			data[69459] <= 8'h10 ;
			data[69460] <= 8'h10 ;
			data[69461] <= 8'h10 ;
			data[69462] <= 8'h10 ;
			data[69463] <= 8'h10 ;
			data[69464] <= 8'h10 ;
			data[69465] <= 8'h10 ;
			data[69466] <= 8'h10 ;
			data[69467] <= 8'h10 ;
			data[69468] <= 8'h10 ;
			data[69469] <= 8'h10 ;
			data[69470] <= 8'h10 ;
			data[69471] <= 8'h10 ;
			data[69472] <= 8'h10 ;
			data[69473] <= 8'h10 ;
			data[69474] <= 8'h10 ;
			data[69475] <= 8'h10 ;
			data[69476] <= 8'h10 ;
			data[69477] <= 8'h10 ;
			data[69478] <= 8'h10 ;
			data[69479] <= 8'h10 ;
			data[69480] <= 8'h10 ;
			data[69481] <= 8'h10 ;
			data[69482] <= 8'h10 ;
			data[69483] <= 8'h10 ;
			data[69484] <= 8'h10 ;
			data[69485] <= 8'h10 ;
			data[69486] <= 8'h10 ;
			data[69487] <= 8'h10 ;
			data[69488] <= 8'h10 ;
			data[69489] <= 8'h10 ;
			data[69490] <= 8'h10 ;
			data[69491] <= 8'h10 ;
			data[69492] <= 8'h10 ;
			data[69493] <= 8'h10 ;
			data[69494] <= 8'h10 ;
			data[69495] <= 8'h10 ;
			data[69496] <= 8'h10 ;
			data[69497] <= 8'h10 ;
			data[69498] <= 8'h10 ;
			data[69499] <= 8'h10 ;
			data[69500] <= 8'h10 ;
			data[69501] <= 8'h10 ;
			data[69502] <= 8'h10 ;
			data[69503] <= 8'h10 ;
			data[69504] <= 8'h10 ;
			data[69505] <= 8'h10 ;
			data[69506] <= 8'h10 ;
			data[69507] <= 8'h10 ;
			data[69508] <= 8'h10 ;
			data[69509] <= 8'h10 ;
			data[69510] <= 8'h10 ;
			data[69511] <= 8'h10 ;
			data[69512] <= 8'h10 ;
			data[69513] <= 8'h10 ;
			data[69514] <= 8'h10 ;
			data[69515] <= 8'h10 ;
			data[69516] <= 8'h10 ;
			data[69517] <= 8'h10 ;
			data[69518] <= 8'h10 ;
			data[69519] <= 8'h10 ;
			data[69520] <= 8'h10 ;
			data[69521] <= 8'h10 ;
			data[69522] <= 8'h10 ;
			data[69523] <= 8'h10 ;
			data[69524] <= 8'h10 ;
			data[69525] <= 8'h10 ;
			data[69526] <= 8'h10 ;
			data[69527] <= 8'h10 ;
			data[69528] <= 8'h10 ;
			data[69529] <= 8'h10 ;
			data[69530] <= 8'h10 ;
			data[69531] <= 8'h10 ;
			data[69532] <= 8'h10 ;
			data[69533] <= 8'h10 ;
			data[69534] <= 8'h10 ;
			data[69535] <= 8'h10 ;
			data[69536] <= 8'h10 ;
			data[69537] <= 8'h10 ;
			data[69538] <= 8'h10 ;
			data[69539] <= 8'h10 ;
			data[69540] <= 8'h10 ;
			data[69541] <= 8'h10 ;
			data[69542] <= 8'h10 ;
			data[69543] <= 8'h10 ;
			data[69544] <= 8'h10 ;
			data[69545] <= 8'h10 ;
			data[69546] <= 8'h10 ;
			data[69547] <= 8'h10 ;
			data[69548] <= 8'h10 ;
			data[69549] <= 8'h10 ;
			data[69550] <= 8'h10 ;
			data[69551] <= 8'h10 ;
			data[69552] <= 8'h10 ;
			data[69553] <= 8'h10 ;
			data[69554] <= 8'h10 ;
			data[69555] <= 8'h10 ;
			data[69556] <= 8'h10 ;
			data[69557] <= 8'h10 ;
			data[69558] <= 8'h10 ;
			data[69559] <= 8'h10 ;
			data[69560] <= 8'h10 ;
			data[69561] <= 8'h10 ;
			data[69562] <= 8'h10 ;
			data[69563] <= 8'h10 ;
			data[69564] <= 8'h10 ;
			data[69565] <= 8'h10 ;
			data[69566] <= 8'h10 ;
			data[69567] <= 8'h10 ;
			data[69568] <= 8'h10 ;
			data[69569] <= 8'h10 ;
			data[69570] <= 8'h10 ;
			data[69571] <= 8'h10 ;
			data[69572] <= 8'h10 ;
			data[69573] <= 8'h10 ;
			data[69574] <= 8'h10 ;
			data[69575] <= 8'h10 ;
			data[69576] <= 8'h10 ;
			data[69577] <= 8'h10 ;
			data[69578] <= 8'h10 ;
			data[69579] <= 8'h10 ;
			data[69580] <= 8'h10 ;
			data[69581] <= 8'h10 ;
			data[69582] <= 8'h10 ;
			data[69583] <= 8'h10 ;
			data[69584] <= 8'h10 ;
			data[69585] <= 8'h10 ;
			data[69586] <= 8'h10 ;
			data[69587] <= 8'h10 ;
			data[69588] <= 8'h10 ;
			data[69589] <= 8'h10 ;
			data[69590] <= 8'h10 ;
			data[69591] <= 8'h10 ;
			data[69592] <= 8'h10 ;
			data[69593] <= 8'h10 ;
			data[69594] <= 8'h10 ;
			data[69595] <= 8'h10 ;
			data[69596] <= 8'h10 ;
			data[69597] <= 8'h10 ;
			data[69598] <= 8'h10 ;
			data[69599] <= 8'h10 ;
			data[69600] <= 8'h10 ;
			data[69601] <= 8'h10 ;
			data[69602] <= 8'h10 ;
			data[69603] <= 8'h10 ;
			data[69604] <= 8'h10 ;
			data[69605] <= 8'h10 ;
			data[69606] <= 8'h10 ;
			data[69607] <= 8'h10 ;
			data[69608] <= 8'h10 ;
			data[69609] <= 8'h10 ;
			data[69610] <= 8'h10 ;
			data[69611] <= 8'h10 ;
			data[69612] <= 8'h10 ;
			data[69613] <= 8'h10 ;
			data[69614] <= 8'h10 ;
			data[69615] <= 8'h10 ;
			data[69616] <= 8'h10 ;
			data[69617] <= 8'h10 ;
			data[69618] <= 8'h10 ;
			data[69619] <= 8'h10 ;
			data[69620] <= 8'h10 ;
			data[69621] <= 8'h10 ;
			data[69622] <= 8'h10 ;
			data[69623] <= 8'h10 ;
			data[69624] <= 8'h10 ;
			data[69625] <= 8'h10 ;
			data[69626] <= 8'h10 ;
			data[69627] <= 8'h10 ;
			data[69628] <= 8'h10 ;
			data[69629] <= 8'h10 ;
			data[69630] <= 8'h10 ;
			data[69631] <= 8'h10 ;
			data[69632] <= 8'h10 ;
			data[69633] <= 8'h10 ;
			data[69634] <= 8'h10 ;
			data[69635] <= 8'h10 ;
			data[69636] <= 8'h10 ;
			data[69637] <= 8'h10 ;
			data[69638] <= 8'h10 ;
			data[69639] <= 8'h10 ;
			data[69640] <= 8'h10 ;
			data[69641] <= 8'h10 ;
			data[69642] <= 8'h10 ;
			data[69643] <= 8'h10 ;
			data[69644] <= 8'h10 ;
			data[69645] <= 8'h10 ;
			data[69646] <= 8'h10 ;
			data[69647] <= 8'h10 ;
			data[69648] <= 8'h10 ;
			data[69649] <= 8'h10 ;
			data[69650] <= 8'h10 ;
			data[69651] <= 8'h10 ;
			data[69652] <= 8'h10 ;
			data[69653] <= 8'h10 ;
			data[69654] <= 8'h10 ;
			data[69655] <= 8'h10 ;
			data[69656] <= 8'h10 ;
			data[69657] <= 8'h10 ;
			data[69658] <= 8'h10 ;
			data[69659] <= 8'h10 ;
			data[69660] <= 8'h10 ;
			data[69661] <= 8'h10 ;
			data[69662] <= 8'h10 ;
			data[69663] <= 8'h10 ;
			data[69664] <= 8'h10 ;
			data[69665] <= 8'h10 ;
			data[69666] <= 8'h10 ;
			data[69667] <= 8'h10 ;
			data[69668] <= 8'h10 ;
			data[69669] <= 8'h10 ;
			data[69670] <= 8'h10 ;
			data[69671] <= 8'h10 ;
			data[69672] <= 8'h10 ;
			data[69673] <= 8'h10 ;
			data[69674] <= 8'h10 ;
			data[69675] <= 8'h10 ;
			data[69676] <= 8'h10 ;
			data[69677] <= 8'h10 ;
			data[69678] <= 8'h10 ;
			data[69679] <= 8'h10 ;
			data[69680] <= 8'h10 ;
			data[69681] <= 8'h10 ;
			data[69682] <= 8'h10 ;
			data[69683] <= 8'h10 ;
			data[69684] <= 8'h10 ;
			data[69685] <= 8'h10 ;
			data[69686] <= 8'h10 ;
			data[69687] <= 8'h10 ;
			data[69688] <= 8'h10 ;
			data[69689] <= 8'h10 ;
			data[69690] <= 8'h10 ;
			data[69691] <= 8'h10 ;
			data[69692] <= 8'h10 ;
			data[69693] <= 8'h10 ;
			data[69694] <= 8'h10 ;
			data[69695] <= 8'h10 ;
			data[69696] <= 8'h10 ;
			data[69697] <= 8'h10 ;
			data[69698] <= 8'h10 ;
			data[69699] <= 8'h10 ;
			data[69700] <= 8'h10 ;
			data[69701] <= 8'h10 ;
			data[69702] <= 8'h10 ;
			data[69703] <= 8'h10 ;
			data[69704] <= 8'h10 ;
			data[69705] <= 8'h10 ;
			data[69706] <= 8'h10 ;
			data[69707] <= 8'h10 ;
			data[69708] <= 8'h10 ;
			data[69709] <= 8'h10 ;
			data[69710] <= 8'h10 ;
			data[69711] <= 8'h10 ;
			data[69712] <= 8'h10 ;
			data[69713] <= 8'h10 ;
			data[69714] <= 8'h10 ;
			data[69715] <= 8'h10 ;
			data[69716] <= 8'h10 ;
			data[69717] <= 8'h10 ;
			data[69718] <= 8'h10 ;
			data[69719] <= 8'h10 ;
			data[69720] <= 8'h10 ;
			data[69721] <= 8'h10 ;
			data[69722] <= 8'h10 ;
			data[69723] <= 8'h10 ;
			data[69724] <= 8'h10 ;
			data[69725] <= 8'h10 ;
			data[69726] <= 8'h10 ;
			data[69727] <= 8'h10 ;
			data[69728] <= 8'h10 ;
			data[69729] <= 8'h10 ;
			data[69730] <= 8'h10 ;
			data[69731] <= 8'h10 ;
			data[69732] <= 8'h10 ;
			data[69733] <= 8'h10 ;
			data[69734] <= 8'h10 ;
			data[69735] <= 8'h10 ;
			data[69736] <= 8'h10 ;
			data[69737] <= 8'h10 ;
			data[69738] <= 8'h10 ;
			data[69739] <= 8'h10 ;
			data[69740] <= 8'h10 ;
			data[69741] <= 8'h10 ;
			data[69742] <= 8'h10 ;
			data[69743] <= 8'h10 ;
			data[69744] <= 8'h10 ;
			data[69745] <= 8'h10 ;
			data[69746] <= 8'h10 ;
			data[69747] <= 8'h10 ;
			data[69748] <= 8'h10 ;
			data[69749] <= 8'h10 ;
			data[69750] <= 8'h10 ;
			data[69751] <= 8'h10 ;
			data[69752] <= 8'h10 ;
			data[69753] <= 8'h10 ;
			data[69754] <= 8'h10 ;
			data[69755] <= 8'h10 ;
			data[69756] <= 8'h10 ;
			data[69757] <= 8'h10 ;
			data[69758] <= 8'h10 ;
			data[69759] <= 8'h10 ;
			data[69760] <= 8'h10 ;
			data[69761] <= 8'h10 ;
			data[69762] <= 8'h10 ;
			data[69763] <= 8'h10 ;
			data[69764] <= 8'h10 ;
			data[69765] <= 8'h10 ;
			data[69766] <= 8'h10 ;
			data[69767] <= 8'h10 ;
			data[69768] <= 8'h10 ;
			data[69769] <= 8'h10 ;
			data[69770] <= 8'h10 ;
			data[69771] <= 8'h10 ;
			data[69772] <= 8'h10 ;
			data[69773] <= 8'h10 ;
			data[69774] <= 8'h10 ;
			data[69775] <= 8'h10 ;
			data[69776] <= 8'h10 ;
			data[69777] <= 8'h10 ;
			data[69778] <= 8'h10 ;
			data[69779] <= 8'h10 ;
			data[69780] <= 8'h10 ;
			data[69781] <= 8'h10 ;
			data[69782] <= 8'h10 ;
			data[69783] <= 8'h10 ;
			data[69784] <= 8'h10 ;
			data[69785] <= 8'h10 ;
			data[69786] <= 8'h10 ;
			data[69787] <= 8'h10 ;
			data[69788] <= 8'h10 ;
			data[69789] <= 8'h10 ;
			data[69790] <= 8'h10 ;
			data[69791] <= 8'h10 ;
			data[69792] <= 8'h10 ;
			data[69793] <= 8'h10 ;
			data[69794] <= 8'h10 ;
			data[69795] <= 8'h10 ;
			data[69796] <= 8'h10 ;
			data[69797] <= 8'h10 ;
			data[69798] <= 8'h10 ;
			data[69799] <= 8'h10 ;
			data[69800] <= 8'h10 ;
			data[69801] <= 8'h10 ;
			data[69802] <= 8'h10 ;
			data[69803] <= 8'h10 ;
			data[69804] <= 8'h10 ;
			data[69805] <= 8'h10 ;
			data[69806] <= 8'h10 ;
			data[69807] <= 8'h10 ;
			data[69808] <= 8'h10 ;
			data[69809] <= 8'h10 ;
			data[69810] <= 8'h10 ;
			data[69811] <= 8'h10 ;
			data[69812] <= 8'h10 ;
			data[69813] <= 8'h10 ;
			data[69814] <= 8'h10 ;
			data[69815] <= 8'h10 ;
			data[69816] <= 8'h10 ;
			data[69817] <= 8'h10 ;
			data[69818] <= 8'h10 ;
			data[69819] <= 8'h10 ;
			data[69820] <= 8'h10 ;
			data[69821] <= 8'h10 ;
			data[69822] <= 8'h10 ;
			data[69823] <= 8'h10 ;
			data[69824] <= 8'h10 ;
			data[69825] <= 8'h10 ;
			data[69826] <= 8'h10 ;
			data[69827] <= 8'h10 ;
			data[69828] <= 8'h10 ;
			data[69829] <= 8'h10 ;
			data[69830] <= 8'h10 ;
			data[69831] <= 8'h10 ;
			data[69832] <= 8'h10 ;
			data[69833] <= 8'h10 ;
			data[69834] <= 8'h10 ;
			data[69835] <= 8'h10 ;
			data[69836] <= 8'h10 ;
			data[69837] <= 8'h10 ;
			data[69838] <= 8'h10 ;
			data[69839] <= 8'h10 ;
			data[69840] <= 8'h10 ;
			data[69841] <= 8'h10 ;
			data[69842] <= 8'h10 ;
			data[69843] <= 8'h10 ;
			data[69844] <= 8'h10 ;
			data[69845] <= 8'h10 ;
			data[69846] <= 8'h10 ;
			data[69847] <= 8'h10 ;
			data[69848] <= 8'h10 ;
			data[69849] <= 8'h10 ;
			data[69850] <= 8'h10 ;
			data[69851] <= 8'h10 ;
			data[69852] <= 8'h10 ;
			data[69853] <= 8'h10 ;
			data[69854] <= 8'h10 ;
			data[69855] <= 8'h10 ;
			data[69856] <= 8'h10 ;
			data[69857] <= 8'h10 ;
			data[69858] <= 8'h10 ;
			data[69859] <= 8'h10 ;
			data[69860] <= 8'h10 ;
			data[69861] <= 8'h10 ;
			data[69862] <= 8'h10 ;
			data[69863] <= 8'h10 ;
			data[69864] <= 8'h10 ;
			data[69865] <= 8'h10 ;
			data[69866] <= 8'h10 ;
			data[69867] <= 8'h10 ;
			data[69868] <= 8'h10 ;
			data[69869] <= 8'h10 ;
			data[69870] <= 8'h10 ;
			data[69871] <= 8'h10 ;
			data[69872] <= 8'h10 ;
			data[69873] <= 8'h10 ;
			data[69874] <= 8'h10 ;
			data[69875] <= 8'h10 ;
			data[69876] <= 8'h10 ;
			data[69877] <= 8'h10 ;
			data[69878] <= 8'h10 ;
			data[69879] <= 8'h10 ;
			data[69880] <= 8'h10 ;
			data[69881] <= 8'h10 ;
			data[69882] <= 8'h10 ;
			data[69883] <= 8'h10 ;
			data[69884] <= 8'h10 ;
			data[69885] <= 8'h10 ;
			data[69886] <= 8'h10 ;
			data[69887] <= 8'h10 ;
			data[69888] <= 8'h10 ;
			data[69889] <= 8'h10 ;
			data[69890] <= 8'h10 ;
			data[69891] <= 8'h10 ;
			data[69892] <= 8'h10 ;
			data[69893] <= 8'h10 ;
			data[69894] <= 8'h10 ;
			data[69895] <= 8'h10 ;
			data[69896] <= 8'h10 ;
			data[69897] <= 8'h10 ;
			data[69898] <= 8'h10 ;
			data[69899] <= 8'h10 ;
			data[69900] <= 8'h10 ;
			data[69901] <= 8'h10 ;
			data[69902] <= 8'h10 ;
			data[69903] <= 8'h10 ;
			data[69904] <= 8'h10 ;
			data[69905] <= 8'h10 ;
			data[69906] <= 8'h10 ;
			data[69907] <= 8'h10 ;
			data[69908] <= 8'h10 ;
			data[69909] <= 8'h10 ;
			data[69910] <= 8'h10 ;
			data[69911] <= 8'h10 ;
			data[69912] <= 8'h10 ;
			data[69913] <= 8'h10 ;
			data[69914] <= 8'h10 ;
			data[69915] <= 8'h10 ;
			data[69916] <= 8'h10 ;
			data[69917] <= 8'h10 ;
			data[69918] <= 8'h10 ;
			data[69919] <= 8'h10 ;
			data[69920] <= 8'h10 ;
			data[69921] <= 8'h10 ;
			data[69922] <= 8'h10 ;
			data[69923] <= 8'h10 ;
			data[69924] <= 8'h10 ;
			data[69925] <= 8'h10 ;
			data[69926] <= 8'h10 ;
			data[69927] <= 8'h10 ;
			data[69928] <= 8'h10 ;
			data[69929] <= 8'h10 ;
			data[69930] <= 8'h10 ;
			data[69931] <= 8'h10 ;
			data[69932] <= 8'h10 ;
			data[69933] <= 8'h10 ;
			data[69934] <= 8'h10 ;
			data[69935] <= 8'h10 ;
			data[69936] <= 8'h10 ;
			data[69937] <= 8'h10 ;
			data[69938] <= 8'h10 ;
			data[69939] <= 8'h10 ;
			data[69940] <= 8'h10 ;
			data[69941] <= 8'h10 ;
			data[69942] <= 8'h10 ;
			data[69943] <= 8'h10 ;
			data[69944] <= 8'h10 ;
			data[69945] <= 8'h10 ;
			data[69946] <= 8'h10 ;
			data[69947] <= 8'h10 ;
			data[69948] <= 8'h10 ;
			data[69949] <= 8'h10 ;
			data[69950] <= 8'h10 ;
			data[69951] <= 8'h10 ;
			data[69952] <= 8'h10 ;
			data[69953] <= 8'h10 ;
			data[69954] <= 8'h10 ;
			data[69955] <= 8'h10 ;
			data[69956] <= 8'h10 ;
			data[69957] <= 8'h10 ;
			data[69958] <= 8'h10 ;
			data[69959] <= 8'h10 ;
			data[69960] <= 8'h10 ;
			data[69961] <= 8'h10 ;
			data[69962] <= 8'h10 ;
			data[69963] <= 8'h10 ;
			data[69964] <= 8'h10 ;
			data[69965] <= 8'h10 ;
			data[69966] <= 8'h10 ;
			data[69967] <= 8'h10 ;
			data[69968] <= 8'h10 ;
			data[69969] <= 8'h10 ;
			data[69970] <= 8'h10 ;
			data[69971] <= 8'h10 ;
			data[69972] <= 8'h10 ;
			data[69973] <= 8'h10 ;
			data[69974] <= 8'h10 ;
			data[69975] <= 8'h10 ;
			data[69976] <= 8'h10 ;
			data[69977] <= 8'h10 ;
			data[69978] <= 8'h10 ;
			data[69979] <= 8'h10 ;
			data[69980] <= 8'h10 ;
			data[69981] <= 8'h10 ;
			data[69982] <= 8'h10 ;
			data[69983] <= 8'h10 ;
			data[69984] <= 8'h10 ;
			data[69985] <= 8'h10 ;
			data[69986] <= 8'h10 ;
			data[69987] <= 8'h10 ;
			data[69988] <= 8'h10 ;
			data[69989] <= 8'h10 ;
			data[69990] <= 8'h10 ;
			data[69991] <= 8'h10 ;
			data[69992] <= 8'h10 ;
			data[69993] <= 8'h10 ;
			data[69994] <= 8'h10 ;
			data[69995] <= 8'h10 ;
			data[69996] <= 8'h10 ;
			data[69997] <= 8'h10 ;
			data[69998] <= 8'h10 ;
			data[69999] <= 8'h10 ;
			data[70000] <= 8'h10 ;
			data[70001] <= 8'h10 ;
			data[70002] <= 8'h10 ;
			data[70003] <= 8'h10 ;
			data[70004] <= 8'h10 ;
			data[70005] <= 8'h10 ;
			data[70006] <= 8'h10 ;
			data[70007] <= 8'h10 ;
			data[70008] <= 8'h10 ;
			data[70009] <= 8'h10 ;
			data[70010] <= 8'h10 ;
			data[70011] <= 8'h10 ;
			data[70012] <= 8'h10 ;
			data[70013] <= 8'h10 ;
			data[70014] <= 8'h10 ;
			data[70015] <= 8'h10 ;
			data[70016] <= 8'h10 ;
			data[70017] <= 8'h10 ;
			data[70018] <= 8'h10 ;
			data[70019] <= 8'h10 ;
			data[70020] <= 8'h10 ;
			data[70021] <= 8'h10 ;
			data[70022] <= 8'h10 ;
			data[70023] <= 8'h10 ;
			data[70024] <= 8'h10 ;
			data[70025] <= 8'h10 ;
			data[70026] <= 8'h10 ;
			data[70027] <= 8'h10 ;
			data[70028] <= 8'h10 ;
			data[70029] <= 8'h10 ;
			data[70030] <= 8'h10 ;
			data[70031] <= 8'h10 ;
			data[70032] <= 8'h10 ;
			data[70033] <= 8'h10 ;
			data[70034] <= 8'h10 ;
			data[70035] <= 8'h10 ;
			data[70036] <= 8'h10 ;
			data[70037] <= 8'h10 ;
			data[70038] <= 8'h10 ;
			data[70039] <= 8'h10 ;
			data[70040] <= 8'h10 ;
			data[70041] <= 8'h10 ;
			data[70042] <= 8'h10 ;
			data[70043] <= 8'h10 ;
			data[70044] <= 8'h10 ;
			data[70045] <= 8'h10 ;
			data[70046] <= 8'h10 ;
			data[70047] <= 8'h10 ;
			data[70048] <= 8'h10 ;
			data[70049] <= 8'h10 ;
			data[70050] <= 8'h10 ;
			data[70051] <= 8'h10 ;
			data[70052] <= 8'h10 ;
			data[70053] <= 8'h10 ;
			data[70054] <= 8'h10 ;
			data[70055] <= 8'h10 ;
			data[70056] <= 8'h10 ;
			data[70057] <= 8'h10 ;
			data[70058] <= 8'h10 ;
			data[70059] <= 8'h10 ;
			data[70060] <= 8'h10 ;
			data[70061] <= 8'h10 ;
			data[70062] <= 8'h10 ;
			data[70063] <= 8'h10 ;
			data[70064] <= 8'h10 ;
			data[70065] <= 8'h10 ;
			data[70066] <= 8'h10 ;
			data[70067] <= 8'h10 ;
			data[70068] <= 8'h10 ;
			data[70069] <= 8'h10 ;
			data[70070] <= 8'h10 ;
			data[70071] <= 8'h10 ;
			data[70072] <= 8'h10 ;
			data[70073] <= 8'h10 ;
			data[70074] <= 8'h10 ;
			data[70075] <= 8'h10 ;
			data[70076] <= 8'h10 ;
			data[70077] <= 8'h10 ;
			data[70078] <= 8'h10 ;
			data[70079] <= 8'h10 ;
			data[70080] <= 8'h10 ;
			data[70081] <= 8'h10 ;
			data[70082] <= 8'h10 ;
			data[70083] <= 8'h10 ;
			data[70084] <= 8'h10 ;
			data[70085] <= 8'h10 ;
			data[70086] <= 8'h10 ;
			data[70087] <= 8'h10 ;
			data[70088] <= 8'h10 ;
			data[70089] <= 8'h10 ;
			data[70090] <= 8'h10 ;
			data[70091] <= 8'h10 ;
			data[70092] <= 8'h10 ;
			data[70093] <= 8'h10 ;
			data[70094] <= 8'h10 ;
			data[70095] <= 8'h10 ;
			data[70096] <= 8'h10 ;
			data[70097] <= 8'h10 ;
			data[70098] <= 8'h10 ;
			data[70099] <= 8'h10 ;
			data[70100] <= 8'h10 ;
			data[70101] <= 8'h10 ;
			data[70102] <= 8'h10 ;
			data[70103] <= 8'h10 ;
			data[70104] <= 8'h10 ;
			data[70105] <= 8'h10 ;
			data[70106] <= 8'h10 ;
			data[70107] <= 8'h10 ;
			data[70108] <= 8'h10 ;
			data[70109] <= 8'h10 ;
			data[70110] <= 8'h10 ;
			data[70111] <= 8'h10 ;
			data[70112] <= 8'h10 ;
			data[70113] <= 8'h10 ;
			data[70114] <= 8'h10 ;
			data[70115] <= 8'h10 ;
			data[70116] <= 8'h10 ;
			data[70117] <= 8'h10 ;
			data[70118] <= 8'h10 ;
			data[70119] <= 8'h10 ;
			data[70120] <= 8'h10 ;
			data[70121] <= 8'h10 ;
			data[70122] <= 8'h10 ;
			data[70123] <= 8'h10 ;
			data[70124] <= 8'h10 ;
			data[70125] <= 8'h10 ;
			data[70126] <= 8'h10 ;
			data[70127] <= 8'h10 ;
			data[70128] <= 8'h10 ;
			data[70129] <= 8'h10 ;
			data[70130] <= 8'h10 ;
			data[70131] <= 8'h10 ;
			data[70132] <= 8'h10 ;
			data[70133] <= 8'h10 ;
			data[70134] <= 8'h10 ;
			data[70135] <= 8'h10 ;
			data[70136] <= 8'h10 ;
			data[70137] <= 8'h10 ;
			data[70138] <= 8'h10 ;
			data[70139] <= 8'h10 ;
			data[70140] <= 8'h10 ;
			data[70141] <= 8'h10 ;
			data[70142] <= 8'h10 ;
			data[70143] <= 8'h10 ;
			data[70144] <= 8'h10 ;
			data[70145] <= 8'h10 ;
			data[70146] <= 8'h10 ;
			data[70147] <= 8'h10 ;
			data[70148] <= 8'h10 ;
			data[70149] <= 8'h10 ;
			data[70150] <= 8'h10 ;
			data[70151] <= 8'h10 ;
			data[70152] <= 8'h10 ;
			data[70153] <= 8'h10 ;
			data[70154] <= 8'h10 ;
			data[70155] <= 8'h10 ;
			data[70156] <= 8'h10 ;
			data[70157] <= 8'h10 ;
			data[70158] <= 8'h10 ;
			data[70159] <= 8'h10 ;
			data[70160] <= 8'h10 ;
			data[70161] <= 8'h10 ;
			data[70162] <= 8'h10 ;
			data[70163] <= 8'h10 ;
			data[70164] <= 8'h10 ;
			data[70165] <= 8'h10 ;
			data[70166] <= 8'h10 ;
			data[70167] <= 8'h10 ;
			data[70168] <= 8'h10 ;
			data[70169] <= 8'h10 ;
			data[70170] <= 8'h10 ;
			data[70171] <= 8'h10 ;
			data[70172] <= 8'h10 ;
			data[70173] <= 8'h10 ;
			data[70174] <= 8'h10 ;
			data[70175] <= 8'h10 ;
			data[70176] <= 8'h10 ;
			data[70177] <= 8'h10 ;
			data[70178] <= 8'h10 ;
			data[70179] <= 8'h10 ;
			data[70180] <= 8'h10 ;
			data[70181] <= 8'h10 ;
			data[70182] <= 8'h10 ;
			data[70183] <= 8'h10 ;
			data[70184] <= 8'h10 ;
			data[70185] <= 8'h10 ;
			data[70186] <= 8'h10 ;
			data[70187] <= 8'h10 ;
			data[70188] <= 8'h10 ;
			data[70189] <= 8'h10 ;
			data[70190] <= 8'h10 ;
			data[70191] <= 8'h10 ;
			data[70192] <= 8'h10 ;
			data[70193] <= 8'h10 ;
			data[70194] <= 8'h10 ;
			data[70195] <= 8'h10 ;
			data[70196] <= 8'h10 ;
			data[70197] <= 8'h10 ;
			data[70198] <= 8'h10 ;
			data[70199] <= 8'h10 ;
			data[70200] <= 8'h10 ;
			data[70201] <= 8'h10 ;
			data[70202] <= 8'h10 ;
			data[70203] <= 8'h10 ;
			data[70204] <= 8'h10 ;
			data[70205] <= 8'h10 ;
			data[70206] <= 8'h10 ;
			data[70207] <= 8'h10 ;
			data[70208] <= 8'h10 ;
			data[70209] <= 8'h10 ;
			data[70210] <= 8'h10 ;
			data[70211] <= 8'h10 ;
			data[70212] <= 8'h10 ;
			data[70213] <= 8'h10 ;
			data[70214] <= 8'h10 ;
			data[70215] <= 8'h10 ;
			data[70216] <= 8'h10 ;
			data[70217] <= 8'h10 ;
			data[70218] <= 8'h10 ;
			data[70219] <= 8'h10 ;
			data[70220] <= 8'h10 ;
			data[70221] <= 8'h10 ;
			data[70222] <= 8'h10 ;
			data[70223] <= 8'h10 ;
			data[70224] <= 8'h10 ;
			data[70225] <= 8'h10 ;
			data[70226] <= 8'h10 ;
			data[70227] <= 8'h10 ;
			data[70228] <= 8'h10 ;
			data[70229] <= 8'h10 ;
			data[70230] <= 8'h10 ;
			data[70231] <= 8'h10 ;
			data[70232] <= 8'h10 ;
			data[70233] <= 8'h10 ;
			data[70234] <= 8'h10 ;
			data[70235] <= 8'h10 ;
			data[70236] <= 8'h10 ;
			data[70237] <= 8'h10 ;
			data[70238] <= 8'h10 ;
			data[70239] <= 8'h10 ;
			data[70240] <= 8'h10 ;
			data[70241] <= 8'h10 ;
			data[70242] <= 8'h10 ;
			data[70243] <= 8'h10 ;
			data[70244] <= 8'h10 ;
			data[70245] <= 8'h10 ;
			data[70246] <= 8'h10 ;
			data[70247] <= 8'h10 ;
			data[70248] <= 8'h10 ;
			data[70249] <= 8'h10 ;
			data[70250] <= 8'h10 ;
			data[70251] <= 8'h10 ;
			data[70252] <= 8'h10 ;
			data[70253] <= 8'h10 ;
			data[70254] <= 8'h10 ;
			data[70255] <= 8'h10 ;
			data[70256] <= 8'h10 ;
			data[70257] <= 8'h10 ;
			data[70258] <= 8'h10 ;
			data[70259] <= 8'h10 ;
			data[70260] <= 8'h10 ;
			data[70261] <= 8'h10 ;
			data[70262] <= 8'h10 ;
			data[70263] <= 8'h10 ;
			data[70264] <= 8'h10 ;
			data[70265] <= 8'h10 ;
			data[70266] <= 8'h10 ;
			data[70267] <= 8'h10 ;
			data[70268] <= 8'h10 ;
			data[70269] <= 8'h10 ;
			data[70270] <= 8'h10 ;
			data[70271] <= 8'h10 ;
			data[70272] <= 8'h10 ;
			data[70273] <= 8'h10 ;
			data[70274] <= 8'h10 ;
			data[70275] <= 8'h10 ;
			data[70276] <= 8'h10 ;
			data[70277] <= 8'h10 ;
			data[70278] <= 8'h10 ;
			data[70279] <= 8'h10 ;
			data[70280] <= 8'h10 ;
			data[70281] <= 8'h10 ;
			data[70282] <= 8'h10 ;
			data[70283] <= 8'h10 ;
			data[70284] <= 8'h10 ;
			data[70285] <= 8'h10 ;
			data[70286] <= 8'h10 ;
			data[70287] <= 8'h10 ;
			data[70288] <= 8'h10 ;
			data[70289] <= 8'h10 ;
			data[70290] <= 8'h10 ;
			data[70291] <= 8'h10 ;
			data[70292] <= 8'h10 ;
			data[70293] <= 8'h10 ;
			data[70294] <= 8'h10 ;
			data[70295] <= 8'h10 ;
			data[70296] <= 8'h10 ;
			data[70297] <= 8'h10 ;
			data[70298] <= 8'h10 ;
			data[70299] <= 8'h10 ;
			data[70300] <= 8'h10 ;
			data[70301] <= 8'h10 ;
			data[70302] <= 8'h10 ;
			data[70303] <= 8'h10 ;
			data[70304] <= 8'h10 ;
			data[70305] <= 8'h10 ;
			data[70306] <= 8'h10 ;
			data[70307] <= 8'h10 ;
			data[70308] <= 8'h10 ;
			data[70309] <= 8'h10 ;
			data[70310] <= 8'h10 ;
			data[70311] <= 8'h10 ;
			data[70312] <= 8'h10 ;
			data[70313] <= 8'h10 ;
			data[70314] <= 8'h10 ;
			data[70315] <= 8'h10 ;
			data[70316] <= 8'h10 ;
			data[70317] <= 8'h10 ;
			data[70318] <= 8'h10 ;
			data[70319] <= 8'h10 ;
			data[70320] <= 8'h10 ;
			data[70321] <= 8'h10 ;
			data[70322] <= 8'h10 ;
			data[70323] <= 8'h10 ;
			data[70324] <= 8'h10 ;
			data[70325] <= 8'h10 ;
			data[70326] <= 8'h10 ;
			data[70327] <= 8'h10 ;
			data[70328] <= 8'h10 ;
			data[70329] <= 8'h10 ;
			data[70330] <= 8'h10 ;
			data[70331] <= 8'h10 ;
			data[70332] <= 8'h10 ;
			data[70333] <= 8'h10 ;
			data[70334] <= 8'h10 ;
			data[70335] <= 8'h10 ;
			data[70336] <= 8'h10 ;
			data[70337] <= 8'h10 ;
			data[70338] <= 8'h10 ;
			data[70339] <= 8'h10 ;
			data[70340] <= 8'h10 ;
			data[70341] <= 8'h10 ;
			data[70342] <= 8'h10 ;
			data[70343] <= 8'h10 ;
			data[70344] <= 8'h10 ;
			data[70345] <= 8'h10 ;
			data[70346] <= 8'h10 ;
			data[70347] <= 8'h10 ;
			data[70348] <= 8'h10 ;
			data[70349] <= 8'h10 ;
			data[70350] <= 8'h10 ;
			data[70351] <= 8'h10 ;
			data[70352] <= 8'h10 ;
			data[70353] <= 8'h10 ;
			data[70354] <= 8'h10 ;
			data[70355] <= 8'h10 ;
			data[70356] <= 8'h10 ;
			data[70357] <= 8'h10 ;
			data[70358] <= 8'h10 ;
			data[70359] <= 8'h10 ;
			data[70360] <= 8'h10 ;
			data[70361] <= 8'h10 ;
			data[70362] <= 8'h10 ;
			data[70363] <= 8'h10 ;
			data[70364] <= 8'h10 ;
			data[70365] <= 8'h10 ;
			data[70366] <= 8'h10 ;
			data[70367] <= 8'h10 ;
			data[70368] <= 8'h10 ;
			data[70369] <= 8'h10 ;
			data[70370] <= 8'h10 ;
			data[70371] <= 8'h10 ;
			data[70372] <= 8'h10 ;
			data[70373] <= 8'h10 ;
			data[70374] <= 8'h10 ;
			data[70375] <= 8'h10 ;
			data[70376] <= 8'h10 ;
			data[70377] <= 8'h10 ;
			data[70378] <= 8'h10 ;
			data[70379] <= 8'h10 ;
			data[70380] <= 8'h10 ;
			data[70381] <= 8'h10 ;
			data[70382] <= 8'h10 ;
			data[70383] <= 8'h10 ;
			data[70384] <= 8'h10 ;
			data[70385] <= 8'h10 ;
			data[70386] <= 8'h10 ;
			data[70387] <= 8'h10 ;
			data[70388] <= 8'h10 ;
			data[70389] <= 8'h10 ;
			data[70390] <= 8'h10 ;
			data[70391] <= 8'h10 ;
			data[70392] <= 8'h10 ;
			data[70393] <= 8'h10 ;
			data[70394] <= 8'h10 ;
			data[70395] <= 8'h10 ;
			data[70396] <= 8'h10 ;
			data[70397] <= 8'h10 ;
			data[70398] <= 8'h10 ;
			data[70399] <= 8'h10 ;
			data[70400] <= 8'h10 ;
			data[70401] <= 8'h10 ;
			data[70402] <= 8'h10 ;
			data[70403] <= 8'h10 ;
			data[70404] <= 8'h10 ;
			data[70405] <= 8'h10 ;
			data[70406] <= 8'h10 ;
			data[70407] <= 8'h10 ;
			data[70408] <= 8'h10 ;
			data[70409] <= 8'h10 ;
			data[70410] <= 8'h10 ;
			data[70411] <= 8'h10 ;
			data[70412] <= 8'h10 ;
			data[70413] <= 8'h10 ;
			data[70414] <= 8'h10 ;
			data[70415] <= 8'h10 ;
			data[70416] <= 8'h10 ;
			data[70417] <= 8'h10 ;
			data[70418] <= 8'h10 ;
			data[70419] <= 8'h10 ;
			data[70420] <= 8'h10 ;
			data[70421] <= 8'h10 ;
			data[70422] <= 8'h10 ;
			data[70423] <= 8'h10 ;
			data[70424] <= 8'h10 ;
			data[70425] <= 8'h10 ;
			data[70426] <= 8'h10 ;
			data[70427] <= 8'h10 ;
			data[70428] <= 8'h10 ;
			data[70429] <= 8'h10 ;
			data[70430] <= 8'h10 ;
			data[70431] <= 8'h10 ;
			data[70432] <= 8'h10 ;
			data[70433] <= 8'h10 ;
			data[70434] <= 8'h10 ;
			data[70435] <= 8'h10 ;
			data[70436] <= 8'h10 ;
			data[70437] <= 8'h10 ;
			data[70438] <= 8'h10 ;
			data[70439] <= 8'h10 ;
			data[70440] <= 8'h10 ;
			data[70441] <= 8'h10 ;
			data[70442] <= 8'h10 ;
			data[70443] <= 8'h10 ;
			data[70444] <= 8'h10 ;
			data[70445] <= 8'h10 ;
			data[70446] <= 8'h10 ;
			data[70447] <= 8'h10 ;
			data[70448] <= 8'h10 ;
			data[70449] <= 8'h10 ;
			data[70450] <= 8'h10 ;
			data[70451] <= 8'h10 ;
			data[70452] <= 8'h10 ;
			data[70453] <= 8'h10 ;
			data[70454] <= 8'h10 ;
			data[70455] <= 8'h10 ;
			data[70456] <= 8'h10 ;
			data[70457] <= 8'h10 ;
			data[70458] <= 8'h10 ;
			data[70459] <= 8'h10 ;
			data[70460] <= 8'h10 ;
			data[70461] <= 8'h10 ;
			data[70462] <= 8'h10 ;
			data[70463] <= 8'h10 ;
			data[70464] <= 8'h10 ;
			data[70465] <= 8'h10 ;
			data[70466] <= 8'h10 ;
			data[70467] <= 8'h10 ;
			data[70468] <= 8'h10 ;
			data[70469] <= 8'h10 ;
			data[70470] <= 8'h10 ;
			data[70471] <= 8'h10 ;
			data[70472] <= 8'h10 ;
			data[70473] <= 8'h10 ;
			data[70474] <= 8'h10 ;
			data[70475] <= 8'h10 ;
			data[70476] <= 8'h10 ;
			data[70477] <= 8'h10 ;
			data[70478] <= 8'h10 ;
			data[70479] <= 8'h10 ;
			data[70480] <= 8'h10 ;
			data[70481] <= 8'h10 ;
			data[70482] <= 8'h10 ;
			data[70483] <= 8'h10 ;
			data[70484] <= 8'h10 ;
			data[70485] <= 8'h10 ;
			data[70486] <= 8'h10 ;
			data[70487] <= 8'h10 ;
			data[70488] <= 8'h10 ;
			data[70489] <= 8'h10 ;
			data[70490] <= 8'h10 ;
			data[70491] <= 8'h10 ;
			data[70492] <= 8'h10 ;
			data[70493] <= 8'h10 ;
			data[70494] <= 8'h10 ;
			data[70495] <= 8'h10 ;
			data[70496] <= 8'h10 ;
			data[70497] <= 8'h10 ;
			data[70498] <= 8'h10 ;
			data[70499] <= 8'h10 ;
			data[70500] <= 8'h10 ;
			data[70501] <= 8'h10 ;
			data[70502] <= 8'h10 ;
			data[70503] <= 8'h10 ;
			data[70504] <= 8'h10 ;
			data[70505] <= 8'h10 ;
			data[70506] <= 8'h10 ;
			data[70507] <= 8'h10 ;
			data[70508] <= 8'h10 ;
			data[70509] <= 8'h10 ;
			data[70510] <= 8'h10 ;
			data[70511] <= 8'h10 ;
			data[70512] <= 8'h10 ;
			data[70513] <= 8'h10 ;
			data[70514] <= 8'h10 ;
			data[70515] <= 8'h10 ;
			data[70516] <= 8'h10 ;
			data[70517] <= 8'h10 ;
			data[70518] <= 8'h10 ;
			data[70519] <= 8'h10 ;
			data[70520] <= 8'h10 ;
			data[70521] <= 8'h10 ;
			data[70522] <= 8'h10 ;
			data[70523] <= 8'h10 ;
			data[70524] <= 8'h10 ;
			data[70525] <= 8'h10 ;
			data[70526] <= 8'h10 ;
			data[70527] <= 8'h10 ;
			data[70528] <= 8'h10 ;
			data[70529] <= 8'h10 ;
			data[70530] <= 8'h10 ;
			data[70531] <= 8'h10 ;
			data[70532] <= 8'h10 ;
			data[70533] <= 8'h10 ;
			data[70534] <= 8'h10 ;
			data[70535] <= 8'h10 ;
			data[70536] <= 8'h10 ;
			data[70537] <= 8'h10 ;
			data[70538] <= 8'h10 ;
			data[70539] <= 8'h10 ;
			data[70540] <= 8'h10 ;
			data[70541] <= 8'h10 ;
			data[70542] <= 8'h10 ;
			data[70543] <= 8'h10 ;
			data[70544] <= 8'h10 ;
			data[70545] <= 8'h10 ;
			data[70546] <= 8'h10 ;
			data[70547] <= 8'h10 ;
			data[70548] <= 8'h10 ;
			data[70549] <= 8'h10 ;
			data[70550] <= 8'h10 ;
			data[70551] <= 8'h10 ;
			data[70552] <= 8'h10 ;
			data[70553] <= 8'h10 ;
			data[70554] <= 8'h10 ;
			data[70555] <= 8'h10 ;
			data[70556] <= 8'h10 ;
			data[70557] <= 8'h10 ;
			data[70558] <= 8'h10 ;
			data[70559] <= 8'h10 ;
			data[70560] <= 8'h10 ;
			data[70561] <= 8'h10 ;
			data[70562] <= 8'h10 ;
			data[70563] <= 8'h10 ;
			data[70564] <= 8'h10 ;
			data[70565] <= 8'h10 ;
			data[70566] <= 8'h10 ;
			data[70567] <= 8'h10 ;
			data[70568] <= 8'h10 ;
			data[70569] <= 8'h10 ;
			data[70570] <= 8'h10 ;
			data[70571] <= 8'h10 ;
			data[70572] <= 8'h10 ;
			data[70573] <= 8'h10 ;
			data[70574] <= 8'h10 ;
			data[70575] <= 8'h10 ;
			data[70576] <= 8'h10 ;
			data[70577] <= 8'h10 ;
			data[70578] <= 8'h10 ;
			data[70579] <= 8'h10 ;
			data[70580] <= 8'h10 ;
			data[70581] <= 8'h10 ;
			data[70582] <= 8'h10 ;
			data[70583] <= 8'h10 ;
			data[70584] <= 8'h10 ;
			data[70585] <= 8'h10 ;
			data[70586] <= 8'h10 ;
			data[70587] <= 8'h10 ;
			data[70588] <= 8'h10 ;
			data[70589] <= 8'h10 ;
			data[70590] <= 8'h10 ;
			data[70591] <= 8'h10 ;
			data[70592] <= 8'h10 ;
			data[70593] <= 8'h10 ;
			data[70594] <= 8'h10 ;
			data[70595] <= 8'h10 ;
			data[70596] <= 8'h10 ;
			data[70597] <= 8'h10 ;
			data[70598] <= 8'h10 ;
			data[70599] <= 8'h10 ;
			data[70600] <= 8'h10 ;
			data[70601] <= 8'h10 ;
			data[70602] <= 8'h10 ;
			data[70603] <= 8'h10 ;
			data[70604] <= 8'h10 ;
			data[70605] <= 8'h10 ;
			data[70606] <= 8'h10 ;
			data[70607] <= 8'h10 ;
			data[70608] <= 8'h10 ;
			data[70609] <= 8'h10 ;
			data[70610] <= 8'h10 ;
			data[70611] <= 8'h10 ;
			data[70612] <= 8'h10 ;
			data[70613] <= 8'h10 ;
			data[70614] <= 8'h10 ;
			data[70615] <= 8'h10 ;
			data[70616] <= 8'h10 ;
			data[70617] <= 8'h10 ;
			data[70618] <= 8'h10 ;
			data[70619] <= 8'h10 ;
			data[70620] <= 8'h10 ;
			data[70621] <= 8'h10 ;
			data[70622] <= 8'h10 ;
			data[70623] <= 8'h10 ;
			data[70624] <= 8'h10 ;
			data[70625] <= 8'h10 ;
			data[70626] <= 8'h10 ;
			data[70627] <= 8'h10 ;
			data[70628] <= 8'h10 ;
			data[70629] <= 8'h10 ;
			data[70630] <= 8'h10 ;
			data[70631] <= 8'h10 ;
			data[70632] <= 8'h10 ;
			data[70633] <= 8'h10 ;
			data[70634] <= 8'h10 ;
			data[70635] <= 8'h10 ;
			data[70636] <= 8'h10 ;
			data[70637] <= 8'h10 ;
			data[70638] <= 8'h10 ;
			data[70639] <= 8'h10 ;
			data[70640] <= 8'h10 ;
			data[70641] <= 8'h10 ;
			data[70642] <= 8'h10 ;
			data[70643] <= 8'h10 ;
			data[70644] <= 8'h10 ;
			data[70645] <= 8'h10 ;
			data[70646] <= 8'h10 ;
			data[70647] <= 8'h10 ;
			data[70648] <= 8'h10 ;
			data[70649] <= 8'h10 ;
			data[70650] <= 8'h10 ;
			data[70651] <= 8'h10 ;
			data[70652] <= 8'h10 ;
			data[70653] <= 8'h10 ;
			data[70654] <= 8'h10 ;
			data[70655] <= 8'h10 ;
			data[70656] <= 8'h10 ;
			data[70657] <= 8'h10 ;
			data[70658] <= 8'h10 ;
			data[70659] <= 8'h10 ;
			data[70660] <= 8'h10 ;
			data[70661] <= 8'h10 ;
			data[70662] <= 8'h10 ;
			data[70663] <= 8'h10 ;
			data[70664] <= 8'h10 ;
			data[70665] <= 8'h10 ;
			data[70666] <= 8'h10 ;
			data[70667] <= 8'h10 ;
			data[70668] <= 8'h10 ;
			data[70669] <= 8'h10 ;
			data[70670] <= 8'h10 ;
			data[70671] <= 8'h10 ;
			data[70672] <= 8'h10 ;
			data[70673] <= 8'h10 ;
			data[70674] <= 8'h10 ;
			data[70675] <= 8'h10 ;
			data[70676] <= 8'h10 ;
			data[70677] <= 8'h10 ;
			data[70678] <= 8'h10 ;
			data[70679] <= 8'h10 ;
			data[70680] <= 8'h10 ;
			data[70681] <= 8'h10 ;
			data[70682] <= 8'h10 ;
			data[70683] <= 8'h10 ;
			data[70684] <= 8'h10 ;
			data[70685] <= 8'h10 ;
			data[70686] <= 8'h10 ;
			data[70687] <= 8'h10 ;
			data[70688] <= 8'h10 ;
			data[70689] <= 8'h10 ;
			data[70690] <= 8'h10 ;
			data[70691] <= 8'h10 ;
			data[70692] <= 8'h10 ;
			data[70693] <= 8'h10 ;
			data[70694] <= 8'h10 ;
			data[70695] <= 8'h10 ;
			data[70696] <= 8'h10 ;
			data[70697] <= 8'h10 ;
			data[70698] <= 8'h10 ;
			data[70699] <= 8'h10 ;
			data[70700] <= 8'h10 ;
			data[70701] <= 8'h10 ;
			data[70702] <= 8'h10 ;
			data[70703] <= 8'h10 ;
			data[70704] <= 8'h10 ;
			data[70705] <= 8'h10 ;
			data[70706] <= 8'h10 ;
			data[70707] <= 8'h10 ;
			data[70708] <= 8'h10 ;
			data[70709] <= 8'h10 ;
			data[70710] <= 8'h10 ;
			data[70711] <= 8'h10 ;
			data[70712] <= 8'h10 ;
			data[70713] <= 8'h10 ;
			data[70714] <= 8'h10 ;
			data[70715] <= 8'h10 ;
			data[70716] <= 8'h10 ;
			data[70717] <= 8'h10 ;
			data[70718] <= 8'h10 ;
			data[70719] <= 8'h10 ;
			data[70720] <= 8'h10 ;
			data[70721] <= 8'h10 ;
			data[70722] <= 8'h10 ;
			data[70723] <= 8'h10 ;
			data[70724] <= 8'h10 ;
			data[70725] <= 8'h10 ;
			data[70726] <= 8'h10 ;
			data[70727] <= 8'h10 ;
			data[70728] <= 8'h10 ;
			data[70729] <= 8'h10 ;
			data[70730] <= 8'h10 ;
			data[70731] <= 8'h10 ;
			data[70732] <= 8'h10 ;
			data[70733] <= 8'h10 ;
			data[70734] <= 8'h10 ;
			data[70735] <= 8'h10 ;
			data[70736] <= 8'h10 ;
			data[70737] <= 8'h10 ;
			data[70738] <= 8'h10 ;
			data[70739] <= 8'h10 ;
			data[70740] <= 8'h10 ;
			data[70741] <= 8'h10 ;
			data[70742] <= 8'h10 ;
			data[70743] <= 8'h10 ;
			data[70744] <= 8'h10 ;
			data[70745] <= 8'h10 ;
			data[70746] <= 8'h10 ;
			data[70747] <= 8'h10 ;
			data[70748] <= 8'h10 ;
			data[70749] <= 8'h10 ;
			data[70750] <= 8'h10 ;
			data[70751] <= 8'h10 ;
			data[70752] <= 8'h10 ;
			data[70753] <= 8'h10 ;
			data[70754] <= 8'h10 ;
			data[70755] <= 8'h10 ;
			data[70756] <= 8'h10 ;
			data[70757] <= 8'h10 ;
			data[70758] <= 8'h10 ;
			data[70759] <= 8'h10 ;
			data[70760] <= 8'h10 ;
			data[70761] <= 8'h10 ;
			data[70762] <= 8'h10 ;
			data[70763] <= 8'h10 ;
			data[70764] <= 8'h10 ;
			data[70765] <= 8'h10 ;
			data[70766] <= 8'h10 ;
			data[70767] <= 8'h10 ;
			data[70768] <= 8'h10 ;
			data[70769] <= 8'h10 ;
			data[70770] <= 8'h10 ;
			data[70771] <= 8'h10 ;
			data[70772] <= 8'h10 ;
			data[70773] <= 8'h10 ;
			data[70774] <= 8'h10 ;
			data[70775] <= 8'h10 ;
			data[70776] <= 8'h10 ;
			data[70777] <= 8'h10 ;
			data[70778] <= 8'h10 ;
			data[70779] <= 8'h10 ;
			data[70780] <= 8'h10 ;
			data[70781] <= 8'h10 ;
			data[70782] <= 8'h10 ;
			data[70783] <= 8'h10 ;
			data[70784] <= 8'h10 ;
			data[70785] <= 8'h10 ;
			data[70786] <= 8'h10 ;
			data[70787] <= 8'h10 ;
			data[70788] <= 8'h10 ;
			data[70789] <= 8'h10 ;
			data[70790] <= 8'h10 ;
			data[70791] <= 8'h10 ;
			data[70792] <= 8'h10 ;
			data[70793] <= 8'h10 ;
			data[70794] <= 8'h10 ;
			data[70795] <= 8'h10 ;
			data[70796] <= 8'h10 ;
			data[70797] <= 8'h10 ;
			data[70798] <= 8'h10 ;
			data[70799] <= 8'h10 ;
			data[70800] <= 8'h10 ;
			data[70801] <= 8'h10 ;
			data[70802] <= 8'h10 ;
			data[70803] <= 8'h10 ;
			data[70804] <= 8'h10 ;
			data[70805] <= 8'h10 ;
			data[70806] <= 8'h10 ;
			data[70807] <= 8'h10 ;
			data[70808] <= 8'h10 ;
			data[70809] <= 8'h10 ;
			data[70810] <= 8'h10 ;
			data[70811] <= 8'h10 ;
			data[70812] <= 8'h10 ;
			data[70813] <= 8'h10 ;
			data[70814] <= 8'h10 ;
			data[70815] <= 8'h10 ;
			data[70816] <= 8'h10 ;
			data[70817] <= 8'h10 ;
			data[70818] <= 8'h10 ;
			data[70819] <= 8'h10 ;
			data[70820] <= 8'h10 ;
			data[70821] <= 8'h10 ;
			data[70822] <= 8'h10 ;
			data[70823] <= 8'h10 ;
			data[70824] <= 8'h10 ;
			data[70825] <= 8'h10 ;
			data[70826] <= 8'h10 ;
			data[70827] <= 8'h10 ;
			data[70828] <= 8'h10 ;
			data[70829] <= 8'h10 ;
			data[70830] <= 8'h10 ;
			data[70831] <= 8'h10 ;
			data[70832] <= 8'h10 ;
			data[70833] <= 8'h10 ;
			data[70834] <= 8'h10 ;
			data[70835] <= 8'h10 ;
			data[70836] <= 8'h10 ;
			data[70837] <= 8'h10 ;
			data[70838] <= 8'h10 ;
			data[70839] <= 8'h10 ;
			data[70840] <= 8'h10 ;
			data[70841] <= 8'h10 ;
			data[70842] <= 8'h10 ;
			data[70843] <= 8'h10 ;
			data[70844] <= 8'h10 ;
			data[70845] <= 8'h10 ;
			data[70846] <= 8'h10 ;
			data[70847] <= 8'h10 ;
			data[70848] <= 8'h10 ;
			data[70849] <= 8'h10 ;
			data[70850] <= 8'h10 ;
			data[70851] <= 8'h10 ;
			data[70852] <= 8'h10 ;
			data[70853] <= 8'h10 ;
			data[70854] <= 8'h10 ;
			data[70855] <= 8'h10 ;
			data[70856] <= 8'h10 ;
			data[70857] <= 8'h10 ;
			data[70858] <= 8'h10 ;
			data[70859] <= 8'h10 ;
			data[70860] <= 8'h10 ;
			data[70861] <= 8'h10 ;
			data[70862] <= 8'h10 ;
			data[70863] <= 8'h10 ;
			data[70864] <= 8'h10 ;
			data[70865] <= 8'h10 ;
			data[70866] <= 8'h10 ;
			data[70867] <= 8'h10 ;
			data[70868] <= 8'h10 ;
			data[70869] <= 8'h10 ;
			data[70870] <= 8'h10 ;
			data[70871] <= 8'h10 ;
			data[70872] <= 8'h10 ;
			data[70873] <= 8'h10 ;
			data[70874] <= 8'h10 ;
			data[70875] <= 8'h10 ;
			data[70876] <= 8'h10 ;
			data[70877] <= 8'h10 ;
			data[70878] <= 8'h10 ;
			data[70879] <= 8'h10 ;
			data[70880] <= 8'h10 ;
			data[70881] <= 8'h10 ;
			data[70882] <= 8'h10 ;
			data[70883] <= 8'h10 ;
			data[70884] <= 8'h10 ;
			data[70885] <= 8'h10 ;
			data[70886] <= 8'h10 ;
			data[70887] <= 8'h10 ;
			data[70888] <= 8'h10 ;
			data[70889] <= 8'h10 ;
			data[70890] <= 8'h10 ;
			data[70891] <= 8'h10 ;
			data[70892] <= 8'h10 ;
			data[70893] <= 8'h10 ;
			data[70894] <= 8'h10 ;
			data[70895] <= 8'h10 ;
			data[70896] <= 8'h10 ;
			data[70897] <= 8'h10 ;
			data[70898] <= 8'h10 ;
			data[70899] <= 8'h10 ;
			data[70900] <= 8'h10 ;
			data[70901] <= 8'h10 ;
			data[70902] <= 8'h10 ;
			data[70903] <= 8'h10 ;
			data[70904] <= 8'h10 ;
			data[70905] <= 8'h10 ;
			data[70906] <= 8'h10 ;
			data[70907] <= 8'h10 ;
			data[70908] <= 8'h10 ;
			data[70909] <= 8'h10 ;
			data[70910] <= 8'h10 ;
			data[70911] <= 8'h10 ;
			data[70912] <= 8'h10 ;
			data[70913] <= 8'h10 ;
			data[70914] <= 8'h10 ;
			data[70915] <= 8'h10 ;
			data[70916] <= 8'h10 ;
			data[70917] <= 8'h10 ;
			data[70918] <= 8'h10 ;
			data[70919] <= 8'h10 ;
			data[70920] <= 8'h10 ;
			data[70921] <= 8'h10 ;
			data[70922] <= 8'h10 ;
			data[70923] <= 8'h10 ;
			data[70924] <= 8'h10 ;
			data[70925] <= 8'h10 ;
			data[70926] <= 8'h10 ;
			data[70927] <= 8'h10 ;
			data[70928] <= 8'h10 ;
			data[70929] <= 8'h10 ;
			data[70930] <= 8'h10 ;
			data[70931] <= 8'h10 ;
			data[70932] <= 8'h10 ;
			data[70933] <= 8'h10 ;
			data[70934] <= 8'h10 ;
			data[70935] <= 8'h10 ;
			data[70936] <= 8'h10 ;
			data[70937] <= 8'h10 ;
			data[70938] <= 8'h10 ;
			data[70939] <= 8'h10 ;
			data[70940] <= 8'h10 ;
			data[70941] <= 8'h10 ;
			data[70942] <= 8'h10 ;
			data[70943] <= 8'h10 ;
			data[70944] <= 8'h10 ;
			data[70945] <= 8'h10 ;
			data[70946] <= 8'h10 ;
			data[70947] <= 8'h10 ;
			data[70948] <= 8'h10 ;
			data[70949] <= 8'h10 ;
			data[70950] <= 8'h10 ;
			data[70951] <= 8'h10 ;
			data[70952] <= 8'h10 ;
			data[70953] <= 8'h10 ;
			data[70954] <= 8'h10 ;
			data[70955] <= 8'h10 ;
			data[70956] <= 8'h10 ;
			data[70957] <= 8'h10 ;
			data[70958] <= 8'h10 ;
			data[70959] <= 8'h10 ;
			data[70960] <= 8'h10 ;
			data[70961] <= 8'h10 ;
			data[70962] <= 8'h10 ;
			data[70963] <= 8'h10 ;
			data[70964] <= 8'h10 ;
			data[70965] <= 8'h10 ;
			data[70966] <= 8'h10 ;
			data[70967] <= 8'h10 ;
			data[70968] <= 8'h10 ;
			data[70969] <= 8'h10 ;
			data[70970] <= 8'h10 ;
			data[70971] <= 8'h10 ;
			data[70972] <= 8'h10 ;
			data[70973] <= 8'h10 ;
			data[70974] <= 8'h10 ;
			data[70975] <= 8'h10 ;
			data[70976] <= 8'h10 ;
			data[70977] <= 8'h10 ;
			data[70978] <= 8'h10 ;
			data[70979] <= 8'h10 ;
			data[70980] <= 8'h10 ;
			data[70981] <= 8'h10 ;
			data[70982] <= 8'h10 ;
			data[70983] <= 8'h10 ;
			data[70984] <= 8'h10 ;
			data[70985] <= 8'h10 ;
			data[70986] <= 8'h10 ;
			data[70987] <= 8'h10 ;
			data[70988] <= 8'h10 ;
			data[70989] <= 8'h10 ;
			data[70990] <= 8'h10 ;
			data[70991] <= 8'h10 ;
			data[70992] <= 8'h10 ;
			data[70993] <= 8'h10 ;
			data[70994] <= 8'h10 ;
			data[70995] <= 8'h10 ;
			data[70996] <= 8'h10 ;
			data[70997] <= 8'h10 ;
			data[70998] <= 8'h10 ;
			data[70999] <= 8'h10 ;
			data[71000] <= 8'h10 ;
			data[71001] <= 8'h10 ;
			data[71002] <= 8'h10 ;
			data[71003] <= 8'h10 ;
			data[71004] <= 8'h10 ;
			data[71005] <= 8'h10 ;
			data[71006] <= 8'h10 ;
			data[71007] <= 8'h10 ;
			data[71008] <= 8'h10 ;
			data[71009] <= 8'h10 ;
			data[71010] <= 8'h10 ;
			data[71011] <= 8'h10 ;
			data[71012] <= 8'h10 ;
			data[71013] <= 8'h10 ;
			data[71014] <= 8'h10 ;
			data[71015] <= 8'h10 ;
			data[71016] <= 8'h10 ;
			data[71017] <= 8'h10 ;
			data[71018] <= 8'h10 ;
			data[71019] <= 8'h10 ;
			data[71020] <= 8'h10 ;
			data[71021] <= 8'h10 ;
			data[71022] <= 8'h10 ;
			data[71023] <= 8'h10 ;
			data[71024] <= 8'h10 ;
			data[71025] <= 8'h10 ;
			data[71026] <= 8'h10 ;
			data[71027] <= 8'h10 ;
			data[71028] <= 8'h10 ;
			data[71029] <= 8'h10 ;
			data[71030] <= 8'h10 ;
			data[71031] <= 8'h10 ;
			data[71032] <= 8'h10 ;
			data[71033] <= 8'h10 ;
			data[71034] <= 8'h10 ;
			data[71035] <= 8'h10 ;
			data[71036] <= 8'h10 ;
			data[71037] <= 8'h10 ;
			data[71038] <= 8'h10 ;
			data[71039] <= 8'h10 ;
			data[71040] <= 8'h10 ;
			data[71041] <= 8'h10 ;
			data[71042] <= 8'h10 ;
			data[71043] <= 8'h10 ;
			data[71044] <= 8'h10 ;
			data[71045] <= 8'h10 ;
			data[71046] <= 8'h10 ;
			data[71047] <= 8'h10 ;
			data[71048] <= 8'h10 ;
			data[71049] <= 8'h10 ;
			data[71050] <= 8'h10 ;
			data[71051] <= 8'h10 ;
			data[71052] <= 8'h10 ;
			data[71053] <= 8'h10 ;
			data[71054] <= 8'h10 ;
			data[71055] <= 8'h10 ;
			data[71056] <= 8'h10 ;
			data[71057] <= 8'h10 ;
			data[71058] <= 8'h10 ;
			data[71059] <= 8'h10 ;
			data[71060] <= 8'h10 ;
			data[71061] <= 8'h10 ;
			data[71062] <= 8'h10 ;
			data[71063] <= 8'h10 ;
			data[71064] <= 8'h10 ;
			data[71065] <= 8'h10 ;
			data[71066] <= 8'h10 ;
			data[71067] <= 8'h10 ;
			data[71068] <= 8'h10 ;
			data[71069] <= 8'h10 ;
			data[71070] <= 8'h10 ;
			data[71071] <= 8'h10 ;
			data[71072] <= 8'h10 ;
			data[71073] <= 8'h10 ;
			data[71074] <= 8'h10 ;
			data[71075] <= 8'h10 ;
			data[71076] <= 8'h10 ;
			data[71077] <= 8'h10 ;
			data[71078] <= 8'h10 ;
			data[71079] <= 8'h10 ;
			data[71080] <= 8'h10 ;
			data[71081] <= 8'h10 ;
			data[71082] <= 8'h10 ;
			data[71083] <= 8'h10 ;
			data[71084] <= 8'h10 ;
			data[71085] <= 8'h10 ;
			data[71086] <= 8'h10 ;
			data[71087] <= 8'h10 ;
			data[71088] <= 8'h10 ;
			data[71089] <= 8'h10 ;
			data[71090] <= 8'h10 ;
			data[71091] <= 8'h10 ;
			data[71092] <= 8'h10 ;
			data[71093] <= 8'h10 ;
			data[71094] <= 8'h10 ;
			data[71095] <= 8'h10 ;
			data[71096] <= 8'h10 ;
			data[71097] <= 8'h10 ;
			data[71098] <= 8'h10 ;
			data[71099] <= 8'h10 ;
			data[71100] <= 8'h10 ;
			data[71101] <= 8'h10 ;
			data[71102] <= 8'h10 ;
			data[71103] <= 8'h10 ;
			data[71104] <= 8'h10 ;
			data[71105] <= 8'h10 ;
			data[71106] <= 8'h10 ;
			data[71107] <= 8'h10 ;
			data[71108] <= 8'h10 ;
			data[71109] <= 8'h10 ;
			data[71110] <= 8'h10 ;
			data[71111] <= 8'h10 ;
			data[71112] <= 8'h10 ;
			data[71113] <= 8'h10 ;
			data[71114] <= 8'h10 ;
			data[71115] <= 8'h10 ;
			data[71116] <= 8'h10 ;
			data[71117] <= 8'h10 ;
			data[71118] <= 8'h10 ;
			data[71119] <= 8'h10 ;
			data[71120] <= 8'h10 ;
			data[71121] <= 8'h10 ;
			data[71122] <= 8'h10 ;
			data[71123] <= 8'h10 ;
			data[71124] <= 8'h10 ;
			data[71125] <= 8'h10 ;
			data[71126] <= 8'h10 ;
			data[71127] <= 8'h10 ;
			data[71128] <= 8'h10 ;
			data[71129] <= 8'h10 ;
			data[71130] <= 8'h10 ;
			data[71131] <= 8'h10 ;
			data[71132] <= 8'h10 ;
			data[71133] <= 8'h10 ;
			data[71134] <= 8'h10 ;
			data[71135] <= 8'h10 ;
			data[71136] <= 8'h10 ;
			data[71137] <= 8'h10 ;
			data[71138] <= 8'h10 ;
			data[71139] <= 8'h10 ;
			data[71140] <= 8'h10 ;
			data[71141] <= 8'h10 ;
			data[71142] <= 8'h10 ;
			data[71143] <= 8'h10 ;
			data[71144] <= 8'h10 ;
			data[71145] <= 8'h10 ;
			data[71146] <= 8'h10 ;
			data[71147] <= 8'h10 ;
			data[71148] <= 8'h10 ;
			data[71149] <= 8'h10 ;
			data[71150] <= 8'h10 ;
			data[71151] <= 8'h10 ;
			data[71152] <= 8'h10 ;
			data[71153] <= 8'h10 ;
			data[71154] <= 8'h10 ;
			data[71155] <= 8'h10 ;
			data[71156] <= 8'h10 ;
			data[71157] <= 8'h10 ;
			data[71158] <= 8'h10 ;
			data[71159] <= 8'h10 ;
			data[71160] <= 8'h10 ;
			data[71161] <= 8'h10 ;
			data[71162] <= 8'h10 ;
			data[71163] <= 8'h10 ;
			data[71164] <= 8'h10 ;
			data[71165] <= 8'h10 ;
			data[71166] <= 8'h10 ;
			data[71167] <= 8'h10 ;
			data[71168] <= 8'h10 ;
			data[71169] <= 8'h10 ;
			data[71170] <= 8'h10 ;
			data[71171] <= 8'h10 ;
			data[71172] <= 8'h10 ;
			data[71173] <= 8'h10 ;
			data[71174] <= 8'h10 ;
			data[71175] <= 8'h10 ;
			data[71176] <= 8'h10 ;
			data[71177] <= 8'h10 ;
			data[71178] <= 8'h10 ;
			data[71179] <= 8'h10 ;
			data[71180] <= 8'h10 ;
			data[71181] <= 8'h10 ;
			data[71182] <= 8'h10 ;
			data[71183] <= 8'h10 ;
			data[71184] <= 8'h10 ;
			data[71185] <= 8'h10 ;
			data[71186] <= 8'h10 ;
			data[71187] <= 8'h10 ;
			data[71188] <= 8'h10 ;
			data[71189] <= 8'h10 ;
			data[71190] <= 8'h10 ;
			data[71191] <= 8'h10 ;
			data[71192] <= 8'h10 ;
			data[71193] <= 8'h10 ;
			data[71194] <= 8'h10 ;
			data[71195] <= 8'h10 ;
			data[71196] <= 8'h10 ;
			data[71197] <= 8'h10 ;
			data[71198] <= 8'h10 ;
			data[71199] <= 8'h10 ;
			data[71200] <= 8'h10 ;
			data[71201] <= 8'h10 ;
			data[71202] <= 8'h10 ;
			data[71203] <= 8'h10 ;
			data[71204] <= 8'h10 ;
			data[71205] <= 8'h10 ;
			data[71206] <= 8'h10 ;
			data[71207] <= 8'h10 ;
			data[71208] <= 8'h10 ;
			data[71209] <= 8'h10 ;
			data[71210] <= 8'h10 ;
			data[71211] <= 8'h10 ;
			data[71212] <= 8'h10 ;
			data[71213] <= 8'h10 ;
			data[71214] <= 8'h10 ;
			data[71215] <= 8'h10 ;
			data[71216] <= 8'h10 ;
			data[71217] <= 8'h10 ;
			data[71218] <= 8'h10 ;
			data[71219] <= 8'h10 ;
			data[71220] <= 8'h10 ;
			data[71221] <= 8'h10 ;
			data[71222] <= 8'h10 ;
			data[71223] <= 8'h10 ;
			data[71224] <= 8'h10 ;
			data[71225] <= 8'h10 ;
			data[71226] <= 8'h10 ;
			data[71227] <= 8'h10 ;
			data[71228] <= 8'h10 ;
			data[71229] <= 8'h10 ;
			data[71230] <= 8'h10 ;
			data[71231] <= 8'h10 ;
			data[71232] <= 8'h10 ;
			data[71233] <= 8'h10 ;
			data[71234] <= 8'h10 ;
			data[71235] <= 8'h10 ;
			data[71236] <= 8'h10 ;
			data[71237] <= 8'h10 ;
			data[71238] <= 8'h10 ;
			data[71239] <= 8'h10 ;
			data[71240] <= 8'h10 ;
			data[71241] <= 8'h10 ;
			data[71242] <= 8'h10 ;
			data[71243] <= 8'h10 ;
			data[71244] <= 8'h10 ;
			data[71245] <= 8'h10 ;
			data[71246] <= 8'h10 ;
			data[71247] <= 8'h10 ;
			data[71248] <= 8'h10 ;
			data[71249] <= 8'h10 ;
			data[71250] <= 8'h10 ;
			data[71251] <= 8'h10 ;
			data[71252] <= 8'h10 ;
			data[71253] <= 8'h10 ;
			data[71254] <= 8'h10 ;
			data[71255] <= 8'h10 ;
			data[71256] <= 8'h10 ;
			data[71257] <= 8'h10 ;
			data[71258] <= 8'h10 ;
			data[71259] <= 8'h10 ;
			data[71260] <= 8'h10 ;
			data[71261] <= 8'h10 ;
			data[71262] <= 8'h10 ;
			data[71263] <= 8'h10 ;
			data[71264] <= 8'h10 ;
			data[71265] <= 8'h10 ;
			data[71266] <= 8'h10 ;
			data[71267] <= 8'h10 ;
			data[71268] <= 8'h10 ;
			data[71269] <= 8'h10 ;
			data[71270] <= 8'h10 ;
			data[71271] <= 8'h10 ;
			data[71272] <= 8'h10 ;
			data[71273] <= 8'h10 ;
			data[71274] <= 8'h10 ;
			data[71275] <= 8'h10 ;
			data[71276] <= 8'h10 ;
			data[71277] <= 8'h10 ;
			data[71278] <= 8'h10 ;
			data[71279] <= 8'h10 ;
			data[71280] <= 8'h10 ;
			data[71281] <= 8'h10 ;
			data[71282] <= 8'h10 ;
			data[71283] <= 8'h10 ;
			data[71284] <= 8'h10 ;
			data[71285] <= 8'h10 ;
			data[71286] <= 8'h10 ;
			data[71287] <= 8'h10 ;
			data[71288] <= 8'h10 ;
			data[71289] <= 8'h10 ;
			data[71290] <= 8'h10 ;
			data[71291] <= 8'h10 ;
			data[71292] <= 8'h10 ;
			data[71293] <= 8'h10 ;
			data[71294] <= 8'h10 ;
			data[71295] <= 8'h10 ;
			data[71296] <= 8'h10 ;
			data[71297] <= 8'h10 ;
			data[71298] <= 8'h10 ;
			data[71299] <= 8'h10 ;
			data[71300] <= 8'h10 ;
			data[71301] <= 8'h10 ;
			data[71302] <= 8'h10 ;
			data[71303] <= 8'h10 ;
			data[71304] <= 8'h10 ;
			data[71305] <= 8'h10 ;
			data[71306] <= 8'h10 ;
			data[71307] <= 8'h10 ;
			data[71308] <= 8'h10 ;
			data[71309] <= 8'h10 ;
			data[71310] <= 8'h10 ;
			data[71311] <= 8'h10 ;
			data[71312] <= 8'h10 ;
			data[71313] <= 8'h10 ;
			data[71314] <= 8'h10 ;
			data[71315] <= 8'h10 ;
			data[71316] <= 8'h10 ;
			data[71317] <= 8'h10 ;
			data[71318] <= 8'h10 ;
			data[71319] <= 8'h10 ;
			data[71320] <= 8'h10 ;
			data[71321] <= 8'h10 ;
			data[71322] <= 8'h10 ;
			data[71323] <= 8'h10 ;
			data[71324] <= 8'h10 ;
			data[71325] <= 8'h10 ;
			data[71326] <= 8'h10 ;
			data[71327] <= 8'h10 ;
			data[71328] <= 8'h10 ;
			data[71329] <= 8'h10 ;
			data[71330] <= 8'h10 ;
			data[71331] <= 8'h10 ;
			data[71332] <= 8'h10 ;
			data[71333] <= 8'h10 ;
			data[71334] <= 8'h10 ;
			data[71335] <= 8'h10 ;
			data[71336] <= 8'h10 ;
			data[71337] <= 8'h10 ;
			data[71338] <= 8'h10 ;
			data[71339] <= 8'h10 ;
			data[71340] <= 8'h10 ;
			data[71341] <= 8'h10 ;
			data[71342] <= 8'h10 ;
			data[71343] <= 8'h10 ;
			data[71344] <= 8'h10 ;
			data[71345] <= 8'h10 ;
			data[71346] <= 8'h10 ;
			data[71347] <= 8'h10 ;
			data[71348] <= 8'h10 ;
			data[71349] <= 8'h10 ;
			data[71350] <= 8'h10 ;
			data[71351] <= 8'h10 ;
			data[71352] <= 8'h10 ;
			data[71353] <= 8'h10 ;
			data[71354] <= 8'h10 ;
			data[71355] <= 8'h10 ;
			data[71356] <= 8'h10 ;
			data[71357] <= 8'h10 ;
			data[71358] <= 8'h10 ;
			data[71359] <= 8'h10 ;
			data[71360] <= 8'h10 ;
			data[71361] <= 8'h10 ;
			data[71362] <= 8'h10 ;
			data[71363] <= 8'h10 ;
			data[71364] <= 8'h10 ;
			data[71365] <= 8'h10 ;
			data[71366] <= 8'h10 ;
			data[71367] <= 8'h10 ;
			data[71368] <= 8'h10 ;
			data[71369] <= 8'h10 ;
			data[71370] <= 8'h10 ;
			data[71371] <= 8'h10 ;
			data[71372] <= 8'h10 ;
			data[71373] <= 8'h10 ;
			data[71374] <= 8'h10 ;
			data[71375] <= 8'h10 ;
			data[71376] <= 8'h10 ;
			data[71377] <= 8'h10 ;
			data[71378] <= 8'h10 ;
			data[71379] <= 8'h10 ;
			data[71380] <= 8'h10 ;
			data[71381] <= 8'h10 ;
			data[71382] <= 8'h10 ;
			data[71383] <= 8'h10 ;
			data[71384] <= 8'h10 ;
			data[71385] <= 8'h10 ;
			data[71386] <= 8'h10 ;
			data[71387] <= 8'h10 ;
			data[71388] <= 8'h10 ;
			data[71389] <= 8'h10 ;
			data[71390] <= 8'h10 ;
			data[71391] <= 8'h10 ;
			data[71392] <= 8'h10 ;
			data[71393] <= 8'h10 ;
			data[71394] <= 8'h10 ;
			data[71395] <= 8'h10 ;
			data[71396] <= 8'h10 ;
			data[71397] <= 8'h10 ;
			data[71398] <= 8'h10 ;
			data[71399] <= 8'h10 ;
			data[71400] <= 8'h10 ;
			data[71401] <= 8'h10 ;
			data[71402] <= 8'h10 ;
			data[71403] <= 8'h10 ;
			data[71404] <= 8'h10 ;
			data[71405] <= 8'h10 ;
			data[71406] <= 8'h10 ;
			data[71407] <= 8'h10 ;
			data[71408] <= 8'h10 ;
			data[71409] <= 8'h10 ;
			data[71410] <= 8'h10 ;
			data[71411] <= 8'h10 ;
			data[71412] <= 8'h10 ;
			data[71413] <= 8'h10 ;
			data[71414] <= 8'h10 ;
			data[71415] <= 8'h10 ;
			data[71416] <= 8'h10 ;
			data[71417] <= 8'h10 ;
			data[71418] <= 8'h10 ;
			data[71419] <= 8'h10 ;
			data[71420] <= 8'h10 ;
			data[71421] <= 8'h10 ;
			data[71422] <= 8'h10 ;
			data[71423] <= 8'h10 ;
			data[71424] <= 8'h10 ;
			data[71425] <= 8'h10 ;
			data[71426] <= 8'h10 ;
			data[71427] <= 8'h10 ;
			data[71428] <= 8'h10 ;
			data[71429] <= 8'h10 ;
			data[71430] <= 8'h10 ;
			data[71431] <= 8'h10 ;
			data[71432] <= 8'h10 ;
			data[71433] <= 8'h10 ;
			data[71434] <= 8'h10 ;
			data[71435] <= 8'h10 ;
			data[71436] <= 8'h10 ;
			data[71437] <= 8'h10 ;
			data[71438] <= 8'h10 ;
			data[71439] <= 8'h10 ;
			data[71440] <= 8'h10 ;
			data[71441] <= 8'h10 ;
			data[71442] <= 8'h10 ;
			data[71443] <= 8'h10 ;
			data[71444] <= 8'h10 ;
			data[71445] <= 8'h10 ;
			data[71446] <= 8'h10 ;
			data[71447] <= 8'h10 ;
			data[71448] <= 8'h10 ;
			data[71449] <= 8'h10 ;
			data[71450] <= 8'h10 ;
			data[71451] <= 8'h10 ;
			data[71452] <= 8'h10 ;
			data[71453] <= 8'h10 ;
			data[71454] <= 8'h10 ;
			data[71455] <= 8'h10 ;
			data[71456] <= 8'h10 ;
			data[71457] <= 8'h10 ;
			data[71458] <= 8'h10 ;
			data[71459] <= 8'h10 ;
			data[71460] <= 8'h10 ;
			data[71461] <= 8'h10 ;
			data[71462] <= 8'h10 ;
			data[71463] <= 8'h10 ;
			data[71464] <= 8'h10 ;
			data[71465] <= 8'h10 ;
			data[71466] <= 8'h10 ;
			data[71467] <= 8'h10 ;
			data[71468] <= 8'h10 ;
			data[71469] <= 8'h10 ;
			data[71470] <= 8'h10 ;
			data[71471] <= 8'h10 ;
			data[71472] <= 8'h10 ;
			data[71473] <= 8'h10 ;
			data[71474] <= 8'h10 ;
			data[71475] <= 8'h10 ;
			data[71476] <= 8'h10 ;
			data[71477] <= 8'h10 ;
			data[71478] <= 8'h10 ;
			data[71479] <= 8'h10 ;
			data[71480] <= 8'h10 ;
			data[71481] <= 8'h10 ;
			data[71482] <= 8'h10 ;
			data[71483] <= 8'h10 ;
			data[71484] <= 8'h10 ;
			data[71485] <= 8'h10 ;
			data[71486] <= 8'h10 ;
			data[71487] <= 8'h10 ;
			data[71488] <= 8'h10 ;
			data[71489] <= 8'h10 ;
			data[71490] <= 8'h10 ;
			data[71491] <= 8'h10 ;
			data[71492] <= 8'h10 ;
			data[71493] <= 8'h10 ;
			data[71494] <= 8'h10 ;
			data[71495] <= 8'h10 ;
			data[71496] <= 8'h10 ;
			data[71497] <= 8'h10 ;
			data[71498] <= 8'h10 ;
			data[71499] <= 8'h10 ;
			data[71500] <= 8'h10 ;
			data[71501] <= 8'h10 ;
			data[71502] <= 8'h10 ;
			data[71503] <= 8'h10 ;
			data[71504] <= 8'h10 ;
			data[71505] <= 8'h10 ;
			data[71506] <= 8'h10 ;
			data[71507] <= 8'h10 ;
			data[71508] <= 8'h10 ;
			data[71509] <= 8'h10 ;
			data[71510] <= 8'h10 ;
			data[71511] <= 8'h10 ;
			data[71512] <= 8'h10 ;
			data[71513] <= 8'h10 ;
			data[71514] <= 8'h10 ;
			data[71515] <= 8'h10 ;
			data[71516] <= 8'h10 ;
			data[71517] <= 8'h10 ;
			data[71518] <= 8'h10 ;
			data[71519] <= 8'h10 ;
			data[71520] <= 8'h10 ;
			data[71521] <= 8'h10 ;
			data[71522] <= 8'h10 ;
			data[71523] <= 8'h10 ;
			data[71524] <= 8'h10 ;
			data[71525] <= 8'h10 ;
			data[71526] <= 8'h10 ;
			data[71527] <= 8'h10 ;
			data[71528] <= 8'h10 ;
			data[71529] <= 8'h10 ;
			data[71530] <= 8'h10 ;
			data[71531] <= 8'h10 ;
			data[71532] <= 8'h10 ;
			data[71533] <= 8'h10 ;
			data[71534] <= 8'h10 ;
			data[71535] <= 8'h10 ;
			data[71536] <= 8'h10 ;
			data[71537] <= 8'h10 ;
			data[71538] <= 8'h10 ;
			data[71539] <= 8'h10 ;
			data[71540] <= 8'h10 ;
			data[71541] <= 8'h10 ;
			data[71542] <= 8'h10 ;
			data[71543] <= 8'h10 ;
			data[71544] <= 8'h10 ;
			data[71545] <= 8'h10 ;
			data[71546] <= 8'h10 ;
			data[71547] <= 8'h10 ;
			data[71548] <= 8'h10 ;
			data[71549] <= 8'h10 ;
			data[71550] <= 8'h10 ;
			data[71551] <= 8'h10 ;
			data[71552] <= 8'h10 ;
			data[71553] <= 8'h10 ;
			data[71554] <= 8'h10 ;
			data[71555] <= 8'h10 ;
			data[71556] <= 8'h10 ;
			data[71557] <= 8'h10 ;
			data[71558] <= 8'h10 ;
			data[71559] <= 8'h10 ;
			data[71560] <= 8'h10 ;
			data[71561] <= 8'h10 ;
			data[71562] <= 8'h10 ;
			data[71563] <= 8'h10 ;
			data[71564] <= 8'h10 ;
			data[71565] <= 8'h10 ;
			data[71566] <= 8'h10 ;
			data[71567] <= 8'h10 ;
			data[71568] <= 8'h10 ;
			data[71569] <= 8'h10 ;
			data[71570] <= 8'h10 ;
			data[71571] <= 8'h10 ;
			data[71572] <= 8'h10 ;
			data[71573] <= 8'h10 ;
			data[71574] <= 8'h10 ;
			data[71575] <= 8'h10 ;
			data[71576] <= 8'h10 ;
			data[71577] <= 8'h10 ;
			data[71578] <= 8'h10 ;
			data[71579] <= 8'h10 ;
			data[71580] <= 8'h10 ;
			data[71581] <= 8'h10 ;
			data[71582] <= 8'h10 ;
			data[71583] <= 8'h10 ;
			data[71584] <= 8'h10 ;
			data[71585] <= 8'h10 ;
			data[71586] <= 8'h10 ;
			data[71587] <= 8'h10 ;
			data[71588] <= 8'h10 ;
			data[71589] <= 8'h10 ;
			data[71590] <= 8'h10 ;
			data[71591] <= 8'h10 ;
			data[71592] <= 8'h10 ;
			data[71593] <= 8'h10 ;
			data[71594] <= 8'h10 ;
			data[71595] <= 8'h10 ;
			data[71596] <= 8'h10 ;
			data[71597] <= 8'h10 ;
			data[71598] <= 8'h10 ;
			data[71599] <= 8'h10 ;
			data[71600] <= 8'h10 ;
			data[71601] <= 8'h10 ;
			data[71602] <= 8'h10 ;
			data[71603] <= 8'h10 ;
			data[71604] <= 8'h10 ;
			data[71605] <= 8'h10 ;
			data[71606] <= 8'h10 ;
			data[71607] <= 8'h10 ;
			data[71608] <= 8'h10 ;
			data[71609] <= 8'h10 ;
			data[71610] <= 8'h10 ;
			data[71611] <= 8'h10 ;
			data[71612] <= 8'h10 ;
			data[71613] <= 8'h10 ;
			data[71614] <= 8'h10 ;
			data[71615] <= 8'h10 ;
			data[71616] <= 8'h10 ;
			data[71617] <= 8'h10 ;
			data[71618] <= 8'h10 ;
			data[71619] <= 8'h10 ;
			data[71620] <= 8'h10 ;
			data[71621] <= 8'h10 ;
			data[71622] <= 8'h10 ;
			data[71623] <= 8'h10 ;
			data[71624] <= 8'h10 ;
			data[71625] <= 8'h10 ;
			data[71626] <= 8'h10 ;
			data[71627] <= 8'h10 ;
			data[71628] <= 8'h10 ;
			data[71629] <= 8'h10 ;
			data[71630] <= 8'h10 ;
			data[71631] <= 8'h10 ;
			data[71632] <= 8'h10 ;
			data[71633] <= 8'h10 ;
			data[71634] <= 8'h10 ;
			data[71635] <= 8'h10 ;
			data[71636] <= 8'h10 ;
			data[71637] <= 8'h10 ;
			data[71638] <= 8'h10 ;
			data[71639] <= 8'h10 ;
			data[71640] <= 8'h10 ;
			data[71641] <= 8'h10 ;
			data[71642] <= 8'h10 ;
			data[71643] <= 8'h10 ;
			data[71644] <= 8'h10 ;
			data[71645] <= 8'h10 ;
			data[71646] <= 8'h10 ;
			data[71647] <= 8'h10 ;
			data[71648] <= 8'h10 ;
			data[71649] <= 8'h10 ;
			data[71650] <= 8'h10 ;
			data[71651] <= 8'h10 ;
			data[71652] <= 8'h10 ;
			data[71653] <= 8'h10 ;
			data[71654] <= 8'h10 ;
			data[71655] <= 8'h10 ;
			data[71656] <= 8'h10 ;
			data[71657] <= 8'h10 ;
			data[71658] <= 8'h10 ;
			data[71659] <= 8'h10 ;
			data[71660] <= 8'h10 ;
			data[71661] <= 8'h10 ;
			data[71662] <= 8'h10 ;
			data[71663] <= 8'h10 ;
			data[71664] <= 8'h10 ;
			data[71665] <= 8'h10 ;
			data[71666] <= 8'h10 ;
			data[71667] <= 8'h10 ;
			data[71668] <= 8'h10 ;
			data[71669] <= 8'h10 ;
			data[71670] <= 8'h10 ;
			data[71671] <= 8'h10 ;
			data[71672] <= 8'h10 ;
			data[71673] <= 8'h10 ;
			data[71674] <= 8'h10 ;
			data[71675] <= 8'h10 ;
			data[71676] <= 8'h10 ;
			data[71677] <= 8'h10 ;
			data[71678] <= 8'h10 ;
			data[71679] <= 8'h10 ;
			data[71680] <= 8'h10 ;
			data[71681] <= 8'h10 ;
			data[71682] <= 8'h10 ;
			data[71683] <= 8'h10 ;
			data[71684] <= 8'h10 ;
			data[71685] <= 8'h10 ;
			data[71686] <= 8'h10 ;
			data[71687] <= 8'h10 ;
			data[71688] <= 8'h10 ;
			data[71689] <= 8'h10 ;
			data[71690] <= 8'h10 ;
			data[71691] <= 8'h10 ;
			data[71692] <= 8'h10 ;
			data[71693] <= 8'h10 ;
			data[71694] <= 8'h10 ;
			data[71695] <= 8'h10 ;
			data[71696] <= 8'h10 ;
			data[71697] <= 8'h10 ;
			data[71698] <= 8'h10 ;
			data[71699] <= 8'h10 ;
			data[71700] <= 8'h10 ;
			data[71701] <= 8'h10 ;
			data[71702] <= 8'h10 ;
			data[71703] <= 8'h10 ;
			data[71704] <= 8'h10 ;
			data[71705] <= 8'h10 ;
			data[71706] <= 8'h10 ;
			data[71707] <= 8'h10 ;
			data[71708] <= 8'h10 ;
			data[71709] <= 8'h10 ;
			data[71710] <= 8'h10 ;
			data[71711] <= 8'h10 ;
			data[71712] <= 8'h10 ;
			data[71713] <= 8'h10 ;
			data[71714] <= 8'h10 ;
			data[71715] <= 8'h10 ;
			data[71716] <= 8'h10 ;
			data[71717] <= 8'h10 ;
			data[71718] <= 8'h10 ;
			data[71719] <= 8'h10 ;
			data[71720] <= 8'h10 ;
			data[71721] <= 8'h10 ;
			data[71722] <= 8'h10 ;
			data[71723] <= 8'h10 ;
			data[71724] <= 8'h10 ;
			data[71725] <= 8'h10 ;
			data[71726] <= 8'h10 ;
			data[71727] <= 8'h10 ;
			data[71728] <= 8'h10 ;
			data[71729] <= 8'h10 ;
			data[71730] <= 8'h10 ;
			data[71731] <= 8'h10 ;
			data[71732] <= 8'h10 ;
			data[71733] <= 8'h10 ;
			data[71734] <= 8'h10 ;
			data[71735] <= 8'h10 ;
			data[71736] <= 8'h10 ;
			data[71737] <= 8'h10 ;
			data[71738] <= 8'h10 ;
			data[71739] <= 8'h10 ;
			data[71740] <= 8'h10 ;
			data[71741] <= 8'h10 ;
			data[71742] <= 8'h10 ;
			data[71743] <= 8'h10 ;
			data[71744] <= 8'h10 ;
			data[71745] <= 8'h10 ;
			data[71746] <= 8'h10 ;
			data[71747] <= 8'h10 ;
			data[71748] <= 8'h10 ;
			data[71749] <= 8'h10 ;
			data[71750] <= 8'h10 ;
			data[71751] <= 8'h10 ;
			data[71752] <= 8'h10 ;
			data[71753] <= 8'h10 ;
			data[71754] <= 8'h10 ;
			data[71755] <= 8'h10 ;
			data[71756] <= 8'h10 ;
			data[71757] <= 8'h10 ;
			data[71758] <= 8'h10 ;
			data[71759] <= 8'h10 ;
			data[71760] <= 8'h10 ;
			data[71761] <= 8'h10 ;
			data[71762] <= 8'h10 ;
			data[71763] <= 8'h10 ;
			data[71764] <= 8'h10 ;
			data[71765] <= 8'h10 ;
			data[71766] <= 8'h10 ;
			data[71767] <= 8'h10 ;
			data[71768] <= 8'h10 ;
			data[71769] <= 8'h10 ;
			data[71770] <= 8'h10 ;
			data[71771] <= 8'h10 ;
			data[71772] <= 8'h10 ;
			data[71773] <= 8'h10 ;
			data[71774] <= 8'h10 ;
			data[71775] <= 8'h10 ;
			data[71776] <= 8'h10 ;
			data[71777] <= 8'h10 ;
			data[71778] <= 8'h10 ;
			data[71779] <= 8'h10 ;
			data[71780] <= 8'h10 ;
			data[71781] <= 8'h10 ;
			data[71782] <= 8'h10 ;
			data[71783] <= 8'h10 ;
			data[71784] <= 8'h10 ;
			data[71785] <= 8'h10 ;
			data[71786] <= 8'h10 ;
			data[71787] <= 8'h10 ;
			data[71788] <= 8'h10 ;
			data[71789] <= 8'h10 ;
			data[71790] <= 8'h10 ;
			data[71791] <= 8'h10 ;
			data[71792] <= 8'h10 ;
			data[71793] <= 8'h10 ;
			data[71794] <= 8'h10 ;
			data[71795] <= 8'h10 ;
			data[71796] <= 8'h10 ;
			data[71797] <= 8'h10 ;
			data[71798] <= 8'h10 ;
			data[71799] <= 8'h10 ;
			data[71800] <= 8'h10 ;
			data[71801] <= 8'h10 ;
			data[71802] <= 8'h10 ;
			data[71803] <= 8'h10 ;
			data[71804] <= 8'h10 ;
			data[71805] <= 8'h10 ;
			data[71806] <= 8'h10 ;
			data[71807] <= 8'h10 ;
			data[71808] <= 8'h10 ;
			data[71809] <= 8'h10 ;
			data[71810] <= 8'h10 ;
			data[71811] <= 8'h10 ;
			data[71812] <= 8'h10 ;
			data[71813] <= 8'h10 ;
			data[71814] <= 8'h10 ;
			data[71815] <= 8'h10 ;
			data[71816] <= 8'h10 ;
			data[71817] <= 8'h10 ;
			data[71818] <= 8'h10 ;
			data[71819] <= 8'h10 ;
			data[71820] <= 8'h10 ;
			data[71821] <= 8'h10 ;
			data[71822] <= 8'h10 ;
			data[71823] <= 8'h10 ;
			data[71824] <= 8'h10 ;
			data[71825] <= 8'h10 ;
			data[71826] <= 8'h10 ;
			data[71827] <= 8'h10 ;
			data[71828] <= 8'h10 ;
			data[71829] <= 8'h10 ;
			data[71830] <= 8'h10 ;
			data[71831] <= 8'h10 ;
			data[71832] <= 8'h10 ;
			data[71833] <= 8'h10 ;
			data[71834] <= 8'h10 ;
			data[71835] <= 8'h10 ;
			data[71836] <= 8'h10 ;
			data[71837] <= 8'h10 ;
			data[71838] <= 8'h10 ;
			data[71839] <= 8'h10 ;
			data[71840] <= 8'h10 ;
			data[71841] <= 8'h10 ;
			data[71842] <= 8'h10 ;
			data[71843] <= 8'h10 ;
			data[71844] <= 8'h10 ;
			data[71845] <= 8'h10 ;
			data[71846] <= 8'h10 ;
			data[71847] <= 8'h10 ;
			data[71848] <= 8'h10 ;
			data[71849] <= 8'h10 ;
			data[71850] <= 8'h10 ;
			data[71851] <= 8'h10 ;
			data[71852] <= 8'h10 ;
			data[71853] <= 8'h10 ;
			data[71854] <= 8'h10 ;
			data[71855] <= 8'h10 ;
			data[71856] <= 8'h10 ;
			data[71857] <= 8'h10 ;
			data[71858] <= 8'h10 ;
			data[71859] <= 8'h10 ;
			data[71860] <= 8'h10 ;
			data[71861] <= 8'h10 ;
			data[71862] <= 8'h10 ;
			data[71863] <= 8'h10 ;
			data[71864] <= 8'h10 ;
			data[71865] <= 8'h10 ;
			data[71866] <= 8'h10 ;
			data[71867] <= 8'h10 ;
			data[71868] <= 8'h10 ;
			data[71869] <= 8'h10 ;
			data[71870] <= 8'h10 ;
			data[71871] <= 8'h10 ;
			data[71872] <= 8'h10 ;
			data[71873] <= 8'h10 ;
			data[71874] <= 8'h10 ;
			data[71875] <= 8'h10 ;
			data[71876] <= 8'h10 ;
			data[71877] <= 8'h10 ;
			data[71878] <= 8'h10 ;
			data[71879] <= 8'h10 ;
			data[71880] <= 8'h10 ;
			data[71881] <= 8'h10 ;
			data[71882] <= 8'h10 ;
			data[71883] <= 8'h10 ;
			data[71884] <= 8'h10 ;
			data[71885] <= 8'h10 ;
			data[71886] <= 8'h10 ;
			data[71887] <= 8'h10 ;
			data[71888] <= 8'h10 ;
			data[71889] <= 8'h10 ;
			data[71890] <= 8'h10 ;
			data[71891] <= 8'h10 ;
			data[71892] <= 8'h10 ;
			data[71893] <= 8'h10 ;
			data[71894] <= 8'h10 ;
			data[71895] <= 8'h10 ;
			data[71896] <= 8'h10 ;
			data[71897] <= 8'h10 ;
			data[71898] <= 8'h10 ;
			data[71899] <= 8'h10 ;
			data[71900] <= 8'h10 ;
			data[71901] <= 8'h10 ;
			data[71902] <= 8'h10 ;
			data[71903] <= 8'h10 ;
			data[71904] <= 8'h10 ;
			data[71905] <= 8'h10 ;
			data[71906] <= 8'h10 ;
			data[71907] <= 8'h10 ;
			data[71908] <= 8'h10 ;
			data[71909] <= 8'h10 ;
			data[71910] <= 8'h10 ;
			data[71911] <= 8'h10 ;
			data[71912] <= 8'h10 ;
			data[71913] <= 8'h10 ;
			data[71914] <= 8'h10 ;
			data[71915] <= 8'h10 ;
			data[71916] <= 8'h10 ;
			data[71917] <= 8'h10 ;
			data[71918] <= 8'h10 ;
			data[71919] <= 8'h10 ;
			data[71920] <= 8'h10 ;
			data[71921] <= 8'h10 ;
			data[71922] <= 8'h10 ;
			data[71923] <= 8'h10 ;
			data[71924] <= 8'h10 ;
			data[71925] <= 8'h10 ;
			data[71926] <= 8'h10 ;
			data[71927] <= 8'h10 ;
			data[71928] <= 8'h10 ;
			data[71929] <= 8'h10 ;
			data[71930] <= 8'h10 ;
			data[71931] <= 8'h10 ;
			data[71932] <= 8'h10 ;
			data[71933] <= 8'h10 ;
			data[71934] <= 8'h10 ;
			data[71935] <= 8'h10 ;
			data[71936] <= 8'h10 ;
			data[71937] <= 8'h10 ;
			data[71938] <= 8'h10 ;
			data[71939] <= 8'h10 ;
			data[71940] <= 8'h10 ;
			data[71941] <= 8'h10 ;
			data[71942] <= 8'h10 ;
			data[71943] <= 8'h10 ;
			data[71944] <= 8'h10 ;
			data[71945] <= 8'h10 ;
			data[71946] <= 8'h10 ;
			data[71947] <= 8'h10 ;
			data[71948] <= 8'h10 ;
			data[71949] <= 8'h10 ;
			data[71950] <= 8'h10 ;
			data[71951] <= 8'h10 ;
			data[71952] <= 8'h10 ;
			data[71953] <= 8'h10 ;
			data[71954] <= 8'h10 ;
			data[71955] <= 8'h10 ;
			data[71956] <= 8'h10 ;
			data[71957] <= 8'h10 ;
			data[71958] <= 8'h10 ;
			data[71959] <= 8'h10 ;
			data[71960] <= 8'h10 ;
			data[71961] <= 8'h10 ;
			data[71962] <= 8'h10 ;
			data[71963] <= 8'h10 ;
			data[71964] <= 8'h10 ;
			data[71965] <= 8'h10 ;
			data[71966] <= 8'h10 ;
			data[71967] <= 8'h10 ;
			data[71968] <= 8'h10 ;
			data[71969] <= 8'h10 ;
			data[71970] <= 8'h10 ;
			data[71971] <= 8'h10 ;
			data[71972] <= 8'h10 ;
			data[71973] <= 8'h10 ;
			data[71974] <= 8'h10 ;
			data[71975] <= 8'h10 ;
			data[71976] <= 8'h10 ;
			data[71977] <= 8'h10 ;
			data[71978] <= 8'h10 ;
			data[71979] <= 8'h10 ;
			data[71980] <= 8'h10 ;
			data[71981] <= 8'h10 ;
			data[71982] <= 8'h10 ;
			data[71983] <= 8'h10 ;
			data[71984] <= 8'h10 ;
			data[71985] <= 8'h10 ;
			data[71986] <= 8'h10 ;
			data[71987] <= 8'h10 ;
			data[71988] <= 8'h10 ;
			data[71989] <= 8'h10 ;
			data[71990] <= 8'h10 ;
			data[71991] <= 8'h10 ;
			data[71992] <= 8'h10 ;
			data[71993] <= 8'h10 ;
			data[71994] <= 8'h10 ;
			data[71995] <= 8'h10 ;
			data[71996] <= 8'h10 ;
			data[71997] <= 8'h10 ;
			data[71998] <= 8'h10 ;
			data[71999] <= 8'h10 ;
			data[72000] <= 8'h10 ;
			data[72001] <= 8'h10 ;
			data[72002] <= 8'h10 ;
			data[72003] <= 8'h10 ;
			data[72004] <= 8'h10 ;
			data[72005] <= 8'h10 ;
			data[72006] <= 8'h10 ;
			data[72007] <= 8'h10 ;
			data[72008] <= 8'h10 ;
			data[72009] <= 8'h10 ;
			data[72010] <= 8'h10 ;
			data[72011] <= 8'h10 ;
			data[72012] <= 8'h10 ;
			data[72013] <= 8'h10 ;
			data[72014] <= 8'h10 ;
			data[72015] <= 8'h10 ;
			data[72016] <= 8'h10 ;
			data[72017] <= 8'h10 ;
			data[72018] <= 8'h10 ;
			data[72019] <= 8'h10 ;
			data[72020] <= 8'h10 ;
			data[72021] <= 8'h10 ;
			data[72022] <= 8'h10 ;
			data[72023] <= 8'h10 ;
			data[72024] <= 8'h10 ;
			data[72025] <= 8'h10 ;
			data[72026] <= 8'h10 ;
			data[72027] <= 8'h10 ;
			data[72028] <= 8'h10 ;
			data[72029] <= 8'h10 ;
			data[72030] <= 8'h10 ;
			data[72031] <= 8'h10 ;
			data[72032] <= 8'h10 ;
			data[72033] <= 8'h10 ;
			data[72034] <= 8'h10 ;
			data[72035] <= 8'h10 ;
			data[72036] <= 8'h10 ;
			data[72037] <= 8'h10 ;
			data[72038] <= 8'h10 ;
			data[72039] <= 8'h10 ;
			data[72040] <= 8'h10 ;
			data[72041] <= 8'h10 ;
			data[72042] <= 8'h10 ;
			data[72043] <= 8'h10 ;
			data[72044] <= 8'h10 ;
			data[72045] <= 8'h10 ;
			data[72046] <= 8'h10 ;
			data[72047] <= 8'h10 ;
			data[72048] <= 8'h10 ;
			data[72049] <= 8'h10 ;
			data[72050] <= 8'h10 ;
			data[72051] <= 8'h10 ;
			data[72052] <= 8'h10 ;
			data[72053] <= 8'h10 ;
			data[72054] <= 8'h10 ;
			data[72055] <= 8'h10 ;
			data[72056] <= 8'h10 ;
			data[72057] <= 8'h10 ;
			data[72058] <= 8'h10 ;
			data[72059] <= 8'h10 ;
			data[72060] <= 8'h10 ;
			data[72061] <= 8'h10 ;
			data[72062] <= 8'h10 ;
			data[72063] <= 8'h10 ;
			data[72064] <= 8'h10 ;
			data[72065] <= 8'h10 ;
			data[72066] <= 8'h10 ;
			data[72067] <= 8'h10 ;
			data[72068] <= 8'h10 ;
			data[72069] <= 8'h10 ;
			data[72070] <= 8'h10 ;
			data[72071] <= 8'h10 ;
			data[72072] <= 8'h10 ;
			data[72073] <= 8'h10 ;
			data[72074] <= 8'h10 ;
			data[72075] <= 8'h10 ;
			data[72076] <= 8'h10 ;
			data[72077] <= 8'h10 ;
			data[72078] <= 8'h10 ;
			data[72079] <= 8'h10 ;
			data[72080] <= 8'h10 ;
			data[72081] <= 8'h10 ;
			data[72082] <= 8'h10 ;
			data[72083] <= 8'h10 ;
			data[72084] <= 8'h10 ;
			data[72085] <= 8'h10 ;
			data[72086] <= 8'h10 ;
			data[72087] <= 8'h10 ;
			data[72088] <= 8'h10 ;
			data[72089] <= 8'h10 ;
			data[72090] <= 8'h10 ;
			data[72091] <= 8'h10 ;
			data[72092] <= 8'h10 ;
			data[72093] <= 8'h10 ;
			data[72094] <= 8'h10 ;
			data[72095] <= 8'h10 ;
			data[72096] <= 8'h10 ;
			data[72097] <= 8'h10 ;
			data[72098] <= 8'h10 ;
			data[72099] <= 8'h10 ;
			data[72100] <= 8'h10 ;
			data[72101] <= 8'h10 ;
			data[72102] <= 8'h10 ;
			data[72103] <= 8'h10 ;
			data[72104] <= 8'h10 ;
			data[72105] <= 8'h10 ;
			data[72106] <= 8'h10 ;
			data[72107] <= 8'h10 ;
			data[72108] <= 8'h10 ;
			data[72109] <= 8'h10 ;
			data[72110] <= 8'h10 ;
			data[72111] <= 8'h10 ;
			data[72112] <= 8'h10 ;
			data[72113] <= 8'h10 ;
			data[72114] <= 8'h10 ;
			data[72115] <= 8'h10 ;
			data[72116] <= 8'h10 ;
			data[72117] <= 8'h10 ;
			data[72118] <= 8'h10 ;
			data[72119] <= 8'h10 ;
			data[72120] <= 8'h10 ;
			data[72121] <= 8'h10 ;
			data[72122] <= 8'h10 ;
			data[72123] <= 8'h10 ;
			data[72124] <= 8'h10 ;
			data[72125] <= 8'h10 ;
			data[72126] <= 8'h10 ;
			data[72127] <= 8'h10 ;
			data[72128] <= 8'h10 ;
			data[72129] <= 8'h10 ;
			data[72130] <= 8'h10 ;
			data[72131] <= 8'h10 ;
			data[72132] <= 8'h10 ;
			data[72133] <= 8'h10 ;
			data[72134] <= 8'h10 ;
			data[72135] <= 8'h10 ;
			data[72136] <= 8'h10 ;
			data[72137] <= 8'h10 ;
			data[72138] <= 8'h10 ;
			data[72139] <= 8'h10 ;
			data[72140] <= 8'h10 ;
			data[72141] <= 8'h10 ;
			data[72142] <= 8'h10 ;
			data[72143] <= 8'h10 ;
			data[72144] <= 8'h10 ;
			data[72145] <= 8'h10 ;
			data[72146] <= 8'h10 ;
			data[72147] <= 8'h10 ;
			data[72148] <= 8'h10 ;
			data[72149] <= 8'h10 ;
			data[72150] <= 8'h10 ;
			data[72151] <= 8'h10 ;
			data[72152] <= 8'h10 ;
			data[72153] <= 8'h10 ;
			data[72154] <= 8'h10 ;
			data[72155] <= 8'h10 ;
			data[72156] <= 8'h10 ;
			data[72157] <= 8'h10 ;
			data[72158] <= 8'h10 ;
			data[72159] <= 8'h10 ;
			data[72160] <= 8'h10 ;
			data[72161] <= 8'h10 ;
			data[72162] <= 8'h10 ;
			data[72163] <= 8'h10 ;
			data[72164] <= 8'h10 ;
			data[72165] <= 8'h10 ;
			data[72166] <= 8'h10 ;
			data[72167] <= 8'h10 ;
			data[72168] <= 8'h10 ;
			data[72169] <= 8'h10 ;
			data[72170] <= 8'h10 ;
			data[72171] <= 8'h10 ;
			data[72172] <= 8'h10 ;
			data[72173] <= 8'h10 ;
			data[72174] <= 8'h10 ;
			data[72175] <= 8'h10 ;
			data[72176] <= 8'h10 ;
			data[72177] <= 8'h10 ;
			data[72178] <= 8'h10 ;
			data[72179] <= 8'h10 ;
			data[72180] <= 8'h10 ;
			data[72181] <= 8'h10 ;
			data[72182] <= 8'h10 ;
			data[72183] <= 8'h10 ;
			data[72184] <= 8'h10 ;
			data[72185] <= 8'h10 ;
			data[72186] <= 8'h10 ;
			data[72187] <= 8'h10 ;
			data[72188] <= 8'h10 ;
			data[72189] <= 8'h10 ;
			data[72190] <= 8'h10 ;
			data[72191] <= 8'h10 ;
			data[72192] <= 8'h10 ;
			data[72193] <= 8'h10 ;
			data[72194] <= 8'h10 ;
			data[72195] <= 8'h10 ;
			data[72196] <= 8'h10 ;
			data[72197] <= 8'h10 ;
			data[72198] <= 8'h10 ;
			data[72199] <= 8'h10 ;
			data[72200] <= 8'h10 ;
			data[72201] <= 8'h10 ;
			data[72202] <= 8'h10 ;
			data[72203] <= 8'h10 ;
			data[72204] <= 8'h10 ;
			data[72205] <= 8'h10 ;
			data[72206] <= 8'h10 ;
			data[72207] <= 8'h10 ;
			data[72208] <= 8'h10 ;
			data[72209] <= 8'h10 ;
			data[72210] <= 8'h10 ;
			data[72211] <= 8'h10 ;
			data[72212] <= 8'h10 ;
			data[72213] <= 8'h10 ;
			data[72214] <= 8'h10 ;
			data[72215] <= 8'h10 ;
			data[72216] <= 8'h10 ;
			data[72217] <= 8'h10 ;
			data[72218] <= 8'h10 ;
			data[72219] <= 8'h10 ;
			data[72220] <= 8'h10 ;
			data[72221] <= 8'h10 ;
			data[72222] <= 8'h10 ;
			data[72223] <= 8'h10 ;
			data[72224] <= 8'h10 ;
			data[72225] <= 8'h10 ;
			data[72226] <= 8'h10 ;
			data[72227] <= 8'h10 ;
			data[72228] <= 8'h10 ;
			data[72229] <= 8'h10 ;
			data[72230] <= 8'h10 ;
			data[72231] <= 8'h10 ;
			data[72232] <= 8'h10 ;
			data[72233] <= 8'h10 ;
			data[72234] <= 8'h10 ;
			data[72235] <= 8'h10 ;
			data[72236] <= 8'h10 ;
			data[72237] <= 8'h10 ;
			data[72238] <= 8'h10 ;
			data[72239] <= 8'h10 ;
			data[72240] <= 8'h10 ;
			data[72241] <= 8'h10 ;
			data[72242] <= 8'h10 ;
			data[72243] <= 8'h10 ;
			data[72244] <= 8'h10 ;
			data[72245] <= 8'h10 ;
			data[72246] <= 8'h10 ;
			data[72247] <= 8'h10 ;
			data[72248] <= 8'h10 ;
			data[72249] <= 8'h10 ;
			data[72250] <= 8'h10 ;
			data[72251] <= 8'h10 ;
			data[72252] <= 8'h10 ;
			data[72253] <= 8'h10 ;
			data[72254] <= 8'h10 ;
			data[72255] <= 8'h10 ;
			data[72256] <= 8'h10 ;
			data[72257] <= 8'h10 ;
			data[72258] <= 8'h10 ;
			data[72259] <= 8'h10 ;
			data[72260] <= 8'h10 ;
			data[72261] <= 8'h10 ;
			data[72262] <= 8'h10 ;
			data[72263] <= 8'h10 ;
			data[72264] <= 8'h10 ;
			data[72265] <= 8'h10 ;
			data[72266] <= 8'h10 ;
			data[72267] <= 8'h10 ;
			data[72268] <= 8'h10 ;
			data[72269] <= 8'h10 ;
			data[72270] <= 8'h10 ;
			data[72271] <= 8'h10 ;
			data[72272] <= 8'h10 ;
			data[72273] <= 8'h10 ;
			data[72274] <= 8'h10 ;
			data[72275] <= 8'h10 ;
			data[72276] <= 8'h10 ;
			data[72277] <= 8'h10 ;
			data[72278] <= 8'h10 ;
			data[72279] <= 8'h10 ;
			data[72280] <= 8'h10 ;
			data[72281] <= 8'h10 ;
			data[72282] <= 8'h10 ;
			data[72283] <= 8'h10 ;
			data[72284] <= 8'h10 ;
			data[72285] <= 8'h10 ;
			data[72286] <= 8'h10 ;
			data[72287] <= 8'h10 ;
			data[72288] <= 8'h10 ;
			data[72289] <= 8'h10 ;
			data[72290] <= 8'h10 ;
			data[72291] <= 8'h10 ;
			data[72292] <= 8'h10 ;
			data[72293] <= 8'h10 ;
			data[72294] <= 8'h10 ;
			data[72295] <= 8'h10 ;
			data[72296] <= 8'h10 ;
			data[72297] <= 8'h10 ;
			data[72298] <= 8'h10 ;
			data[72299] <= 8'h10 ;
			data[72300] <= 8'h10 ;
			data[72301] <= 8'h10 ;
			data[72302] <= 8'h10 ;
			data[72303] <= 8'h10 ;
			data[72304] <= 8'h10 ;
			data[72305] <= 8'h10 ;
			data[72306] <= 8'h10 ;
			data[72307] <= 8'h10 ;
			data[72308] <= 8'h10 ;
			data[72309] <= 8'h10 ;
			data[72310] <= 8'h10 ;
			data[72311] <= 8'h10 ;
			data[72312] <= 8'h10 ;
			data[72313] <= 8'h10 ;
			data[72314] <= 8'h10 ;
			data[72315] <= 8'h10 ;
			data[72316] <= 8'h10 ;
			data[72317] <= 8'h10 ;
			data[72318] <= 8'h10 ;
			data[72319] <= 8'h10 ;
			data[72320] <= 8'h10 ;
			data[72321] <= 8'h10 ;
			data[72322] <= 8'h10 ;
			data[72323] <= 8'h10 ;
			data[72324] <= 8'h10 ;
			data[72325] <= 8'h10 ;
			data[72326] <= 8'h10 ;
			data[72327] <= 8'h10 ;
			data[72328] <= 8'h10 ;
			data[72329] <= 8'h10 ;
			data[72330] <= 8'h10 ;
			data[72331] <= 8'h10 ;
			data[72332] <= 8'h10 ;
			data[72333] <= 8'h10 ;
			data[72334] <= 8'h10 ;
			data[72335] <= 8'h10 ;
			data[72336] <= 8'h10 ;
			data[72337] <= 8'h10 ;
			data[72338] <= 8'h10 ;
			data[72339] <= 8'h10 ;
			data[72340] <= 8'h10 ;
			data[72341] <= 8'h10 ;
			data[72342] <= 8'h10 ;
			data[72343] <= 8'h10 ;
			data[72344] <= 8'h10 ;
			data[72345] <= 8'h10 ;
			data[72346] <= 8'h10 ;
			data[72347] <= 8'h10 ;
			data[72348] <= 8'h10 ;
			data[72349] <= 8'h10 ;
			data[72350] <= 8'h10 ;
			data[72351] <= 8'h10 ;
			data[72352] <= 8'h10 ;
			data[72353] <= 8'h10 ;
			data[72354] <= 8'h10 ;
			data[72355] <= 8'h10 ;
			data[72356] <= 8'h10 ;
			data[72357] <= 8'h10 ;
			data[72358] <= 8'h10 ;
			data[72359] <= 8'h10 ;
			data[72360] <= 8'h10 ;
			data[72361] <= 8'h10 ;
			data[72362] <= 8'h10 ;
			data[72363] <= 8'h10 ;
			data[72364] <= 8'h10 ;
			data[72365] <= 8'h10 ;
			data[72366] <= 8'h10 ;
			data[72367] <= 8'h10 ;
			data[72368] <= 8'h10 ;
			data[72369] <= 8'h10 ;
			data[72370] <= 8'h10 ;
			data[72371] <= 8'h10 ;
			data[72372] <= 8'h10 ;
			data[72373] <= 8'h10 ;
			data[72374] <= 8'h10 ;
			data[72375] <= 8'h10 ;
			data[72376] <= 8'h10 ;
			data[72377] <= 8'h10 ;
			data[72378] <= 8'h10 ;
			data[72379] <= 8'h10 ;
			data[72380] <= 8'h10 ;
			data[72381] <= 8'h10 ;
			data[72382] <= 8'h10 ;
			data[72383] <= 8'h10 ;
			data[72384] <= 8'h10 ;
			data[72385] <= 8'h10 ;
			data[72386] <= 8'h10 ;
			data[72387] <= 8'h10 ;
			data[72388] <= 8'h10 ;
			data[72389] <= 8'h10 ;
			data[72390] <= 8'h10 ;
			data[72391] <= 8'h10 ;
			data[72392] <= 8'h10 ;
			data[72393] <= 8'h10 ;
			data[72394] <= 8'h10 ;
			data[72395] <= 8'h10 ;
			data[72396] <= 8'h10 ;
			data[72397] <= 8'h10 ;
			data[72398] <= 8'h10 ;
			data[72399] <= 8'h10 ;
			data[72400] <= 8'h10 ;
			data[72401] <= 8'h10 ;
			data[72402] <= 8'h10 ;
			data[72403] <= 8'h10 ;
			data[72404] <= 8'h10 ;
			data[72405] <= 8'h10 ;
			data[72406] <= 8'h10 ;
			data[72407] <= 8'h10 ;
			data[72408] <= 8'h10 ;
			data[72409] <= 8'h10 ;
			data[72410] <= 8'h10 ;
			data[72411] <= 8'h10 ;
			data[72412] <= 8'h10 ;
			data[72413] <= 8'h10 ;
			data[72414] <= 8'h10 ;
			data[72415] <= 8'h10 ;
			data[72416] <= 8'h10 ;
			data[72417] <= 8'h10 ;
			data[72418] <= 8'h10 ;
			data[72419] <= 8'h10 ;
			data[72420] <= 8'h10 ;
			data[72421] <= 8'h10 ;
			data[72422] <= 8'h10 ;
			data[72423] <= 8'h10 ;
			data[72424] <= 8'h10 ;
			data[72425] <= 8'h10 ;
			data[72426] <= 8'h10 ;
			data[72427] <= 8'h10 ;
			data[72428] <= 8'h10 ;
			data[72429] <= 8'h10 ;
			data[72430] <= 8'h10 ;
			data[72431] <= 8'h10 ;
			data[72432] <= 8'h10 ;
			data[72433] <= 8'h10 ;
			data[72434] <= 8'h10 ;
			data[72435] <= 8'h10 ;
			data[72436] <= 8'h10 ;
			data[72437] <= 8'h10 ;
			data[72438] <= 8'h10 ;
			data[72439] <= 8'h10 ;
			data[72440] <= 8'h10 ;
			data[72441] <= 8'h10 ;
			data[72442] <= 8'h10 ;
			data[72443] <= 8'h10 ;
			data[72444] <= 8'h10 ;
			data[72445] <= 8'h10 ;
			data[72446] <= 8'h10 ;
			data[72447] <= 8'h10 ;
			data[72448] <= 8'h10 ;
			data[72449] <= 8'h10 ;
			data[72450] <= 8'h10 ;
			data[72451] <= 8'h10 ;
			data[72452] <= 8'h10 ;
			data[72453] <= 8'h10 ;
			data[72454] <= 8'h10 ;
			data[72455] <= 8'h10 ;
			data[72456] <= 8'h10 ;
			data[72457] <= 8'h10 ;
			data[72458] <= 8'h10 ;
			data[72459] <= 8'h10 ;
			data[72460] <= 8'h10 ;
			data[72461] <= 8'h10 ;
			data[72462] <= 8'h10 ;
			data[72463] <= 8'h10 ;
			data[72464] <= 8'h10 ;
			data[72465] <= 8'h10 ;
			data[72466] <= 8'h10 ;
			data[72467] <= 8'h10 ;
			data[72468] <= 8'h10 ;
			data[72469] <= 8'h10 ;
			data[72470] <= 8'h10 ;
			data[72471] <= 8'h10 ;
			data[72472] <= 8'h10 ;
			data[72473] <= 8'h10 ;
			data[72474] <= 8'h10 ;
			data[72475] <= 8'h10 ;
			data[72476] <= 8'h10 ;
			data[72477] <= 8'h10 ;
			data[72478] <= 8'h10 ;
			data[72479] <= 8'h10 ;
			data[72480] <= 8'h10 ;
			data[72481] <= 8'h10 ;
			data[72482] <= 8'h10 ;
			data[72483] <= 8'h10 ;
			data[72484] <= 8'h10 ;
			data[72485] <= 8'h10 ;
			data[72486] <= 8'h10 ;
			data[72487] <= 8'h10 ;
			data[72488] <= 8'h10 ;
			data[72489] <= 8'h10 ;
			data[72490] <= 8'h10 ;
			data[72491] <= 8'h10 ;
			data[72492] <= 8'h10 ;
			data[72493] <= 8'h10 ;
			data[72494] <= 8'h10 ;
			data[72495] <= 8'h10 ;
			data[72496] <= 8'h10 ;
			data[72497] <= 8'h10 ;
			data[72498] <= 8'h10 ;
			data[72499] <= 8'h10 ;
			data[72500] <= 8'h10 ;
			data[72501] <= 8'h10 ;
			data[72502] <= 8'h10 ;
			data[72503] <= 8'h10 ;
			data[72504] <= 8'h10 ;
			data[72505] <= 8'h10 ;
			data[72506] <= 8'h10 ;
			data[72507] <= 8'h10 ;
			data[72508] <= 8'h10 ;
			data[72509] <= 8'h10 ;
			data[72510] <= 8'h10 ;
			data[72511] <= 8'h10 ;
			data[72512] <= 8'h10 ;
			data[72513] <= 8'h10 ;
			data[72514] <= 8'h10 ;
			data[72515] <= 8'h10 ;
			data[72516] <= 8'h10 ;
			data[72517] <= 8'h10 ;
			data[72518] <= 8'h10 ;
			data[72519] <= 8'h10 ;
			data[72520] <= 8'h10 ;
			data[72521] <= 8'h10 ;
			data[72522] <= 8'h10 ;
			data[72523] <= 8'h10 ;
			data[72524] <= 8'h10 ;
			data[72525] <= 8'h10 ;
			data[72526] <= 8'h10 ;
			data[72527] <= 8'h10 ;
			data[72528] <= 8'h10 ;
			data[72529] <= 8'h10 ;
			data[72530] <= 8'h10 ;
			data[72531] <= 8'h10 ;
			data[72532] <= 8'h10 ;
			data[72533] <= 8'h10 ;
			data[72534] <= 8'h10 ;
			data[72535] <= 8'h10 ;
			data[72536] <= 8'h10 ;
			data[72537] <= 8'h10 ;
			data[72538] <= 8'h10 ;
			data[72539] <= 8'h10 ;
			data[72540] <= 8'h10 ;
			data[72541] <= 8'h10 ;
			data[72542] <= 8'h10 ;
			data[72543] <= 8'h10 ;
			data[72544] <= 8'h10 ;
			data[72545] <= 8'h10 ;
			data[72546] <= 8'h10 ;
			data[72547] <= 8'h10 ;
			data[72548] <= 8'h10 ;
			data[72549] <= 8'h10 ;
			data[72550] <= 8'h10 ;
			data[72551] <= 8'h10 ;
			data[72552] <= 8'h10 ;
			data[72553] <= 8'h10 ;
			data[72554] <= 8'h10 ;
			data[72555] <= 8'h10 ;
			data[72556] <= 8'h10 ;
			data[72557] <= 8'h10 ;
			data[72558] <= 8'h10 ;
			data[72559] <= 8'h10 ;
			data[72560] <= 8'h10 ;
			data[72561] <= 8'h10 ;
			data[72562] <= 8'h10 ;
			data[72563] <= 8'h10 ;
			data[72564] <= 8'h10 ;
			data[72565] <= 8'h10 ;
			data[72566] <= 8'h10 ;
			data[72567] <= 8'h10 ;
			data[72568] <= 8'h10 ;
			data[72569] <= 8'h10 ;
			data[72570] <= 8'h10 ;
			data[72571] <= 8'h10 ;
			data[72572] <= 8'h10 ;
			data[72573] <= 8'h10 ;
			data[72574] <= 8'h10 ;
			data[72575] <= 8'h10 ;
			data[72576] <= 8'h10 ;
			data[72577] <= 8'h10 ;
			data[72578] <= 8'h10 ;
			data[72579] <= 8'h10 ;
			data[72580] <= 8'h10 ;
			data[72581] <= 8'h10 ;
			data[72582] <= 8'h10 ;
			data[72583] <= 8'h10 ;
			data[72584] <= 8'h10 ;
			data[72585] <= 8'h10 ;
			data[72586] <= 8'h10 ;
			data[72587] <= 8'h10 ;
			data[72588] <= 8'h10 ;
			data[72589] <= 8'h10 ;
			data[72590] <= 8'h10 ;
			data[72591] <= 8'h10 ;
			data[72592] <= 8'h10 ;
			data[72593] <= 8'h10 ;
			data[72594] <= 8'h10 ;
			data[72595] <= 8'h10 ;
			data[72596] <= 8'h10 ;
			data[72597] <= 8'h10 ;
			data[72598] <= 8'h10 ;
			data[72599] <= 8'h10 ;
			data[72600] <= 8'h10 ;
			data[72601] <= 8'h10 ;
			data[72602] <= 8'h10 ;
			data[72603] <= 8'h10 ;
			data[72604] <= 8'h10 ;
			data[72605] <= 8'h10 ;
			data[72606] <= 8'h10 ;
			data[72607] <= 8'h10 ;
			data[72608] <= 8'h10 ;
			data[72609] <= 8'h10 ;
			data[72610] <= 8'h10 ;
			data[72611] <= 8'h10 ;
			data[72612] <= 8'h10 ;
			data[72613] <= 8'h10 ;
			data[72614] <= 8'h10 ;
			data[72615] <= 8'h10 ;
			data[72616] <= 8'h10 ;
			data[72617] <= 8'h10 ;
			data[72618] <= 8'h10 ;
			data[72619] <= 8'h10 ;
			data[72620] <= 8'h10 ;
			data[72621] <= 8'h10 ;
			data[72622] <= 8'h10 ;
			data[72623] <= 8'h10 ;
			data[72624] <= 8'h10 ;
			data[72625] <= 8'h10 ;
			data[72626] <= 8'h10 ;
			data[72627] <= 8'h10 ;
			data[72628] <= 8'h10 ;
			data[72629] <= 8'h10 ;
			data[72630] <= 8'h10 ;
			data[72631] <= 8'h10 ;
			data[72632] <= 8'h10 ;
			data[72633] <= 8'h10 ;
			data[72634] <= 8'h10 ;
			data[72635] <= 8'h10 ;
			data[72636] <= 8'h10 ;
			data[72637] <= 8'h10 ;
			data[72638] <= 8'h10 ;
			data[72639] <= 8'h10 ;
			data[72640] <= 8'h10 ;
			data[72641] <= 8'h10 ;
			data[72642] <= 8'h10 ;
			data[72643] <= 8'h10 ;
			data[72644] <= 8'h10 ;
			data[72645] <= 8'h10 ;
			data[72646] <= 8'h10 ;
			data[72647] <= 8'h10 ;
			data[72648] <= 8'h10 ;
			data[72649] <= 8'h10 ;
			data[72650] <= 8'h10 ;
			data[72651] <= 8'h10 ;
			data[72652] <= 8'h10 ;
			data[72653] <= 8'h10 ;
			data[72654] <= 8'h10 ;
			data[72655] <= 8'h10 ;
			data[72656] <= 8'h10 ;
			data[72657] <= 8'h10 ;
			data[72658] <= 8'h10 ;
			data[72659] <= 8'h10 ;
			data[72660] <= 8'h10 ;
			data[72661] <= 8'h10 ;
			data[72662] <= 8'h10 ;
			data[72663] <= 8'h10 ;
			data[72664] <= 8'h10 ;
			data[72665] <= 8'h10 ;
			data[72666] <= 8'h10 ;
			data[72667] <= 8'h10 ;
			data[72668] <= 8'h10 ;
			data[72669] <= 8'h10 ;
			data[72670] <= 8'h10 ;
			data[72671] <= 8'h10 ;
			data[72672] <= 8'h10 ;
			data[72673] <= 8'h10 ;
			data[72674] <= 8'h10 ;
			data[72675] <= 8'h10 ;
			data[72676] <= 8'h10 ;
			data[72677] <= 8'h10 ;
			data[72678] <= 8'h10 ;
			data[72679] <= 8'h10 ;
			data[72680] <= 8'h10 ;
			data[72681] <= 8'h10 ;
			data[72682] <= 8'h10 ;
			data[72683] <= 8'h10 ;
			data[72684] <= 8'h10 ;
			data[72685] <= 8'h10 ;
			data[72686] <= 8'h10 ;
			data[72687] <= 8'h10 ;
			data[72688] <= 8'h10 ;
			data[72689] <= 8'h10 ;
			data[72690] <= 8'h10 ;
			data[72691] <= 8'h10 ;
			data[72692] <= 8'h10 ;
			data[72693] <= 8'h10 ;
			data[72694] <= 8'h10 ;
			data[72695] <= 8'h10 ;
			data[72696] <= 8'h10 ;
			data[72697] <= 8'h10 ;
			data[72698] <= 8'h10 ;
			data[72699] <= 8'h10 ;
			data[72700] <= 8'h10 ;
			data[72701] <= 8'h10 ;
			data[72702] <= 8'h10 ;
			data[72703] <= 8'h10 ;
			data[72704] <= 8'h10 ;
			data[72705] <= 8'h10 ;
			data[72706] <= 8'h10 ;
			data[72707] <= 8'h10 ;
			data[72708] <= 8'h10 ;
			data[72709] <= 8'h10 ;
			data[72710] <= 8'h10 ;
			data[72711] <= 8'h10 ;
			data[72712] <= 8'h10 ;
			data[72713] <= 8'h10 ;
			data[72714] <= 8'h10 ;
			data[72715] <= 8'h10 ;
			data[72716] <= 8'h10 ;
			data[72717] <= 8'h10 ;
			data[72718] <= 8'h10 ;
			data[72719] <= 8'h10 ;
			data[72720] <= 8'h10 ;
			data[72721] <= 8'h10 ;
			data[72722] <= 8'h10 ;
			data[72723] <= 8'h10 ;
			data[72724] <= 8'h10 ;
			data[72725] <= 8'h10 ;
			data[72726] <= 8'h10 ;
			data[72727] <= 8'h10 ;
			data[72728] <= 8'h10 ;
			data[72729] <= 8'h10 ;
			data[72730] <= 8'h10 ;
			data[72731] <= 8'h10 ;
			data[72732] <= 8'h10 ;
			data[72733] <= 8'h10 ;
			data[72734] <= 8'h10 ;
			data[72735] <= 8'h10 ;
			data[72736] <= 8'h10 ;
			data[72737] <= 8'h10 ;
			data[72738] <= 8'h10 ;
			data[72739] <= 8'h10 ;
			data[72740] <= 8'h10 ;
			data[72741] <= 8'h10 ;
			data[72742] <= 8'h10 ;
			data[72743] <= 8'h10 ;
			data[72744] <= 8'h10 ;
			data[72745] <= 8'h10 ;
			data[72746] <= 8'h10 ;
			data[72747] <= 8'h10 ;
			data[72748] <= 8'h10 ;
			data[72749] <= 8'h10 ;
			data[72750] <= 8'h10 ;
			data[72751] <= 8'h10 ;
			data[72752] <= 8'h10 ;
			data[72753] <= 8'h10 ;
			data[72754] <= 8'h10 ;
			data[72755] <= 8'h10 ;
			data[72756] <= 8'h10 ;
			data[72757] <= 8'h10 ;
			data[72758] <= 8'h10 ;
			data[72759] <= 8'h10 ;
			data[72760] <= 8'h10 ;
			data[72761] <= 8'h10 ;
			data[72762] <= 8'h10 ;
			data[72763] <= 8'h10 ;
			data[72764] <= 8'h10 ;
			data[72765] <= 8'h10 ;
			data[72766] <= 8'h10 ;
			data[72767] <= 8'h10 ;
			data[72768] <= 8'h10 ;
			data[72769] <= 8'h10 ;
			data[72770] <= 8'h10 ;
			data[72771] <= 8'h10 ;
			data[72772] <= 8'h10 ;
			data[72773] <= 8'h10 ;
			data[72774] <= 8'h10 ;
			data[72775] <= 8'h10 ;
			data[72776] <= 8'h10 ;
			data[72777] <= 8'h10 ;
			data[72778] <= 8'h10 ;
			data[72779] <= 8'h10 ;
			data[72780] <= 8'h10 ;
			data[72781] <= 8'h10 ;
			data[72782] <= 8'h10 ;
			data[72783] <= 8'h10 ;
			data[72784] <= 8'h10 ;
			data[72785] <= 8'h10 ;
			data[72786] <= 8'h10 ;
			data[72787] <= 8'h10 ;
			data[72788] <= 8'h10 ;
			data[72789] <= 8'h10 ;
			data[72790] <= 8'h10 ;
			data[72791] <= 8'h10 ;
			data[72792] <= 8'h10 ;
			data[72793] <= 8'h10 ;
			data[72794] <= 8'h10 ;
			data[72795] <= 8'h10 ;
			data[72796] <= 8'h10 ;
			data[72797] <= 8'h10 ;
			data[72798] <= 8'h10 ;
			data[72799] <= 8'h10 ;
			data[72800] <= 8'h10 ;
			data[72801] <= 8'h10 ;
			data[72802] <= 8'h10 ;
			data[72803] <= 8'h10 ;
			data[72804] <= 8'h10 ;
			data[72805] <= 8'h10 ;
			data[72806] <= 8'h10 ;
			data[72807] <= 8'h10 ;
			data[72808] <= 8'h10 ;
			data[72809] <= 8'h10 ;
			data[72810] <= 8'h10 ;
			data[72811] <= 8'h10 ;
			data[72812] <= 8'h10 ;
			data[72813] <= 8'h10 ;
			data[72814] <= 8'h10 ;
			data[72815] <= 8'h10 ;
			data[72816] <= 8'h10 ;
			data[72817] <= 8'h10 ;
			data[72818] <= 8'h10 ;
			data[72819] <= 8'h10 ;
			data[72820] <= 8'h10 ;
			data[72821] <= 8'h10 ;
			data[72822] <= 8'h10 ;
			data[72823] <= 8'h10 ;
			data[72824] <= 8'h10 ;
			data[72825] <= 8'h10 ;
			data[72826] <= 8'h10 ;
			data[72827] <= 8'h10 ;
			data[72828] <= 8'h10 ;
			data[72829] <= 8'h10 ;
			data[72830] <= 8'h10 ;
			data[72831] <= 8'h10 ;
			data[72832] <= 8'h10 ;
			data[72833] <= 8'h10 ;
			data[72834] <= 8'h10 ;
			data[72835] <= 8'h10 ;
			data[72836] <= 8'h10 ;
			data[72837] <= 8'h10 ;
			data[72838] <= 8'h10 ;
			data[72839] <= 8'h10 ;
			data[72840] <= 8'h10 ;
			data[72841] <= 8'h10 ;
			data[72842] <= 8'h10 ;
			data[72843] <= 8'h10 ;
			data[72844] <= 8'h10 ;
			data[72845] <= 8'h10 ;
			data[72846] <= 8'h10 ;
			data[72847] <= 8'h10 ;
			data[72848] <= 8'h10 ;
			data[72849] <= 8'h10 ;
			data[72850] <= 8'h10 ;
			data[72851] <= 8'h10 ;
			data[72852] <= 8'h10 ;
			data[72853] <= 8'h10 ;
			data[72854] <= 8'h10 ;
			data[72855] <= 8'h10 ;
			data[72856] <= 8'h10 ;
			data[72857] <= 8'h10 ;
			data[72858] <= 8'h10 ;
			data[72859] <= 8'h10 ;
			data[72860] <= 8'h10 ;
			data[72861] <= 8'h10 ;
			data[72862] <= 8'h10 ;
			data[72863] <= 8'h10 ;
			data[72864] <= 8'h10 ;
			data[72865] <= 8'h10 ;
			data[72866] <= 8'h10 ;
			data[72867] <= 8'h10 ;
			data[72868] <= 8'h10 ;
			data[72869] <= 8'h10 ;
			data[72870] <= 8'h10 ;
			data[72871] <= 8'h10 ;
			data[72872] <= 8'h10 ;
			data[72873] <= 8'h10 ;
			data[72874] <= 8'h10 ;
			data[72875] <= 8'h10 ;
			data[72876] <= 8'h10 ;
			data[72877] <= 8'h10 ;
			data[72878] <= 8'h10 ;
			data[72879] <= 8'h10 ;
			data[72880] <= 8'h10 ;
			data[72881] <= 8'h10 ;
			data[72882] <= 8'h10 ;
			data[72883] <= 8'h10 ;
			data[72884] <= 8'h10 ;
			data[72885] <= 8'h10 ;
			data[72886] <= 8'h10 ;
			data[72887] <= 8'h10 ;
			data[72888] <= 8'h10 ;
			data[72889] <= 8'h10 ;
			data[72890] <= 8'h10 ;
			data[72891] <= 8'h10 ;
			data[72892] <= 8'h10 ;
			data[72893] <= 8'h10 ;
			data[72894] <= 8'h10 ;
			data[72895] <= 8'h10 ;
			data[72896] <= 8'h10 ;
			data[72897] <= 8'h10 ;
			data[72898] <= 8'h10 ;
			data[72899] <= 8'h10 ;
			data[72900] <= 8'h10 ;
			data[72901] <= 8'h10 ;
			data[72902] <= 8'h10 ;
			data[72903] <= 8'h10 ;
			data[72904] <= 8'h10 ;
			data[72905] <= 8'h10 ;
			data[72906] <= 8'h10 ;
			data[72907] <= 8'h10 ;
			data[72908] <= 8'h10 ;
			data[72909] <= 8'h10 ;
			data[72910] <= 8'h10 ;
			data[72911] <= 8'h10 ;
			data[72912] <= 8'h10 ;
			data[72913] <= 8'h10 ;
			data[72914] <= 8'h10 ;
			data[72915] <= 8'h10 ;
			data[72916] <= 8'h10 ;
			data[72917] <= 8'h10 ;
			data[72918] <= 8'h10 ;
			data[72919] <= 8'h10 ;
			data[72920] <= 8'h10 ;
			data[72921] <= 8'h10 ;
			data[72922] <= 8'h10 ;
			data[72923] <= 8'h10 ;
			data[72924] <= 8'h10 ;
			data[72925] <= 8'h10 ;
			data[72926] <= 8'h10 ;
			data[72927] <= 8'h10 ;
			data[72928] <= 8'h10 ;
			data[72929] <= 8'h10 ;
			data[72930] <= 8'h10 ;
			data[72931] <= 8'h10 ;
			data[72932] <= 8'h10 ;
			data[72933] <= 8'h10 ;
			data[72934] <= 8'h10 ;
			data[72935] <= 8'h10 ;
			data[72936] <= 8'h10 ;
			data[72937] <= 8'h10 ;
			data[72938] <= 8'h10 ;
			data[72939] <= 8'h10 ;
			data[72940] <= 8'h10 ;
			data[72941] <= 8'h10 ;
			data[72942] <= 8'h10 ;
			data[72943] <= 8'h10 ;
			data[72944] <= 8'h10 ;
			data[72945] <= 8'h10 ;
			data[72946] <= 8'h10 ;
			data[72947] <= 8'h10 ;
			data[72948] <= 8'h10 ;
			data[72949] <= 8'h10 ;
			data[72950] <= 8'h10 ;
			data[72951] <= 8'h10 ;
			data[72952] <= 8'h10 ;
			data[72953] <= 8'h10 ;
			data[72954] <= 8'h10 ;
			data[72955] <= 8'h10 ;
			data[72956] <= 8'h10 ;
			data[72957] <= 8'h10 ;
			data[72958] <= 8'h10 ;
			data[72959] <= 8'h10 ;
			data[72960] <= 8'h10 ;
			data[72961] <= 8'h10 ;
			data[72962] <= 8'h10 ;
			data[72963] <= 8'h10 ;
			data[72964] <= 8'h10 ;
			data[72965] <= 8'h10 ;
			data[72966] <= 8'h10 ;
			data[72967] <= 8'h10 ;
			data[72968] <= 8'h10 ;
			data[72969] <= 8'h10 ;
			data[72970] <= 8'h10 ;
			data[72971] <= 8'h10 ;
			data[72972] <= 8'h10 ;
			data[72973] <= 8'h10 ;
			data[72974] <= 8'h10 ;
			data[72975] <= 8'h10 ;
			data[72976] <= 8'h10 ;
			data[72977] <= 8'h10 ;
			data[72978] <= 8'h10 ;
			data[72979] <= 8'h10 ;
			data[72980] <= 8'h10 ;
			data[72981] <= 8'h10 ;
			data[72982] <= 8'h10 ;
			data[72983] <= 8'h10 ;
			data[72984] <= 8'h10 ;
			data[72985] <= 8'h10 ;
			data[72986] <= 8'h10 ;
			data[72987] <= 8'h10 ;
			data[72988] <= 8'h10 ;
			data[72989] <= 8'h10 ;
			data[72990] <= 8'h10 ;
			data[72991] <= 8'h10 ;
			data[72992] <= 8'h10 ;
			data[72993] <= 8'h10 ;
			data[72994] <= 8'h10 ;
			data[72995] <= 8'h10 ;
			data[72996] <= 8'h10 ;
			data[72997] <= 8'h10 ;
			data[72998] <= 8'h10 ;
			data[72999] <= 8'h10 ;
			data[73000] <= 8'h10 ;
			data[73001] <= 8'h10 ;
			data[73002] <= 8'h10 ;
			data[73003] <= 8'h10 ;
			data[73004] <= 8'h10 ;
			data[73005] <= 8'h10 ;
			data[73006] <= 8'h10 ;
			data[73007] <= 8'h10 ;
			data[73008] <= 8'h10 ;
			data[73009] <= 8'h10 ;
			data[73010] <= 8'h10 ;
			data[73011] <= 8'h10 ;
			data[73012] <= 8'h10 ;
			data[73013] <= 8'h10 ;
			data[73014] <= 8'h10 ;
			data[73015] <= 8'h10 ;
			data[73016] <= 8'h10 ;
			data[73017] <= 8'h10 ;
			data[73018] <= 8'h10 ;
			data[73019] <= 8'h10 ;
			data[73020] <= 8'h10 ;
			data[73021] <= 8'h10 ;
			data[73022] <= 8'h10 ;
			data[73023] <= 8'h10 ;
			data[73024] <= 8'h10 ;
			data[73025] <= 8'h10 ;
			data[73026] <= 8'h10 ;
			data[73027] <= 8'h10 ;
			data[73028] <= 8'h10 ;
			data[73029] <= 8'h10 ;
			data[73030] <= 8'h10 ;
			data[73031] <= 8'h10 ;
			data[73032] <= 8'h10 ;
			data[73033] <= 8'h10 ;
			data[73034] <= 8'h10 ;
			data[73035] <= 8'h10 ;
			data[73036] <= 8'h10 ;
			data[73037] <= 8'h10 ;
			data[73038] <= 8'h10 ;
			data[73039] <= 8'h10 ;
			data[73040] <= 8'h10 ;
			data[73041] <= 8'h10 ;
			data[73042] <= 8'h10 ;
			data[73043] <= 8'h10 ;
			data[73044] <= 8'h10 ;
			data[73045] <= 8'h10 ;
			data[73046] <= 8'h10 ;
			data[73047] <= 8'h10 ;
			data[73048] <= 8'h10 ;
			data[73049] <= 8'h10 ;
			data[73050] <= 8'h10 ;
			data[73051] <= 8'h10 ;
			data[73052] <= 8'h10 ;
			data[73053] <= 8'h10 ;
			data[73054] <= 8'h10 ;
			data[73055] <= 8'h10 ;
			data[73056] <= 8'h10 ;
			data[73057] <= 8'h10 ;
			data[73058] <= 8'h10 ;
			data[73059] <= 8'h10 ;
			data[73060] <= 8'h10 ;
			data[73061] <= 8'h10 ;
			data[73062] <= 8'h10 ;
			data[73063] <= 8'h10 ;
			data[73064] <= 8'h10 ;
			data[73065] <= 8'h10 ;
			data[73066] <= 8'h10 ;
			data[73067] <= 8'h10 ;
			data[73068] <= 8'h10 ;
			data[73069] <= 8'h10 ;
			data[73070] <= 8'h10 ;
			data[73071] <= 8'h10 ;
			data[73072] <= 8'h10 ;
			data[73073] <= 8'h10 ;
			data[73074] <= 8'h10 ;
			data[73075] <= 8'h10 ;
			data[73076] <= 8'h10 ;
			data[73077] <= 8'h10 ;
			data[73078] <= 8'h10 ;
			data[73079] <= 8'h10 ;
			data[73080] <= 8'h10 ;
			data[73081] <= 8'h10 ;
			data[73082] <= 8'h10 ;
			data[73083] <= 8'h10 ;
			data[73084] <= 8'h10 ;
			data[73085] <= 8'h10 ;
			data[73086] <= 8'h10 ;
			data[73087] <= 8'h10 ;
			data[73088] <= 8'h10 ;
			data[73089] <= 8'h10 ;
			data[73090] <= 8'h10 ;
			data[73091] <= 8'h10 ;
			data[73092] <= 8'h10 ;
			data[73093] <= 8'h10 ;
			data[73094] <= 8'h10 ;
			data[73095] <= 8'h10 ;
			data[73096] <= 8'h10 ;
			data[73097] <= 8'h10 ;
			data[73098] <= 8'h10 ;
			data[73099] <= 8'h10 ;
			data[73100] <= 8'h10 ;
			data[73101] <= 8'h10 ;
			data[73102] <= 8'h10 ;
			data[73103] <= 8'h10 ;
			data[73104] <= 8'h10 ;
			data[73105] <= 8'h10 ;
			data[73106] <= 8'h10 ;
			data[73107] <= 8'h10 ;
			data[73108] <= 8'h10 ;
			data[73109] <= 8'h10 ;
			data[73110] <= 8'h10 ;
			data[73111] <= 8'h10 ;
			data[73112] <= 8'h10 ;
			data[73113] <= 8'h10 ;
			data[73114] <= 8'h10 ;
			data[73115] <= 8'h10 ;
			data[73116] <= 8'h10 ;
			data[73117] <= 8'h10 ;
			data[73118] <= 8'h10 ;
			data[73119] <= 8'h10 ;
			data[73120] <= 8'h10 ;
			data[73121] <= 8'h10 ;
			data[73122] <= 8'h10 ;
			data[73123] <= 8'h10 ;
			data[73124] <= 8'h10 ;
			data[73125] <= 8'h10 ;
			data[73126] <= 8'h10 ;
			data[73127] <= 8'h10 ;
			data[73128] <= 8'h10 ;
			data[73129] <= 8'h10 ;
			data[73130] <= 8'h10 ;
			data[73131] <= 8'h10 ;
			data[73132] <= 8'h10 ;
			data[73133] <= 8'h10 ;
			data[73134] <= 8'h10 ;
			data[73135] <= 8'h10 ;
			data[73136] <= 8'h10 ;
			data[73137] <= 8'h10 ;
			data[73138] <= 8'h10 ;
			data[73139] <= 8'h10 ;
			data[73140] <= 8'h10 ;
			data[73141] <= 8'h10 ;
			data[73142] <= 8'h10 ;
			data[73143] <= 8'h10 ;
			data[73144] <= 8'h10 ;
			data[73145] <= 8'h10 ;
			data[73146] <= 8'h10 ;
			data[73147] <= 8'h10 ;
			data[73148] <= 8'h10 ;
			data[73149] <= 8'h10 ;
			data[73150] <= 8'h10 ;
			data[73151] <= 8'h10 ;
			data[73152] <= 8'h10 ;
			data[73153] <= 8'h10 ;
			data[73154] <= 8'h10 ;
			data[73155] <= 8'h10 ;
			data[73156] <= 8'h10 ;
			data[73157] <= 8'h10 ;
			data[73158] <= 8'h10 ;
			data[73159] <= 8'h10 ;
			data[73160] <= 8'h10 ;
			data[73161] <= 8'h10 ;
			data[73162] <= 8'h10 ;
			data[73163] <= 8'h10 ;
			data[73164] <= 8'h10 ;
			data[73165] <= 8'h10 ;
			data[73166] <= 8'h10 ;
			data[73167] <= 8'h10 ;
			data[73168] <= 8'h10 ;
			data[73169] <= 8'h10 ;
			data[73170] <= 8'h10 ;
			data[73171] <= 8'h10 ;
			data[73172] <= 8'h10 ;
			data[73173] <= 8'h10 ;
			data[73174] <= 8'h10 ;
			data[73175] <= 8'h10 ;
			data[73176] <= 8'h10 ;
			data[73177] <= 8'h10 ;
			data[73178] <= 8'h10 ;
			data[73179] <= 8'h10 ;
			data[73180] <= 8'h10 ;
			data[73181] <= 8'h10 ;
			data[73182] <= 8'h10 ;
			data[73183] <= 8'h10 ;
			data[73184] <= 8'h10 ;
			data[73185] <= 8'h10 ;
			data[73186] <= 8'h10 ;
			data[73187] <= 8'h10 ;
			data[73188] <= 8'h10 ;
			data[73189] <= 8'h10 ;
			data[73190] <= 8'h10 ;
			data[73191] <= 8'h10 ;
			data[73192] <= 8'h10 ;
			data[73193] <= 8'h10 ;
			data[73194] <= 8'h10 ;
			data[73195] <= 8'h10 ;
			data[73196] <= 8'h10 ;
			data[73197] <= 8'h10 ;
			data[73198] <= 8'h10 ;
			data[73199] <= 8'h10 ;
			data[73200] <= 8'h10 ;
			data[73201] <= 8'h10 ;
			data[73202] <= 8'h10 ;
			data[73203] <= 8'h10 ;
			data[73204] <= 8'h10 ;
			data[73205] <= 8'h10 ;
			data[73206] <= 8'h10 ;
			data[73207] <= 8'h10 ;
			data[73208] <= 8'h10 ;
			data[73209] <= 8'h10 ;
			data[73210] <= 8'h10 ;
			data[73211] <= 8'h10 ;
			data[73212] <= 8'h10 ;
			data[73213] <= 8'h10 ;
			data[73214] <= 8'h10 ;
			data[73215] <= 8'h10 ;
			data[73216] <= 8'h10 ;
			data[73217] <= 8'h10 ;
			data[73218] <= 8'h10 ;
			data[73219] <= 8'h10 ;
			data[73220] <= 8'h10 ;
			data[73221] <= 8'h10 ;
			data[73222] <= 8'h10 ;
			data[73223] <= 8'h10 ;
			data[73224] <= 8'h10 ;
			data[73225] <= 8'h10 ;
			data[73226] <= 8'h10 ;
			data[73227] <= 8'h10 ;
			data[73228] <= 8'h10 ;
			data[73229] <= 8'h10 ;
			data[73230] <= 8'h10 ;
			data[73231] <= 8'h10 ;
			data[73232] <= 8'h10 ;
			data[73233] <= 8'h10 ;
			data[73234] <= 8'h10 ;
			data[73235] <= 8'h10 ;
			data[73236] <= 8'h10 ;
			data[73237] <= 8'h10 ;
			data[73238] <= 8'h10 ;
			data[73239] <= 8'h10 ;
			data[73240] <= 8'h10 ;
			data[73241] <= 8'h10 ;
			data[73242] <= 8'h10 ;
			data[73243] <= 8'h10 ;
			data[73244] <= 8'h10 ;
			data[73245] <= 8'h10 ;
			data[73246] <= 8'h10 ;
			data[73247] <= 8'h10 ;
			data[73248] <= 8'h10 ;
			data[73249] <= 8'h10 ;
			data[73250] <= 8'h10 ;
			data[73251] <= 8'h10 ;
			data[73252] <= 8'h10 ;
			data[73253] <= 8'h10 ;
			data[73254] <= 8'h10 ;
			data[73255] <= 8'h10 ;
			data[73256] <= 8'h10 ;
			data[73257] <= 8'h10 ;
			data[73258] <= 8'h10 ;
			data[73259] <= 8'h10 ;
			data[73260] <= 8'h10 ;
			data[73261] <= 8'h10 ;
			data[73262] <= 8'h10 ;
			data[73263] <= 8'h10 ;
			data[73264] <= 8'h10 ;
			data[73265] <= 8'h10 ;
			data[73266] <= 8'h10 ;
			data[73267] <= 8'h10 ;
			data[73268] <= 8'h10 ;
			data[73269] <= 8'h10 ;
			data[73270] <= 8'h10 ;
			data[73271] <= 8'h10 ;
			data[73272] <= 8'h10 ;
			data[73273] <= 8'h10 ;
			data[73274] <= 8'h10 ;
			data[73275] <= 8'h10 ;
			data[73276] <= 8'h10 ;
			data[73277] <= 8'h10 ;
			data[73278] <= 8'h10 ;
			data[73279] <= 8'h10 ;
			data[73280] <= 8'h10 ;
			data[73281] <= 8'h10 ;
			data[73282] <= 8'h10 ;
			data[73283] <= 8'h10 ;
			data[73284] <= 8'h10 ;
			data[73285] <= 8'h10 ;
			data[73286] <= 8'h10 ;
			data[73287] <= 8'h10 ;
			data[73288] <= 8'h10 ;
			data[73289] <= 8'h10 ;
			data[73290] <= 8'h10 ;
			data[73291] <= 8'h10 ;
			data[73292] <= 8'h10 ;
			data[73293] <= 8'h10 ;
			data[73294] <= 8'h10 ;
			data[73295] <= 8'h10 ;
			data[73296] <= 8'h10 ;
			data[73297] <= 8'h10 ;
			data[73298] <= 8'h10 ;
			data[73299] <= 8'h10 ;
			data[73300] <= 8'h10 ;
			data[73301] <= 8'h10 ;
			data[73302] <= 8'h10 ;
			data[73303] <= 8'h10 ;
			data[73304] <= 8'h10 ;
			data[73305] <= 8'h10 ;
			data[73306] <= 8'h10 ;
			data[73307] <= 8'h10 ;
			data[73308] <= 8'h10 ;
			data[73309] <= 8'h10 ;
			data[73310] <= 8'h10 ;
			data[73311] <= 8'h10 ;
			data[73312] <= 8'h10 ;
			data[73313] <= 8'h10 ;
			data[73314] <= 8'h10 ;
			data[73315] <= 8'h10 ;
			data[73316] <= 8'h10 ;
			data[73317] <= 8'h10 ;
			data[73318] <= 8'h10 ;
			data[73319] <= 8'h10 ;
			data[73320] <= 8'h10 ;
			data[73321] <= 8'h10 ;
			data[73322] <= 8'h10 ;
			data[73323] <= 8'h10 ;
			data[73324] <= 8'h10 ;
			data[73325] <= 8'h10 ;
			data[73326] <= 8'h10 ;
			data[73327] <= 8'h10 ;
			data[73328] <= 8'h10 ;
			data[73329] <= 8'h10 ;
			data[73330] <= 8'h10 ;
			data[73331] <= 8'h10 ;
			data[73332] <= 8'h10 ;
			data[73333] <= 8'h10 ;
			data[73334] <= 8'h10 ;
			data[73335] <= 8'h10 ;
			data[73336] <= 8'h10 ;
			data[73337] <= 8'h10 ;
			data[73338] <= 8'h10 ;
			data[73339] <= 8'h10 ;
			data[73340] <= 8'h10 ;
			data[73341] <= 8'h10 ;
			data[73342] <= 8'h10 ;
			data[73343] <= 8'h10 ;
			data[73344] <= 8'h10 ;
			data[73345] <= 8'h10 ;
			data[73346] <= 8'h10 ;
			data[73347] <= 8'h10 ;
			data[73348] <= 8'h10 ;
			data[73349] <= 8'h10 ;
			data[73350] <= 8'h10 ;
			data[73351] <= 8'h10 ;
			data[73352] <= 8'h10 ;
			data[73353] <= 8'h10 ;
			data[73354] <= 8'h10 ;
			data[73355] <= 8'h10 ;
			data[73356] <= 8'h10 ;
			data[73357] <= 8'h10 ;
			data[73358] <= 8'h10 ;
			data[73359] <= 8'h10 ;
			data[73360] <= 8'h10 ;
			data[73361] <= 8'h10 ;
			data[73362] <= 8'h10 ;
			data[73363] <= 8'h10 ;
			data[73364] <= 8'h10 ;
			data[73365] <= 8'h10 ;
			data[73366] <= 8'h10 ;
			data[73367] <= 8'h10 ;
			data[73368] <= 8'h10 ;
			data[73369] <= 8'h10 ;
			data[73370] <= 8'h10 ;
			data[73371] <= 8'h10 ;
			data[73372] <= 8'h10 ;
			data[73373] <= 8'h10 ;
			data[73374] <= 8'h10 ;
			data[73375] <= 8'h10 ;
			data[73376] <= 8'h10 ;
			data[73377] <= 8'h10 ;
			data[73378] <= 8'h10 ;
			data[73379] <= 8'h10 ;
			data[73380] <= 8'h10 ;
			data[73381] <= 8'h10 ;
			data[73382] <= 8'h10 ;
			data[73383] <= 8'h10 ;
			data[73384] <= 8'h10 ;
			data[73385] <= 8'h10 ;
			data[73386] <= 8'h10 ;
			data[73387] <= 8'h10 ;
			data[73388] <= 8'h10 ;
			data[73389] <= 8'h10 ;
			data[73390] <= 8'h10 ;
			data[73391] <= 8'h10 ;
			data[73392] <= 8'h10 ;
			data[73393] <= 8'h10 ;
			data[73394] <= 8'h10 ;
			data[73395] <= 8'h10 ;
			data[73396] <= 8'h10 ;
			data[73397] <= 8'h10 ;
			data[73398] <= 8'h10 ;
			data[73399] <= 8'h10 ;
			data[73400] <= 8'h10 ;
			data[73401] <= 8'h10 ;
			data[73402] <= 8'h10 ;
			data[73403] <= 8'h10 ;
			data[73404] <= 8'h10 ;
			data[73405] <= 8'h10 ;
			data[73406] <= 8'h10 ;
			data[73407] <= 8'h10 ;
			data[73408] <= 8'h10 ;
			data[73409] <= 8'h10 ;
			data[73410] <= 8'h10 ;
			data[73411] <= 8'h10 ;
			data[73412] <= 8'h10 ;
			data[73413] <= 8'h10 ;
			data[73414] <= 8'h10 ;
			data[73415] <= 8'h10 ;
			data[73416] <= 8'h10 ;
			data[73417] <= 8'h10 ;
			data[73418] <= 8'h10 ;
			data[73419] <= 8'h10 ;
			data[73420] <= 8'h10 ;
			data[73421] <= 8'h10 ;
			data[73422] <= 8'h10 ;
			data[73423] <= 8'h10 ;
			data[73424] <= 8'h10 ;
			data[73425] <= 8'h10 ;
			data[73426] <= 8'h10 ;
			data[73427] <= 8'h10 ;
			data[73428] <= 8'h10 ;
			data[73429] <= 8'h10 ;
			data[73430] <= 8'h10 ;
			data[73431] <= 8'h10 ;
			data[73432] <= 8'h10 ;
			data[73433] <= 8'h10 ;
			data[73434] <= 8'h10 ;
			data[73435] <= 8'h10 ;
			data[73436] <= 8'h10 ;
			data[73437] <= 8'h10 ;
			data[73438] <= 8'h10 ;
			data[73439] <= 8'h10 ;
			data[73440] <= 8'h10 ;
			data[73441] <= 8'h10 ;
			data[73442] <= 8'h10 ;
			data[73443] <= 8'h10 ;
			data[73444] <= 8'h10 ;
			data[73445] <= 8'h10 ;
			data[73446] <= 8'h10 ;
			data[73447] <= 8'h10 ;
			data[73448] <= 8'h10 ;
			data[73449] <= 8'h10 ;
			data[73450] <= 8'h10 ;
			data[73451] <= 8'h10 ;
			data[73452] <= 8'h10 ;
			data[73453] <= 8'h10 ;
			data[73454] <= 8'h10 ;
			data[73455] <= 8'h10 ;
			data[73456] <= 8'h10 ;
			data[73457] <= 8'h10 ;
			data[73458] <= 8'h10 ;
			data[73459] <= 8'h10 ;
			data[73460] <= 8'h10 ;
			data[73461] <= 8'h10 ;
			data[73462] <= 8'h10 ;
			data[73463] <= 8'h10 ;
			data[73464] <= 8'h10 ;
			data[73465] <= 8'h10 ;
			data[73466] <= 8'h10 ;
			data[73467] <= 8'h10 ;
			data[73468] <= 8'h10 ;
			data[73469] <= 8'h10 ;
			data[73470] <= 8'h10 ;
			data[73471] <= 8'h10 ;
			data[73472] <= 8'h10 ;
			data[73473] <= 8'h10 ;
			data[73474] <= 8'h10 ;
			data[73475] <= 8'h10 ;
			data[73476] <= 8'h10 ;
			data[73477] <= 8'h10 ;
			data[73478] <= 8'h10 ;
			data[73479] <= 8'h10 ;
			data[73480] <= 8'h10 ;
			data[73481] <= 8'h10 ;
			data[73482] <= 8'h10 ;
			data[73483] <= 8'h10 ;
			data[73484] <= 8'h10 ;
			data[73485] <= 8'h10 ;
			data[73486] <= 8'h10 ;
			data[73487] <= 8'h10 ;
			data[73488] <= 8'h10 ;
			data[73489] <= 8'h10 ;
			data[73490] <= 8'h10 ;
			data[73491] <= 8'h10 ;
			data[73492] <= 8'h10 ;
			data[73493] <= 8'h10 ;
			data[73494] <= 8'h10 ;
			data[73495] <= 8'h10 ;
			data[73496] <= 8'h10 ;
			data[73497] <= 8'h10 ;
			data[73498] <= 8'h10 ;
			data[73499] <= 8'h10 ;
			data[73500] <= 8'h10 ;
			data[73501] <= 8'h10 ;
			data[73502] <= 8'h10 ;
			data[73503] <= 8'h10 ;
			data[73504] <= 8'h10 ;
			data[73505] <= 8'h10 ;
			data[73506] <= 8'h10 ;
			data[73507] <= 8'h10 ;
			data[73508] <= 8'h10 ;
			data[73509] <= 8'h10 ;
			data[73510] <= 8'h10 ;
			data[73511] <= 8'h10 ;
			data[73512] <= 8'h10 ;
			data[73513] <= 8'h10 ;
			data[73514] <= 8'h10 ;
			data[73515] <= 8'h10 ;
			data[73516] <= 8'h10 ;
			data[73517] <= 8'h10 ;
			data[73518] <= 8'h10 ;
			data[73519] <= 8'h10 ;
			data[73520] <= 8'h10 ;
			data[73521] <= 8'h10 ;
			data[73522] <= 8'h10 ;
			data[73523] <= 8'h10 ;
			data[73524] <= 8'h10 ;
			data[73525] <= 8'h10 ;
			data[73526] <= 8'h10 ;
			data[73527] <= 8'h10 ;
			data[73528] <= 8'h10 ;
			data[73529] <= 8'h10 ;
			data[73530] <= 8'h10 ;
			data[73531] <= 8'h10 ;
			data[73532] <= 8'h10 ;
			data[73533] <= 8'h10 ;
			data[73534] <= 8'h10 ;
			data[73535] <= 8'h10 ;
			data[73536] <= 8'h10 ;
			data[73537] <= 8'h10 ;
			data[73538] <= 8'h10 ;
			data[73539] <= 8'h10 ;
			data[73540] <= 8'h10 ;
			data[73541] <= 8'h10 ;
			data[73542] <= 8'h10 ;
			data[73543] <= 8'h10 ;
			data[73544] <= 8'h10 ;
			data[73545] <= 8'h10 ;
			data[73546] <= 8'h10 ;
			data[73547] <= 8'h10 ;
			data[73548] <= 8'h10 ;
			data[73549] <= 8'h10 ;
			data[73550] <= 8'h10 ;
			data[73551] <= 8'h10 ;
			data[73552] <= 8'h10 ;
			data[73553] <= 8'h10 ;
			data[73554] <= 8'h10 ;
			data[73555] <= 8'h10 ;
			data[73556] <= 8'h10 ;
			data[73557] <= 8'h10 ;
			data[73558] <= 8'h10 ;
			data[73559] <= 8'h10 ;
			data[73560] <= 8'h10 ;
			data[73561] <= 8'h10 ;
			data[73562] <= 8'h10 ;
			data[73563] <= 8'h10 ;
			data[73564] <= 8'h10 ;
			data[73565] <= 8'h10 ;
			data[73566] <= 8'h10 ;
			data[73567] <= 8'h10 ;
			data[73568] <= 8'h10 ;
			data[73569] <= 8'h10 ;
			data[73570] <= 8'h10 ;
			data[73571] <= 8'h10 ;
			data[73572] <= 8'h10 ;
			data[73573] <= 8'h10 ;
			data[73574] <= 8'h10 ;
			data[73575] <= 8'h10 ;
			data[73576] <= 8'h10 ;
			data[73577] <= 8'h10 ;
			data[73578] <= 8'h10 ;
			data[73579] <= 8'h10 ;
			data[73580] <= 8'h10 ;
			data[73581] <= 8'h10 ;
			data[73582] <= 8'h10 ;
			data[73583] <= 8'h10 ;
			data[73584] <= 8'h10 ;
			data[73585] <= 8'h10 ;
			data[73586] <= 8'h10 ;
			data[73587] <= 8'h10 ;
			data[73588] <= 8'h10 ;
			data[73589] <= 8'h10 ;
			data[73590] <= 8'h10 ;
			data[73591] <= 8'h10 ;
			data[73592] <= 8'h10 ;
			data[73593] <= 8'h10 ;
			data[73594] <= 8'h10 ;
			data[73595] <= 8'h10 ;
			data[73596] <= 8'h10 ;
			data[73597] <= 8'h10 ;
			data[73598] <= 8'h10 ;
			data[73599] <= 8'h10 ;
			data[73600] <= 8'h10 ;
			data[73601] <= 8'h10 ;
			data[73602] <= 8'h10 ;
			data[73603] <= 8'h10 ;
			data[73604] <= 8'h10 ;
			data[73605] <= 8'h10 ;
			data[73606] <= 8'h10 ;
			data[73607] <= 8'h10 ;
			data[73608] <= 8'h10 ;
			data[73609] <= 8'h10 ;
			data[73610] <= 8'h10 ;
			data[73611] <= 8'h10 ;
			data[73612] <= 8'h10 ;
			data[73613] <= 8'h10 ;
			data[73614] <= 8'h10 ;
			data[73615] <= 8'h10 ;
			data[73616] <= 8'h10 ;
			data[73617] <= 8'h10 ;
			data[73618] <= 8'h10 ;
			data[73619] <= 8'h10 ;
			data[73620] <= 8'h10 ;
			data[73621] <= 8'h10 ;
			data[73622] <= 8'h10 ;
			data[73623] <= 8'h10 ;
			data[73624] <= 8'h10 ;
			data[73625] <= 8'h10 ;
			data[73626] <= 8'h10 ;
			data[73627] <= 8'h10 ;
			data[73628] <= 8'h10 ;
			data[73629] <= 8'h10 ;
			data[73630] <= 8'h10 ;
			data[73631] <= 8'h10 ;
			data[73632] <= 8'h10 ;
			data[73633] <= 8'h10 ;
			data[73634] <= 8'h10 ;
			data[73635] <= 8'h10 ;
			data[73636] <= 8'h10 ;
			data[73637] <= 8'h10 ;
			data[73638] <= 8'h10 ;
			data[73639] <= 8'h10 ;
			data[73640] <= 8'h10 ;
			data[73641] <= 8'h10 ;
			data[73642] <= 8'h10 ;
			data[73643] <= 8'h10 ;
			data[73644] <= 8'h10 ;
			data[73645] <= 8'h10 ;
			data[73646] <= 8'h10 ;
			data[73647] <= 8'h10 ;
			data[73648] <= 8'h10 ;
			data[73649] <= 8'h10 ;
			data[73650] <= 8'h10 ;
			data[73651] <= 8'h10 ;
			data[73652] <= 8'h10 ;
			data[73653] <= 8'h10 ;
			data[73654] <= 8'h10 ;
			data[73655] <= 8'h10 ;
			data[73656] <= 8'h10 ;
			data[73657] <= 8'h10 ;
			data[73658] <= 8'h10 ;
			data[73659] <= 8'h10 ;
			data[73660] <= 8'h10 ;
			data[73661] <= 8'h10 ;
			data[73662] <= 8'h10 ;
			data[73663] <= 8'h10 ;
			data[73664] <= 8'h10 ;
			data[73665] <= 8'h10 ;
			data[73666] <= 8'h10 ;
			data[73667] <= 8'h10 ;
			data[73668] <= 8'h10 ;
			data[73669] <= 8'h10 ;
			data[73670] <= 8'h10 ;
			data[73671] <= 8'h10 ;
			data[73672] <= 8'h10 ;
			data[73673] <= 8'h10 ;
			data[73674] <= 8'h10 ;
			data[73675] <= 8'h10 ;
			data[73676] <= 8'h10 ;
			data[73677] <= 8'h10 ;
			data[73678] <= 8'h10 ;
			data[73679] <= 8'h10 ;
			data[73680] <= 8'h10 ;
			data[73681] <= 8'h10 ;
			data[73682] <= 8'h10 ;
			data[73683] <= 8'h10 ;
			data[73684] <= 8'h10 ;
			data[73685] <= 8'h10 ;
			data[73686] <= 8'h10 ;
			data[73687] <= 8'h10 ;
			data[73688] <= 8'h10 ;
			data[73689] <= 8'h10 ;
			data[73690] <= 8'h10 ;
			data[73691] <= 8'h10 ;
			data[73692] <= 8'h10 ;
			data[73693] <= 8'h10 ;
			data[73694] <= 8'h10 ;
			data[73695] <= 8'h10 ;
			data[73696] <= 8'h10 ;
			data[73697] <= 8'h10 ;
			data[73698] <= 8'h10 ;
			data[73699] <= 8'h10 ;
			data[73700] <= 8'h10 ;
			data[73701] <= 8'h10 ;
			data[73702] <= 8'h10 ;
			data[73703] <= 8'h10 ;
			data[73704] <= 8'h10 ;
			data[73705] <= 8'h10 ;
			data[73706] <= 8'h10 ;
			data[73707] <= 8'h10 ;
			data[73708] <= 8'h10 ;
			data[73709] <= 8'h10 ;
			data[73710] <= 8'h10 ;
			data[73711] <= 8'h10 ;
			data[73712] <= 8'h10 ;
			data[73713] <= 8'h10 ;
			data[73714] <= 8'h10 ;
			data[73715] <= 8'h10 ;
			data[73716] <= 8'h10 ;
			data[73717] <= 8'h10 ;
			data[73718] <= 8'h10 ;
			data[73719] <= 8'h10 ;
			data[73720] <= 8'h10 ;
			data[73721] <= 8'h10 ;
			data[73722] <= 8'h10 ;
			data[73723] <= 8'h10 ;
			data[73724] <= 8'h10 ;
			data[73725] <= 8'h10 ;
			data[73726] <= 8'h10 ;
			data[73727] <= 8'h10 ;
			data[73728] <= 8'h10 ;
			data[73729] <= 8'h10 ;
			data[73730] <= 8'h10 ;
			data[73731] <= 8'h10 ;
			data[73732] <= 8'h10 ;
			data[73733] <= 8'h10 ;
			data[73734] <= 8'h10 ;
			data[73735] <= 8'h10 ;
			data[73736] <= 8'h10 ;
			data[73737] <= 8'h10 ;
			data[73738] <= 8'h10 ;
			data[73739] <= 8'h10 ;
			data[73740] <= 8'h10 ;
			data[73741] <= 8'h10 ;
			data[73742] <= 8'h10 ;
			data[73743] <= 8'h10 ;
			data[73744] <= 8'h10 ;
			data[73745] <= 8'h10 ;
			data[73746] <= 8'h10 ;
			data[73747] <= 8'h10 ;
			data[73748] <= 8'h10 ;
			data[73749] <= 8'h10 ;
			data[73750] <= 8'h10 ;
			data[73751] <= 8'h10 ;
			data[73752] <= 8'h10 ;
			data[73753] <= 8'h10 ;
			data[73754] <= 8'h10 ;
			data[73755] <= 8'h10 ;
			data[73756] <= 8'h10 ;
			data[73757] <= 8'h10 ;
			data[73758] <= 8'h10 ;
			data[73759] <= 8'h10 ;
			data[73760] <= 8'h10 ;
			data[73761] <= 8'h10 ;
			data[73762] <= 8'h10 ;
			data[73763] <= 8'h10 ;
			data[73764] <= 8'h10 ;
			data[73765] <= 8'h10 ;
			data[73766] <= 8'h10 ;
			data[73767] <= 8'h10 ;
			data[73768] <= 8'h10 ;
			data[73769] <= 8'h10 ;
			data[73770] <= 8'h10 ;
			data[73771] <= 8'h10 ;
			data[73772] <= 8'h10 ;
			data[73773] <= 8'h10 ;
			data[73774] <= 8'h10 ;
			data[73775] <= 8'h10 ;
			data[73776] <= 8'h10 ;
			data[73777] <= 8'h10 ;
			data[73778] <= 8'h10 ;
			data[73779] <= 8'h10 ;
			data[73780] <= 8'h10 ;
			data[73781] <= 8'h10 ;
			data[73782] <= 8'h10 ;
			data[73783] <= 8'h10 ;
			data[73784] <= 8'h10 ;
			data[73785] <= 8'h10 ;
			data[73786] <= 8'h10 ;
			data[73787] <= 8'h10 ;
			data[73788] <= 8'h10 ;
			data[73789] <= 8'h10 ;
			data[73790] <= 8'h10 ;
			data[73791] <= 8'h10 ;
			data[73792] <= 8'h10 ;
			data[73793] <= 8'h10 ;
			data[73794] <= 8'h10 ;
			data[73795] <= 8'h10 ;
			data[73796] <= 8'h10 ;
			data[73797] <= 8'h10 ;
			data[73798] <= 8'h10 ;
			data[73799] <= 8'h10 ;
			data[73800] <= 8'h10 ;
			data[73801] <= 8'h10 ;
			data[73802] <= 8'h10 ;
			data[73803] <= 8'h10 ;
			data[73804] <= 8'h10 ;
			data[73805] <= 8'h10 ;
			data[73806] <= 8'h10 ;
			data[73807] <= 8'h10 ;
			data[73808] <= 8'h10 ;
			data[73809] <= 8'h10 ;
			data[73810] <= 8'h10 ;
			data[73811] <= 8'h10 ;
			data[73812] <= 8'h10 ;
			data[73813] <= 8'h10 ;
			data[73814] <= 8'h10 ;
			data[73815] <= 8'h10 ;
			data[73816] <= 8'h10 ;
			data[73817] <= 8'h10 ;
			data[73818] <= 8'h10 ;
			data[73819] <= 8'h10 ;
			data[73820] <= 8'h10 ;
			data[73821] <= 8'h10 ;
			data[73822] <= 8'h10 ;
			data[73823] <= 8'h10 ;
			data[73824] <= 8'h10 ;
			data[73825] <= 8'h10 ;
			data[73826] <= 8'h10 ;
			data[73827] <= 8'h10 ;
			data[73828] <= 8'h10 ;
			data[73829] <= 8'h10 ;
			data[73830] <= 8'h10 ;
			data[73831] <= 8'h10 ;
			data[73832] <= 8'h10 ;
			data[73833] <= 8'h10 ;
			data[73834] <= 8'h10 ;
			data[73835] <= 8'h10 ;
			data[73836] <= 8'h10 ;
			data[73837] <= 8'h10 ;
			data[73838] <= 8'h10 ;
			data[73839] <= 8'h10 ;
			data[73840] <= 8'h10 ;
			data[73841] <= 8'h10 ;
			data[73842] <= 8'h10 ;
			data[73843] <= 8'h10 ;
			data[73844] <= 8'h10 ;
			data[73845] <= 8'h10 ;
			data[73846] <= 8'h10 ;
			data[73847] <= 8'h10 ;
			data[73848] <= 8'h10 ;
			data[73849] <= 8'h10 ;
			data[73850] <= 8'h10 ;
			data[73851] <= 8'h10 ;
			data[73852] <= 8'h10 ;
			data[73853] <= 8'h10 ;
			data[73854] <= 8'h10 ;
			data[73855] <= 8'h10 ;
			data[73856] <= 8'h10 ;
			data[73857] <= 8'h10 ;
			data[73858] <= 8'h10 ;
			data[73859] <= 8'h10 ;
			data[73860] <= 8'h10 ;
			data[73861] <= 8'h10 ;
			data[73862] <= 8'h10 ;
			data[73863] <= 8'h10 ;
			data[73864] <= 8'h10 ;
			data[73865] <= 8'h10 ;
			data[73866] <= 8'h10 ;
			data[73867] <= 8'h10 ;
			data[73868] <= 8'h10 ;
			data[73869] <= 8'h10 ;
			data[73870] <= 8'h10 ;
			data[73871] <= 8'h10 ;
			data[73872] <= 8'h10 ;
			data[73873] <= 8'h10 ;
			data[73874] <= 8'h10 ;
			data[73875] <= 8'h10 ;
			data[73876] <= 8'h10 ;
			data[73877] <= 8'h10 ;
			data[73878] <= 8'h10 ;
			data[73879] <= 8'h10 ;
			data[73880] <= 8'h10 ;
			data[73881] <= 8'h10 ;
			data[73882] <= 8'h10 ;
			data[73883] <= 8'h10 ;
			data[73884] <= 8'h10 ;
			data[73885] <= 8'h10 ;
			data[73886] <= 8'h10 ;
			data[73887] <= 8'h10 ;
			data[73888] <= 8'h10 ;
			data[73889] <= 8'h10 ;
			data[73890] <= 8'h10 ;
			data[73891] <= 8'h10 ;
			data[73892] <= 8'h10 ;
			data[73893] <= 8'h10 ;
			data[73894] <= 8'h10 ;
			data[73895] <= 8'h10 ;
			data[73896] <= 8'h10 ;
			data[73897] <= 8'h10 ;
			data[73898] <= 8'h10 ;
			data[73899] <= 8'h10 ;
			data[73900] <= 8'h10 ;
			data[73901] <= 8'h10 ;
			data[73902] <= 8'h10 ;
			data[73903] <= 8'h10 ;
			data[73904] <= 8'h10 ;
			data[73905] <= 8'h10 ;
			data[73906] <= 8'h10 ;
			data[73907] <= 8'h10 ;
			data[73908] <= 8'h10 ;
			data[73909] <= 8'h10 ;
			data[73910] <= 8'h10 ;
			data[73911] <= 8'h10 ;
			data[73912] <= 8'h10 ;
			data[73913] <= 8'h10 ;
			data[73914] <= 8'h10 ;
			data[73915] <= 8'h10 ;
			data[73916] <= 8'h10 ;
			data[73917] <= 8'h10 ;
			data[73918] <= 8'h10 ;
			data[73919] <= 8'h10 ;
			data[73920] <= 8'h10 ;
			data[73921] <= 8'h10 ;
			data[73922] <= 8'h10 ;
			data[73923] <= 8'h10 ;
			data[73924] <= 8'h10 ;
			data[73925] <= 8'h10 ;
			data[73926] <= 8'h10 ;
			data[73927] <= 8'h10 ;
			data[73928] <= 8'h10 ;
			data[73929] <= 8'h10 ;
			data[73930] <= 8'h10 ;
			data[73931] <= 8'h10 ;
			data[73932] <= 8'h10 ;
			data[73933] <= 8'h10 ;
			data[73934] <= 8'h10 ;
			data[73935] <= 8'h10 ;
			data[73936] <= 8'h10 ;
			data[73937] <= 8'h10 ;
			data[73938] <= 8'h10 ;
			data[73939] <= 8'h10 ;
			data[73940] <= 8'h10 ;
			data[73941] <= 8'h10 ;
			data[73942] <= 8'h10 ;
			data[73943] <= 8'h10 ;
			data[73944] <= 8'h10 ;
			data[73945] <= 8'h10 ;
			data[73946] <= 8'h10 ;
			data[73947] <= 8'h10 ;
			data[73948] <= 8'h10 ;
			data[73949] <= 8'h10 ;
			data[73950] <= 8'h10 ;
			data[73951] <= 8'h10 ;
			data[73952] <= 8'h10 ;
			data[73953] <= 8'h10 ;
			data[73954] <= 8'h10 ;
			data[73955] <= 8'h10 ;
			data[73956] <= 8'h10 ;
			data[73957] <= 8'h10 ;
			data[73958] <= 8'h10 ;
			data[73959] <= 8'h10 ;
			data[73960] <= 8'h10 ;
			data[73961] <= 8'h10 ;
			data[73962] <= 8'h10 ;
			data[73963] <= 8'h10 ;
			data[73964] <= 8'h10 ;
			data[73965] <= 8'h10 ;
			data[73966] <= 8'h10 ;
			data[73967] <= 8'h10 ;
			data[73968] <= 8'h10 ;
			data[73969] <= 8'h10 ;
			data[73970] <= 8'h10 ;
			data[73971] <= 8'h10 ;
			data[73972] <= 8'h10 ;
			data[73973] <= 8'h10 ;
			data[73974] <= 8'h10 ;
			data[73975] <= 8'h10 ;
			data[73976] <= 8'h10 ;
			data[73977] <= 8'h10 ;
			data[73978] <= 8'h10 ;
			data[73979] <= 8'h10 ;
			data[73980] <= 8'h10 ;
			data[73981] <= 8'h10 ;
			data[73982] <= 8'h10 ;
			data[73983] <= 8'h10 ;
			data[73984] <= 8'h10 ;
			data[73985] <= 8'h10 ;
			data[73986] <= 8'h10 ;
			data[73987] <= 8'h10 ;
			data[73988] <= 8'h10 ;
			data[73989] <= 8'h10 ;
			data[73990] <= 8'h10 ;
			data[73991] <= 8'h10 ;
			data[73992] <= 8'h10 ;
			data[73993] <= 8'h10 ;
			data[73994] <= 8'h10 ;
			data[73995] <= 8'h10 ;
			data[73996] <= 8'h10 ;
			data[73997] <= 8'h10 ;
			data[73998] <= 8'h10 ;
			data[73999] <= 8'h10 ;
			data[74000] <= 8'h10 ;
			data[74001] <= 8'h10 ;
			data[74002] <= 8'h10 ;
			data[74003] <= 8'h10 ;
			data[74004] <= 8'h10 ;
			data[74005] <= 8'h10 ;
			data[74006] <= 8'h10 ;
			data[74007] <= 8'h10 ;
			data[74008] <= 8'h10 ;
			data[74009] <= 8'h10 ;
			data[74010] <= 8'h10 ;
			data[74011] <= 8'h10 ;
			data[74012] <= 8'h10 ;
			data[74013] <= 8'h10 ;
			data[74014] <= 8'h10 ;
			data[74015] <= 8'h10 ;
			data[74016] <= 8'h10 ;
			data[74017] <= 8'h10 ;
			data[74018] <= 8'h10 ;
			data[74019] <= 8'h10 ;
			data[74020] <= 8'h10 ;
			data[74021] <= 8'h10 ;
			data[74022] <= 8'h10 ;
			data[74023] <= 8'h10 ;
			data[74024] <= 8'h10 ;
			data[74025] <= 8'h10 ;
			data[74026] <= 8'h10 ;
			data[74027] <= 8'h10 ;
			data[74028] <= 8'h10 ;
			data[74029] <= 8'h10 ;
			data[74030] <= 8'h10 ;
			data[74031] <= 8'h10 ;
			data[74032] <= 8'h10 ;
			data[74033] <= 8'h10 ;
			data[74034] <= 8'h10 ;
			data[74035] <= 8'h10 ;
			data[74036] <= 8'h10 ;
			data[74037] <= 8'h10 ;
			data[74038] <= 8'h10 ;
			data[74039] <= 8'h10 ;
			data[74040] <= 8'h10 ;
			data[74041] <= 8'h10 ;
			data[74042] <= 8'h10 ;
			data[74043] <= 8'h10 ;
			data[74044] <= 8'h10 ;
			data[74045] <= 8'h10 ;
			data[74046] <= 8'h10 ;
			data[74047] <= 8'h10 ;
			data[74048] <= 8'h10 ;
			data[74049] <= 8'h10 ;
			data[74050] <= 8'h10 ;
			data[74051] <= 8'h10 ;
			data[74052] <= 8'h10 ;
			data[74053] <= 8'h10 ;
			data[74054] <= 8'h10 ;
			data[74055] <= 8'h10 ;
			data[74056] <= 8'h10 ;
			data[74057] <= 8'h10 ;
			data[74058] <= 8'h10 ;
			data[74059] <= 8'h10 ;
			data[74060] <= 8'h10 ;
			data[74061] <= 8'h10 ;
			data[74062] <= 8'h10 ;
			data[74063] <= 8'h10 ;
			data[74064] <= 8'h10 ;
			data[74065] <= 8'h10 ;
			data[74066] <= 8'h10 ;
			data[74067] <= 8'h10 ;
			data[74068] <= 8'h10 ;
			data[74069] <= 8'h10 ;
			data[74070] <= 8'h10 ;
			data[74071] <= 8'h10 ;
			data[74072] <= 8'h10 ;
			data[74073] <= 8'h10 ;
			data[74074] <= 8'h10 ;
			data[74075] <= 8'h10 ;
			data[74076] <= 8'h10 ;
			data[74077] <= 8'h10 ;
			data[74078] <= 8'h10 ;
			data[74079] <= 8'h10 ;
			data[74080] <= 8'h10 ;
			data[74081] <= 8'h10 ;
			data[74082] <= 8'h10 ;
			data[74083] <= 8'h10 ;
			data[74084] <= 8'h10 ;
			data[74085] <= 8'h10 ;
			data[74086] <= 8'h10 ;
			data[74087] <= 8'h10 ;
			data[74088] <= 8'h10 ;
			data[74089] <= 8'h10 ;
			data[74090] <= 8'h10 ;
			data[74091] <= 8'h10 ;
			data[74092] <= 8'h10 ;
			data[74093] <= 8'h10 ;
			data[74094] <= 8'h10 ;
			data[74095] <= 8'h10 ;
			data[74096] <= 8'h10 ;
			data[74097] <= 8'h10 ;
			data[74098] <= 8'h10 ;
			data[74099] <= 8'h10 ;
			data[74100] <= 8'h10 ;
			data[74101] <= 8'h10 ;
			data[74102] <= 8'h10 ;
			data[74103] <= 8'h10 ;
			data[74104] <= 8'h10 ;
			data[74105] <= 8'h10 ;
			data[74106] <= 8'h10 ;
			data[74107] <= 8'h10 ;
			data[74108] <= 8'h10 ;
			data[74109] <= 8'h10 ;
			data[74110] <= 8'h10 ;
			data[74111] <= 8'h10 ;
			data[74112] <= 8'h10 ;
			data[74113] <= 8'h10 ;
			data[74114] <= 8'h10 ;
			data[74115] <= 8'h10 ;
			data[74116] <= 8'h10 ;
			data[74117] <= 8'h10 ;
			data[74118] <= 8'h10 ;
			data[74119] <= 8'h10 ;
			data[74120] <= 8'h10 ;
			data[74121] <= 8'h10 ;
			data[74122] <= 8'h10 ;
			data[74123] <= 8'h10 ;
			data[74124] <= 8'h10 ;
			data[74125] <= 8'h10 ;
			data[74126] <= 8'h10 ;
			data[74127] <= 8'h10 ;
			data[74128] <= 8'h10 ;
			data[74129] <= 8'h10 ;
			data[74130] <= 8'h10 ;
			data[74131] <= 8'h10 ;
			data[74132] <= 8'h10 ;
			data[74133] <= 8'h10 ;
			data[74134] <= 8'h10 ;
			data[74135] <= 8'h10 ;
			data[74136] <= 8'h10 ;
			data[74137] <= 8'h10 ;
			data[74138] <= 8'h10 ;
			data[74139] <= 8'h10 ;
			data[74140] <= 8'h10 ;
			data[74141] <= 8'h10 ;
			data[74142] <= 8'h10 ;
			data[74143] <= 8'h10 ;
			data[74144] <= 8'h10 ;
			data[74145] <= 8'h10 ;
			data[74146] <= 8'h10 ;
			data[74147] <= 8'h10 ;
			data[74148] <= 8'h10 ;
			data[74149] <= 8'h10 ;
			data[74150] <= 8'h10 ;
			data[74151] <= 8'h10 ;
			data[74152] <= 8'h10 ;
			data[74153] <= 8'h10 ;
			data[74154] <= 8'h10 ;
			data[74155] <= 8'h10 ;
			data[74156] <= 8'h10 ;
			data[74157] <= 8'h10 ;
			data[74158] <= 8'h10 ;
			data[74159] <= 8'h10 ;
			data[74160] <= 8'h10 ;
			data[74161] <= 8'h10 ;
			data[74162] <= 8'h10 ;
			data[74163] <= 8'h10 ;
			data[74164] <= 8'h10 ;
			data[74165] <= 8'h10 ;
			data[74166] <= 8'h10 ;
			data[74167] <= 8'h10 ;
			data[74168] <= 8'h10 ;
			data[74169] <= 8'h10 ;
			data[74170] <= 8'h10 ;
			data[74171] <= 8'h10 ;
			data[74172] <= 8'h10 ;
			data[74173] <= 8'h10 ;
			data[74174] <= 8'h10 ;
			data[74175] <= 8'h10 ;
			data[74176] <= 8'h10 ;
			data[74177] <= 8'h10 ;
			data[74178] <= 8'h10 ;
			data[74179] <= 8'h10 ;
			data[74180] <= 8'h10 ;
			data[74181] <= 8'h10 ;
			data[74182] <= 8'h10 ;
			data[74183] <= 8'h10 ;
			data[74184] <= 8'h10 ;
			data[74185] <= 8'h10 ;
			data[74186] <= 8'h10 ;
			data[74187] <= 8'h10 ;
			data[74188] <= 8'h10 ;
			data[74189] <= 8'h10 ;
			data[74190] <= 8'h10 ;
			data[74191] <= 8'h10 ;
			data[74192] <= 8'h10 ;
			data[74193] <= 8'h10 ;
			data[74194] <= 8'h10 ;
			data[74195] <= 8'h10 ;
			data[74196] <= 8'h10 ;
			data[74197] <= 8'h10 ;
			data[74198] <= 8'h10 ;
			data[74199] <= 8'h10 ;
			data[74200] <= 8'h10 ;
			data[74201] <= 8'h10 ;
			data[74202] <= 8'h10 ;
			data[74203] <= 8'h10 ;
			data[74204] <= 8'h10 ;
			data[74205] <= 8'h10 ;
			data[74206] <= 8'h10 ;
			data[74207] <= 8'h10 ;
			data[74208] <= 8'h10 ;
			data[74209] <= 8'h10 ;
			data[74210] <= 8'h10 ;
			data[74211] <= 8'h10 ;
			data[74212] <= 8'h10 ;
			data[74213] <= 8'h10 ;
			data[74214] <= 8'h10 ;
			data[74215] <= 8'h10 ;
			data[74216] <= 8'h10 ;
			data[74217] <= 8'h10 ;
			data[74218] <= 8'h10 ;
			data[74219] <= 8'h10 ;
			data[74220] <= 8'h10 ;
			data[74221] <= 8'h10 ;
			data[74222] <= 8'h10 ;
			data[74223] <= 8'h10 ;
			data[74224] <= 8'h10 ;
			data[74225] <= 8'h10 ;
			data[74226] <= 8'h10 ;
			data[74227] <= 8'h10 ;
			data[74228] <= 8'h10 ;
			data[74229] <= 8'h10 ;
			data[74230] <= 8'h10 ;
			data[74231] <= 8'h10 ;
			data[74232] <= 8'h10 ;
			data[74233] <= 8'h10 ;
			data[74234] <= 8'h10 ;
			data[74235] <= 8'h10 ;
			data[74236] <= 8'h10 ;
			data[74237] <= 8'h10 ;
			data[74238] <= 8'h10 ;
			data[74239] <= 8'h10 ;
			data[74240] <= 8'h10 ;
			data[74241] <= 8'h10 ;
			data[74242] <= 8'h10 ;
			data[74243] <= 8'h10 ;
			data[74244] <= 8'h10 ;
			data[74245] <= 8'h10 ;
			data[74246] <= 8'h10 ;
			data[74247] <= 8'h10 ;
			data[74248] <= 8'h10 ;
			data[74249] <= 8'h10 ;
			data[74250] <= 8'h10 ;
			data[74251] <= 8'h10 ;
			data[74252] <= 8'h10 ;
			data[74253] <= 8'h10 ;
			data[74254] <= 8'h10 ;
			data[74255] <= 8'h10 ;
			data[74256] <= 8'h10 ;
			data[74257] <= 8'h10 ;
			data[74258] <= 8'h10 ;
			data[74259] <= 8'h10 ;
			data[74260] <= 8'h10 ;
			data[74261] <= 8'h10 ;
			data[74262] <= 8'h10 ;
			data[74263] <= 8'h10 ;
			data[74264] <= 8'h10 ;
			data[74265] <= 8'h10 ;
			data[74266] <= 8'h10 ;
			data[74267] <= 8'h10 ;
			data[74268] <= 8'h10 ;
			data[74269] <= 8'h10 ;
			data[74270] <= 8'h10 ;
			data[74271] <= 8'h10 ;
			data[74272] <= 8'h10 ;
			data[74273] <= 8'h10 ;
			data[74274] <= 8'h10 ;
			data[74275] <= 8'h10 ;
			data[74276] <= 8'h10 ;
			data[74277] <= 8'h10 ;
			data[74278] <= 8'h10 ;
			data[74279] <= 8'h10 ;
			data[74280] <= 8'h10 ;
			data[74281] <= 8'h10 ;
			data[74282] <= 8'h10 ;
			data[74283] <= 8'h10 ;
			data[74284] <= 8'h10 ;
			data[74285] <= 8'h10 ;
			data[74286] <= 8'h10 ;
			data[74287] <= 8'h10 ;
			data[74288] <= 8'h10 ;
			data[74289] <= 8'h10 ;
			data[74290] <= 8'h10 ;
			data[74291] <= 8'h10 ;
			data[74292] <= 8'h10 ;
			data[74293] <= 8'h10 ;
			data[74294] <= 8'h10 ;
			data[74295] <= 8'h10 ;
			data[74296] <= 8'h10 ;
			data[74297] <= 8'h10 ;
			data[74298] <= 8'h10 ;
			data[74299] <= 8'h10 ;
			data[74300] <= 8'h10 ;
			data[74301] <= 8'h10 ;
			data[74302] <= 8'h10 ;
			data[74303] <= 8'h10 ;
			data[74304] <= 8'h10 ;
			data[74305] <= 8'h10 ;
			data[74306] <= 8'h10 ;
			data[74307] <= 8'h10 ;
			data[74308] <= 8'h10 ;
			data[74309] <= 8'h10 ;
			data[74310] <= 8'h10 ;
			data[74311] <= 8'h10 ;
			data[74312] <= 8'h10 ;
			data[74313] <= 8'h10 ;
			data[74314] <= 8'h10 ;
			data[74315] <= 8'h10 ;
			data[74316] <= 8'h10 ;
			data[74317] <= 8'h10 ;
			data[74318] <= 8'h10 ;
			data[74319] <= 8'h10 ;
			data[74320] <= 8'h10 ;
			data[74321] <= 8'h10 ;
			data[74322] <= 8'h10 ;
			data[74323] <= 8'h10 ;
			data[74324] <= 8'h10 ;
			data[74325] <= 8'h10 ;
			data[74326] <= 8'h10 ;
			data[74327] <= 8'h10 ;
			data[74328] <= 8'h10 ;
			data[74329] <= 8'h10 ;
			data[74330] <= 8'h10 ;
			data[74331] <= 8'h10 ;
			data[74332] <= 8'h10 ;
			data[74333] <= 8'h10 ;
			data[74334] <= 8'h10 ;
			data[74335] <= 8'h10 ;
			data[74336] <= 8'h10 ;
			data[74337] <= 8'h10 ;
			data[74338] <= 8'h10 ;
			data[74339] <= 8'h10 ;
			data[74340] <= 8'h10 ;
			data[74341] <= 8'h10 ;
			data[74342] <= 8'h10 ;
			data[74343] <= 8'h10 ;
			data[74344] <= 8'h10 ;
			data[74345] <= 8'h10 ;
			data[74346] <= 8'h10 ;
			data[74347] <= 8'h10 ;
			data[74348] <= 8'h10 ;
			data[74349] <= 8'h10 ;
			data[74350] <= 8'h10 ;
			data[74351] <= 8'h10 ;
			data[74352] <= 8'h10 ;
			data[74353] <= 8'h10 ;
			data[74354] <= 8'h10 ;
			data[74355] <= 8'h10 ;
			data[74356] <= 8'h10 ;
			data[74357] <= 8'h10 ;
			data[74358] <= 8'h10 ;
			data[74359] <= 8'h10 ;
			data[74360] <= 8'h10 ;
			data[74361] <= 8'h10 ;
			data[74362] <= 8'h10 ;
			data[74363] <= 8'h10 ;
			data[74364] <= 8'h10 ;
			data[74365] <= 8'h10 ;
			data[74366] <= 8'h10 ;
			data[74367] <= 8'h10 ;
			data[74368] <= 8'h10 ;
			data[74369] <= 8'h10 ;
			data[74370] <= 8'h10 ;
			data[74371] <= 8'h10 ;
			data[74372] <= 8'h10 ;
			data[74373] <= 8'h10 ;
			data[74374] <= 8'h10 ;
			data[74375] <= 8'h10 ;
			data[74376] <= 8'h10 ;
			data[74377] <= 8'h10 ;
			data[74378] <= 8'h10 ;
			data[74379] <= 8'h10 ;
			data[74380] <= 8'h10 ;
			data[74381] <= 8'h10 ;
			data[74382] <= 8'h10 ;
			data[74383] <= 8'h10 ;
			data[74384] <= 8'h10 ;
			data[74385] <= 8'h10 ;
			data[74386] <= 8'h10 ;
			data[74387] <= 8'h10 ;
			data[74388] <= 8'h10 ;
			data[74389] <= 8'h10 ;
			data[74390] <= 8'h10 ;
			data[74391] <= 8'h10 ;
			data[74392] <= 8'h10 ;
			data[74393] <= 8'h10 ;
			data[74394] <= 8'h10 ;
			data[74395] <= 8'h10 ;
			data[74396] <= 8'h10 ;
			data[74397] <= 8'h10 ;
			data[74398] <= 8'h10 ;
			data[74399] <= 8'h10 ;
			data[74400] <= 8'h10 ;
			data[74401] <= 8'h10 ;
			data[74402] <= 8'h10 ;
			data[74403] <= 8'h10 ;
			data[74404] <= 8'h10 ;
			data[74405] <= 8'h10 ;
			data[74406] <= 8'h10 ;
			data[74407] <= 8'h10 ;
			data[74408] <= 8'h10 ;
			data[74409] <= 8'h10 ;
			data[74410] <= 8'h10 ;
			data[74411] <= 8'h10 ;
			data[74412] <= 8'h10 ;
			data[74413] <= 8'h10 ;
			data[74414] <= 8'h10 ;
			data[74415] <= 8'h10 ;
			data[74416] <= 8'h10 ;
			data[74417] <= 8'h10 ;
			data[74418] <= 8'h10 ;
			data[74419] <= 8'h10 ;
			data[74420] <= 8'h10 ;
			data[74421] <= 8'h10 ;
			data[74422] <= 8'h10 ;
			data[74423] <= 8'h10 ;
			data[74424] <= 8'h10 ;
			data[74425] <= 8'h10 ;
			data[74426] <= 8'h10 ;
			data[74427] <= 8'h10 ;
			data[74428] <= 8'h10 ;
			data[74429] <= 8'h10 ;
			data[74430] <= 8'h10 ;
			data[74431] <= 8'h10 ;
			data[74432] <= 8'h10 ;
			data[74433] <= 8'h10 ;
			data[74434] <= 8'h10 ;
			data[74435] <= 8'h10 ;
			data[74436] <= 8'h10 ;
			data[74437] <= 8'h10 ;
			data[74438] <= 8'h10 ;
			data[74439] <= 8'h10 ;
			data[74440] <= 8'h10 ;
			data[74441] <= 8'h10 ;
			data[74442] <= 8'h10 ;
			data[74443] <= 8'h10 ;
			data[74444] <= 8'h10 ;
			data[74445] <= 8'h10 ;
			data[74446] <= 8'h10 ;
			data[74447] <= 8'h10 ;
			data[74448] <= 8'h10 ;
			data[74449] <= 8'h10 ;
			data[74450] <= 8'h10 ;
			data[74451] <= 8'h10 ;
			data[74452] <= 8'h10 ;
			data[74453] <= 8'h10 ;
			data[74454] <= 8'h10 ;
			data[74455] <= 8'h10 ;
			data[74456] <= 8'h10 ;
			data[74457] <= 8'h10 ;
			data[74458] <= 8'h10 ;
			data[74459] <= 8'h10 ;
			data[74460] <= 8'h10 ;
			data[74461] <= 8'h10 ;
			data[74462] <= 8'h10 ;
			data[74463] <= 8'h10 ;
			data[74464] <= 8'h10 ;
			data[74465] <= 8'h10 ;
			data[74466] <= 8'h10 ;
			data[74467] <= 8'h10 ;
			data[74468] <= 8'h10 ;
			data[74469] <= 8'h10 ;
			data[74470] <= 8'h10 ;
			data[74471] <= 8'h10 ;
			data[74472] <= 8'h10 ;
			data[74473] <= 8'h10 ;
			data[74474] <= 8'h10 ;
			data[74475] <= 8'h10 ;
			data[74476] <= 8'h10 ;
			data[74477] <= 8'h10 ;
			data[74478] <= 8'h10 ;
			data[74479] <= 8'h10 ;
			data[74480] <= 8'h10 ;
			data[74481] <= 8'h10 ;
			data[74482] <= 8'h10 ;
			data[74483] <= 8'h10 ;
			data[74484] <= 8'h10 ;
			data[74485] <= 8'h10 ;
			data[74486] <= 8'h10 ;
			data[74487] <= 8'h10 ;
			data[74488] <= 8'h10 ;
			data[74489] <= 8'h10 ;
			data[74490] <= 8'h10 ;
			data[74491] <= 8'h10 ;
			data[74492] <= 8'h10 ;
			data[74493] <= 8'h10 ;
			data[74494] <= 8'h10 ;
			data[74495] <= 8'h10 ;
			data[74496] <= 8'h10 ;
			data[74497] <= 8'h10 ;
			data[74498] <= 8'h10 ;
			data[74499] <= 8'h10 ;
			data[74500] <= 8'h10 ;
			data[74501] <= 8'h10 ;
			data[74502] <= 8'h10 ;
			data[74503] <= 8'h10 ;
			data[74504] <= 8'h10 ;
			data[74505] <= 8'h10 ;
			data[74506] <= 8'h10 ;
			data[74507] <= 8'h10 ;
			data[74508] <= 8'h10 ;
			data[74509] <= 8'h10 ;
			data[74510] <= 8'h10 ;
			data[74511] <= 8'h10 ;
			data[74512] <= 8'h10 ;
			data[74513] <= 8'h10 ;
			data[74514] <= 8'h10 ;
			data[74515] <= 8'h10 ;
			data[74516] <= 8'h10 ;
			data[74517] <= 8'h10 ;
			data[74518] <= 8'h10 ;
			data[74519] <= 8'h10 ;
			data[74520] <= 8'h10 ;
			data[74521] <= 8'h10 ;
			data[74522] <= 8'h10 ;
			data[74523] <= 8'h10 ;
			data[74524] <= 8'h10 ;
			data[74525] <= 8'h10 ;
			data[74526] <= 8'h10 ;
			data[74527] <= 8'h10 ;
			data[74528] <= 8'h10 ;
			data[74529] <= 8'h10 ;
			data[74530] <= 8'h10 ;
			data[74531] <= 8'h10 ;
			data[74532] <= 8'h10 ;
			data[74533] <= 8'h10 ;
			data[74534] <= 8'h10 ;
			data[74535] <= 8'h10 ;
			data[74536] <= 8'h10 ;
			data[74537] <= 8'h10 ;
			data[74538] <= 8'h10 ;
			data[74539] <= 8'h10 ;
			data[74540] <= 8'h10 ;
			data[74541] <= 8'h10 ;
			data[74542] <= 8'h10 ;
			data[74543] <= 8'h10 ;
			data[74544] <= 8'h10 ;
			data[74545] <= 8'h10 ;
			data[74546] <= 8'h10 ;
			data[74547] <= 8'h10 ;
			data[74548] <= 8'h10 ;
			data[74549] <= 8'h10 ;
			data[74550] <= 8'h10 ;
			data[74551] <= 8'h10 ;
			data[74552] <= 8'h10 ;
			data[74553] <= 8'h10 ;
			data[74554] <= 8'h10 ;
			data[74555] <= 8'h10 ;
			data[74556] <= 8'h10 ;
			data[74557] <= 8'h10 ;
			data[74558] <= 8'h10 ;
			data[74559] <= 8'h10 ;
			data[74560] <= 8'h10 ;
			data[74561] <= 8'h10 ;
			data[74562] <= 8'h10 ;
			data[74563] <= 8'h10 ;
			data[74564] <= 8'h10 ;
			data[74565] <= 8'h10 ;
			data[74566] <= 8'h10 ;
			data[74567] <= 8'h10 ;
			data[74568] <= 8'h10 ;
			data[74569] <= 8'h10 ;
			data[74570] <= 8'h10 ;
			data[74571] <= 8'h10 ;
			data[74572] <= 8'h10 ;
			data[74573] <= 8'h10 ;
			data[74574] <= 8'h10 ;
			data[74575] <= 8'h10 ;
			data[74576] <= 8'h10 ;
			data[74577] <= 8'h10 ;
			data[74578] <= 8'h10 ;
			data[74579] <= 8'h10 ;
			data[74580] <= 8'h10 ;
			data[74581] <= 8'h10 ;
			data[74582] <= 8'h10 ;
			data[74583] <= 8'h10 ;
			data[74584] <= 8'h10 ;
			data[74585] <= 8'h10 ;
			data[74586] <= 8'h10 ;
			data[74587] <= 8'h10 ;
			data[74588] <= 8'h10 ;
			data[74589] <= 8'h10 ;
			data[74590] <= 8'h10 ;
			data[74591] <= 8'h10 ;
			data[74592] <= 8'h10 ;
			data[74593] <= 8'h10 ;
			data[74594] <= 8'h10 ;
			data[74595] <= 8'h10 ;
			data[74596] <= 8'h10 ;
			data[74597] <= 8'h10 ;
			data[74598] <= 8'h10 ;
			data[74599] <= 8'h10 ;
			data[74600] <= 8'h10 ;
			data[74601] <= 8'h10 ;
			data[74602] <= 8'h10 ;
			data[74603] <= 8'h10 ;
			data[74604] <= 8'h10 ;
			data[74605] <= 8'h10 ;
			data[74606] <= 8'h10 ;
			data[74607] <= 8'h10 ;
			data[74608] <= 8'h10 ;
			data[74609] <= 8'h10 ;
			data[74610] <= 8'h10 ;
			data[74611] <= 8'h10 ;
			data[74612] <= 8'h10 ;
			data[74613] <= 8'h10 ;
			data[74614] <= 8'h10 ;
			data[74615] <= 8'h10 ;
			data[74616] <= 8'h10 ;
			data[74617] <= 8'h10 ;
			data[74618] <= 8'h10 ;
			data[74619] <= 8'h10 ;
			data[74620] <= 8'h10 ;
			data[74621] <= 8'h10 ;
			data[74622] <= 8'h10 ;
			data[74623] <= 8'h10 ;
			data[74624] <= 8'h10 ;
			data[74625] <= 8'h10 ;
			data[74626] <= 8'h10 ;
			data[74627] <= 8'h10 ;
			data[74628] <= 8'h10 ;
			data[74629] <= 8'h10 ;
			data[74630] <= 8'h10 ;
			data[74631] <= 8'h10 ;
			data[74632] <= 8'h10 ;
			data[74633] <= 8'h10 ;
			data[74634] <= 8'h10 ;
			data[74635] <= 8'h10 ;
			data[74636] <= 8'h10 ;
			data[74637] <= 8'h10 ;
			data[74638] <= 8'h10 ;
			data[74639] <= 8'h10 ;
			data[74640] <= 8'h10 ;
			data[74641] <= 8'h10 ;
			data[74642] <= 8'h10 ;
			data[74643] <= 8'h10 ;
			data[74644] <= 8'h10 ;
			data[74645] <= 8'h10 ;
			data[74646] <= 8'h10 ;
			data[74647] <= 8'h10 ;
			data[74648] <= 8'h10 ;
			data[74649] <= 8'h10 ;
			data[74650] <= 8'h10 ;
			data[74651] <= 8'h10 ;
			data[74652] <= 8'h10 ;
			data[74653] <= 8'h10 ;
			data[74654] <= 8'h10 ;
			data[74655] <= 8'h10 ;
			data[74656] <= 8'h10 ;
			data[74657] <= 8'h10 ;
			data[74658] <= 8'h10 ;
			data[74659] <= 8'h10 ;
			data[74660] <= 8'h10 ;
			data[74661] <= 8'h10 ;
			data[74662] <= 8'h10 ;
			data[74663] <= 8'h10 ;
			data[74664] <= 8'h10 ;
			data[74665] <= 8'h10 ;
			data[74666] <= 8'h10 ;
			data[74667] <= 8'h10 ;
			data[74668] <= 8'h10 ;
			data[74669] <= 8'h10 ;
			data[74670] <= 8'h10 ;
			data[74671] <= 8'h10 ;
			data[74672] <= 8'h10 ;
			data[74673] <= 8'h10 ;
			data[74674] <= 8'h10 ;
			data[74675] <= 8'h10 ;
			data[74676] <= 8'h10 ;
			data[74677] <= 8'h10 ;
			data[74678] <= 8'h10 ;
			data[74679] <= 8'h10 ;
			data[74680] <= 8'h10 ;
			data[74681] <= 8'h10 ;
			data[74682] <= 8'h10 ;
			data[74683] <= 8'h10 ;
			data[74684] <= 8'h10 ;
			data[74685] <= 8'h10 ;
			data[74686] <= 8'h10 ;
			data[74687] <= 8'h10 ;
			data[74688] <= 8'h10 ;
			data[74689] <= 8'h10 ;
			data[74690] <= 8'h10 ;
			data[74691] <= 8'h10 ;
			data[74692] <= 8'h10 ;
			data[74693] <= 8'h10 ;
			data[74694] <= 8'h10 ;
			data[74695] <= 8'h10 ;
			data[74696] <= 8'h10 ;
			data[74697] <= 8'h10 ;
			data[74698] <= 8'h10 ;
			data[74699] <= 8'h10 ;
			data[74700] <= 8'h10 ;
			data[74701] <= 8'h10 ;
			data[74702] <= 8'h10 ;
			data[74703] <= 8'h10 ;
			data[74704] <= 8'h10 ;
			data[74705] <= 8'h10 ;
			data[74706] <= 8'h10 ;
			data[74707] <= 8'h10 ;
			data[74708] <= 8'h10 ;
			data[74709] <= 8'h10 ;
			data[74710] <= 8'h10 ;
			data[74711] <= 8'h10 ;
			data[74712] <= 8'h10 ;
			data[74713] <= 8'h10 ;
			data[74714] <= 8'h10 ;
			data[74715] <= 8'h10 ;
			data[74716] <= 8'h10 ;
			data[74717] <= 8'h10 ;
			data[74718] <= 8'h10 ;
			data[74719] <= 8'h10 ;
			data[74720] <= 8'h10 ;
			data[74721] <= 8'h10 ;
			data[74722] <= 8'h10 ;
			data[74723] <= 8'h10 ;
			data[74724] <= 8'h10 ;
			data[74725] <= 8'h10 ;
			data[74726] <= 8'h10 ;
			data[74727] <= 8'h10 ;
			data[74728] <= 8'h10 ;
			data[74729] <= 8'h10 ;
			data[74730] <= 8'h10 ;
			data[74731] <= 8'h10 ;
			data[74732] <= 8'h10 ;
			data[74733] <= 8'h10 ;
			data[74734] <= 8'h10 ;
			data[74735] <= 8'h10 ;
			data[74736] <= 8'h10 ;
			data[74737] <= 8'h10 ;
			data[74738] <= 8'h10 ;
			data[74739] <= 8'h10 ;
			data[74740] <= 8'h10 ;
			data[74741] <= 8'h10 ;
			data[74742] <= 8'h10 ;
			data[74743] <= 8'h10 ;
			data[74744] <= 8'h10 ;
			data[74745] <= 8'h10 ;
			data[74746] <= 8'h10 ;
			data[74747] <= 8'h10 ;
			data[74748] <= 8'h10 ;
			data[74749] <= 8'h10 ;
			data[74750] <= 8'h10 ;
			data[74751] <= 8'h10 ;
			data[74752] <= 8'h10 ;
			data[74753] <= 8'h10 ;
			data[74754] <= 8'h10 ;
			data[74755] <= 8'h10 ;
			data[74756] <= 8'h10 ;
			data[74757] <= 8'h10 ;
			data[74758] <= 8'h10 ;
			data[74759] <= 8'h10 ;
			data[74760] <= 8'h10 ;
			data[74761] <= 8'h10 ;
			data[74762] <= 8'h10 ;
			data[74763] <= 8'h10 ;
			data[74764] <= 8'h10 ;
			data[74765] <= 8'h10 ;
			data[74766] <= 8'h10 ;
			data[74767] <= 8'h10 ;
			data[74768] <= 8'h10 ;
			data[74769] <= 8'h10 ;
			data[74770] <= 8'h10 ;
			data[74771] <= 8'h10 ;
			data[74772] <= 8'h10 ;
			data[74773] <= 8'h10 ;
			data[74774] <= 8'h10 ;
			data[74775] <= 8'h10 ;
			data[74776] <= 8'h10 ;
			data[74777] <= 8'h10 ;
			data[74778] <= 8'h10 ;
			data[74779] <= 8'h10 ;
			data[74780] <= 8'h10 ;
			data[74781] <= 8'h10 ;
			data[74782] <= 8'h10 ;
			data[74783] <= 8'h10 ;
			data[74784] <= 8'h10 ;
			data[74785] <= 8'h10 ;
			data[74786] <= 8'h10 ;
			data[74787] <= 8'h10 ;
			data[74788] <= 8'h10 ;
			data[74789] <= 8'h10 ;
			data[74790] <= 8'h10 ;
			data[74791] <= 8'h10 ;
			data[74792] <= 8'h10 ;
			data[74793] <= 8'h10 ;
			data[74794] <= 8'h10 ;
			data[74795] <= 8'h10 ;
			data[74796] <= 8'h10 ;
			data[74797] <= 8'h10 ;
			data[74798] <= 8'h10 ;
			data[74799] <= 8'h10 ;
			data[74800] <= 8'h10 ;
			data[74801] <= 8'h10 ;
			data[74802] <= 8'h10 ;
			data[74803] <= 8'h10 ;
			data[74804] <= 8'h10 ;
			data[74805] <= 8'h10 ;
			data[74806] <= 8'h10 ;
			data[74807] <= 8'h10 ;
			data[74808] <= 8'h10 ;
			data[74809] <= 8'h10 ;
			data[74810] <= 8'h10 ;
			data[74811] <= 8'h10 ;
			data[74812] <= 8'h10 ;
			data[74813] <= 8'h10 ;
			data[74814] <= 8'h10 ;
			data[74815] <= 8'h10 ;
			data[74816] <= 8'h10 ;
			data[74817] <= 8'h10 ;
			data[74818] <= 8'h10 ;
			data[74819] <= 8'h10 ;
			data[74820] <= 8'h10 ;
			data[74821] <= 8'h10 ;
			data[74822] <= 8'h10 ;
			data[74823] <= 8'h10 ;
			data[74824] <= 8'h10 ;
			data[74825] <= 8'h10 ;
			data[74826] <= 8'h10 ;
			data[74827] <= 8'h10 ;
			data[74828] <= 8'h10 ;
			data[74829] <= 8'h10 ;
			data[74830] <= 8'h10 ;
			data[74831] <= 8'h10 ;
			data[74832] <= 8'h10 ;
			data[74833] <= 8'h10 ;
			data[74834] <= 8'h10 ;
			data[74835] <= 8'h10 ;
			data[74836] <= 8'h10 ;
			data[74837] <= 8'h10 ;
			data[74838] <= 8'h10 ;
			data[74839] <= 8'h10 ;
			data[74840] <= 8'h10 ;
			data[74841] <= 8'h10 ;
			data[74842] <= 8'h10 ;
			data[74843] <= 8'h10 ;
			data[74844] <= 8'h10 ;
			data[74845] <= 8'h10 ;
			data[74846] <= 8'h10 ;
			data[74847] <= 8'h10 ;
			data[74848] <= 8'h10 ;
			data[74849] <= 8'h10 ;
			data[74850] <= 8'h10 ;
			data[74851] <= 8'h10 ;
			data[74852] <= 8'h10 ;
			data[74853] <= 8'h10 ;
			data[74854] <= 8'h10 ;
			data[74855] <= 8'h10 ;
			data[74856] <= 8'h10 ;
			data[74857] <= 8'h10 ;
			data[74858] <= 8'h10 ;
			data[74859] <= 8'h10 ;
			data[74860] <= 8'h10 ;
			data[74861] <= 8'h10 ;
			data[74862] <= 8'h10 ;
			data[74863] <= 8'h10 ;
			data[74864] <= 8'h10 ;
			data[74865] <= 8'h10 ;
			data[74866] <= 8'h10 ;
			data[74867] <= 8'h10 ;
			data[74868] <= 8'h10 ;
			data[74869] <= 8'h10 ;
			data[74870] <= 8'h10 ;
			data[74871] <= 8'h10 ;
			data[74872] <= 8'h10 ;
			data[74873] <= 8'h10 ;
			data[74874] <= 8'h10 ;
			data[74875] <= 8'h10 ;
			data[74876] <= 8'h10 ;
			data[74877] <= 8'h10 ;
			data[74878] <= 8'h10 ;
			data[74879] <= 8'h10 ;
			data[74880] <= 8'h10 ;
			data[74881] <= 8'h10 ;
			data[74882] <= 8'h10 ;
			data[74883] <= 8'h10 ;
			data[74884] <= 8'h10 ;
			data[74885] <= 8'h10 ;
			data[74886] <= 8'h10 ;
			data[74887] <= 8'h10 ;
			data[74888] <= 8'h10 ;
			data[74889] <= 8'h10 ;
			data[74890] <= 8'h10 ;
			data[74891] <= 8'h10 ;
			data[74892] <= 8'h10 ;
			data[74893] <= 8'h10 ;
			data[74894] <= 8'h10 ;
			data[74895] <= 8'h10 ;
			data[74896] <= 8'h10 ;
			data[74897] <= 8'h10 ;
			data[74898] <= 8'h10 ;
			data[74899] <= 8'h10 ;
			data[74900] <= 8'h10 ;
			data[74901] <= 8'h10 ;
			data[74902] <= 8'h10 ;
			data[74903] <= 8'h10 ;
			data[74904] <= 8'h10 ;
			data[74905] <= 8'h10 ;
			data[74906] <= 8'h10 ;
			data[74907] <= 8'h10 ;
			data[74908] <= 8'h10 ;
			data[74909] <= 8'h10 ;
			data[74910] <= 8'h10 ;
			data[74911] <= 8'h10 ;
			data[74912] <= 8'h10 ;
			data[74913] <= 8'h10 ;
			data[74914] <= 8'h10 ;
			data[74915] <= 8'h10 ;
			data[74916] <= 8'h10 ;
			data[74917] <= 8'h10 ;
			data[74918] <= 8'h10 ;
			data[74919] <= 8'h10 ;
			data[74920] <= 8'h10 ;
			data[74921] <= 8'h10 ;
			data[74922] <= 8'h10 ;
			data[74923] <= 8'h10 ;
			data[74924] <= 8'h10 ;
			data[74925] <= 8'h10 ;
			data[74926] <= 8'h10 ;
			data[74927] <= 8'h10 ;
			data[74928] <= 8'h10 ;
			data[74929] <= 8'h10 ;
			data[74930] <= 8'h10 ;
			data[74931] <= 8'h10 ;
			data[74932] <= 8'h10 ;
			data[74933] <= 8'h10 ;
			data[74934] <= 8'h10 ;
			data[74935] <= 8'h10 ;
			data[74936] <= 8'h10 ;
			data[74937] <= 8'h10 ;
			data[74938] <= 8'h10 ;
			data[74939] <= 8'h10 ;
			data[74940] <= 8'h10 ;
			data[74941] <= 8'h10 ;
			data[74942] <= 8'h10 ;
			data[74943] <= 8'h10 ;
			data[74944] <= 8'h10 ;
			data[74945] <= 8'h10 ;
			data[74946] <= 8'h10 ;
			data[74947] <= 8'h10 ;
			data[74948] <= 8'h10 ;
			data[74949] <= 8'h10 ;
			data[74950] <= 8'h10 ;
			data[74951] <= 8'h10 ;
			data[74952] <= 8'h10 ;
			data[74953] <= 8'h10 ;
			data[74954] <= 8'h10 ;
			data[74955] <= 8'h10 ;
			data[74956] <= 8'h10 ;
			data[74957] <= 8'h10 ;
			data[74958] <= 8'h10 ;
			data[74959] <= 8'h10 ;
			data[74960] <= 8'h10 ;
			data[74961] <= 8'h10 ;
			data[74962] <= 8'h10 ;
			data[74963] <= 8'h10 ;
			data[74964] <= 8'h10 ;
			data[74965] <= 8'h10 ;
			data[74966] <= 8'h10 ;
			data[74967] <= 8'h10 ;
			data[74968] <= 8'h10 ;
			data[74969] <= 8'h10 ;
			data[74970] <= 8'h10 ;
			data[74971] <= 8'h10 ;
			data[74972] <= 8'h10 ;
			data[74973] <= 8'h10 ;
			data[74974] <= 8'h10 ;
			data[74975] <= 8'h10 ;
			data[74976] <= 8'h10 ;
			data[74977] <= 8'h10 ;
			data[74978] <= 8'h10 ;
			data[74979] <= 8'h10 ;
			data[74980] <= 8'h10 ;
			data[74981] <= 8'h10 ;
			data[74982] <= 8'h10 ;
			data[74983] <= 8'h10 ;
			data[74984] <= 8'h10 ;
			data[74985] <= 8'h10 ;
			data[74986] <= 8'h10 ;
			data[74987] <= 8'h10 ;
			data[74988] <= 8'h10 ;
			data[74989] <= 8'h10 ;
			data[74990] <= 8'h10 ;
			data[74991] <= 8'h10 ;
			data[74992] <= 8'h10 ;
			data[74993] <= 8'h10 ;
			data[74994] <= 8'h10 ;
			data[74995] <= 8'h10 ;
			data[74996] <= 8'h10 ;
			data[74997] <= 8'h10 ;
			data[74998] <= 8'h10 ;
			data[74999] <= 8'h10 ;
			data[75000] <= 8'h10 ;
			data[75001] <= 8'h10 ;
			data[75002] <= 8'h10 ;
			data[75003] <= 8'h10 ;
			data[75004] <= 8'h10 ;
			data[75005] <= 8'h10 ;
			data[75006] <= 8'h10 ;
			data[75007] <= 8'h10 ;
			data[75008] <= 8'h10 ;
			data[75009] <= 8'h10 ;
			data[75010] <= 8'h10 ;
			data[75011] <= 8'h10 ;
			data[75012] <= 8'h10 ;
			data[75013] <= 8'h10 ;
			data[75014] <= 8'h10 ;
			data[75015] <= 8'h10 ;
			data[75016] <= 8'h10 ;
			data[75017] <= 8'h10 ;
			data[75018] <= 8'h10 ;
			data[75019] <= 8'h10 ;
			data[75020] <= 8'h10 ;
			data[75021] <= 8'h10 ;
			data[75022] <= 8'h10 ;
			data[75023] <= 8'h10 ;
			data[75024] <= 8'h10 ;
			data[75025] <= 8'h10 ;
			data[75026] <= 8'h10 ;
			data[75027] <= 8'h10 ;
			data[75028] <= 8'h10 ;
			data[75029] <= 8'h10 ;
			data[75030] <= 8'h10 ;
			data[75031] <= 8'h10 ;
			data[75032] <= 8'h10 ;
			data[75033] <= 8'h10 ;
			data[75034] <= 8'h10 ;
			data[75035] <= 8'h10 ;
			data[75036] <= 8'h10 ;
			data[75037] <= 8'h10 ;
			data[75038] <= 8'h10 ;
			data[75039] <= 8'h10 ;
			data[75040] <= 8'h10 ;
			data[75041] <= 8'h10 ;
			data[75042] <= 8'h10 ;
			data[75043] <= 8'h10 ;
			data[75044] <= 8'h10 ;
			data[75045] <= 8'h10 ;
			data[75046] <= 8'h10 ;
			data[75047] <= 8'h10 ;
			data[75048] <= 8'h10 ;
			data[75049] <= 8'h10 ;
			data[75050] <= 8'h10 ;
			data[75051] <= 8'h10 ;
			data[75052] <= 8'h10 ;
			data[75053] <= 8'h10 ;
			data[75054] <= 8'h10 ;
			data[75055] <= 8'h10 ;
			data[75056] <= 8'h10 ;
			data[75057] <= 8'h10 ;
			data[75058] <= 8'h10 ;
			data[75059] <= 8'h10 ;
			data[75060] <= 8'h10 ;
			data[75061] <= 8'h10 ;
			data[75062] <= 8'h10 ;
			data[75063] <= 8'h10 ;
			data[75064] <= 8'h10 ;
			data[75065] <= 8'h10 ;
			data[75066] <= 8'h10 ;
			data[75067] <= 8'h10 ;
			data[75068] <= 8'h10 ;
			data[75069] <= 8'h10 ;
			data[75070] <= 8'h10 ;
			data[75071] <= 8'h10 ;
			data[75072] <= 8'h10 ;
			data[75073] <= 8'h10 ;
			data[75074] <= 8'h10 ;
			data[75075] <= 8'h10 ;
			data[75076] <= 8'h10 ;
			data[75077] <= 8'h10 ;
			data[75078] <= 8'h10 ;
			data[75079] <= 8'h10 ;
			data[75080] <= 8'h10 ;
			data[75081] <= 8'h10 ;
			data[75082] <= 8'h10 ;
			data[75083] <= 8'h10 ;
			data[75084] <= 8'h10 ;
			data[75085] <= 8'h10 ;
			data[75086] <= 8'h10 ;
			data[75087] <= 8'h10 ;
			data[75088] <= 8'h10 ;
			data[75089] <= 8'h10 ;
			data[75090] <= 8'h10 ;
			data[75091] <= 8'h10 ;
			data[75092] <= 8'h10 ;
			data[75093] <= 8'h10 ;
			data[75094] <= 8'h10 ;
			data[75095] <= 8'h10 ;
			data[75096] <= 8'h10 ;
			data[75097] <= 8'h10 ;
			data[75098] <= 8'h10 ;
			data[75099] <= 8'h10 ;
			data[75100] <= 8'h10 ;
			data[75101] <= 8'h10 ;
			data[75102] <= 8'h10 ;
			data[75103] <= 8'h10 ;
			data[75104] <= 8'h10 ;
			data[75105] <= 8'h10 ;
			data[75106] <= 8'h10 ;
			data[75107] <= 8'h10 ;
			data[75108] <= 8'h10 ;
			data[75109] <= 8'h10 ;
			data[75110] <= 8'h10 ;
			data[75111] <= 8'h10 ;
			data[75112] <= 8'h10 ;
			data[75113] <= 8'h10 ;
			data[75114] <= 8'h10 ;
			data[75115] <= 8'h10 ;
			data[75116] <= 8'h10 ;
			data[75117] <= 8'h10 ;
			data[75118] <= 8'h10 ;
			data[75119] <= 8'h10 ;
			data[75120] <= 8'h10 ;
			data[75121] <= 8'h10 ;
			data[75122] <= 8'h10 ;
			data[75123] <= 8'h10 ;
			data[75124] <= 8'h10 ;
			data[75125] <= 8'h10 ;
			data[75126] <= 8'h10 ;
			data[75127] <= 8'h10 ;
			data[75128] <= 8'h10 ;
			data[75129] <= 8'h10 ;
			data[75130] <= 8'h10 ;
			data[75131] <= 8'h10 ;
			data[75132] <= 8'h10 ;
			data[75133] <= 8'h10 ;
			data[75134] <= 8'h10 ;
			data[75135] <= 8'h10 ;
			data[75136] <= 8'h10 ;
			data[75137] <= 8'h10 ;
			data[75138] <= 8'h10 ;
			data[75139] <= 8'h10 ;
			data[75140] <= 8'h10 ;
			data[75141] <= 8'h10 ;
			data[75142] <= 8'h10 ;
			data[75143] <= 8'h10 ;
			data[75144] <= 8'h10 ;
			data[75145] <= 8'h10 ;
			data[75146] <= 8'h10 ;
			data[75147] <= 8'h10 ;
			data[75148] <= 8'h10 ;
			data[75149] <= 8'h10 ;
			data[75150] <= 8'h10 ;
			data[75151] <= 8'h10 ;
			data[75152] <= 8'h10 ;
			data[75153] <= 8'h10 ;
			data[75154] <= 8'h10 ;
			data[75155] <= 8'h10 ;
			data[75156] <= 8'h10 ;
			data[75157] <= 8'h10 ;
			data[75158] <= 8'h10 ;
			data[75159] <= 8'h10 ;
			data[75160] <= 8'h10 ;
			data[75161] <= 8'h10 ;
			data[75162] <= 8'h10 ;
			data[75163] <= 8'h10 ;
			data[75164] <= 8'h10 ;
			data[75165] <= 8'h10 ;
			data[75166] <= 8'h10 ;
			data[75167] <= 8'h10 ;
			data[75168] <= 8'h10 ;
			data[75169] <= 8'h10 ;
			data[75170] <= 8'h10 ;
			data[75171] <= 8'h10 ;
			data[75172] <= 8'h10 ;
			data[75173] <= 8'h10 ;
			data[75174] <= 8'h10 ;
			data[75175] <= 8'h10 ;
			data[75176] <= 8'h10 ;
			data[75177] <= 8'h10 ;
			data[75178] <= 8'h10 ;
			data[75179] <= 8'h10 ;
			data[75180] <= 8'h10 ;
			data[75181] <= 8'h10 ;
			data[75182] <= 8'h10 ;
			data[75183] <= 8'h10 ;
			data[75184] <= 8'h10 ;
			data[75185] <= 8'h10 ;
			data[75186] <= 8'h10 ;
			data[75187] <= 8'h10 ;
			data[75188] <= 8'h10 ;
			data[75189] <= 8'h10 ;
			data[75190] <= 8'h10 ;
			data[75191] <= 8'h10 ;
			data[75192] <= 8'h10 ;
			data[75193] <= 8'h10 ;
			data[75194] <= 8'h10 ;
			data[75195] <= 8'h10 ;
			data[75196] <= 8'h10 ;
			data[75197] <= 8'h10 ;
			data[75198] <= 8'h10 ;
			data[75199] <= 8'h10 ;
			data[75200] <= 8'h10 ;
			data[75201] <= 8'h10 ;
			data[75202] <= 8'h10 ;
			data[75203] <= 8'h10 ;
			data[75204] <= 8'h10 ;
			data[75205] <= 8'h10 ;
			data[75206] <= 8'h10 ;
			data[75207] <= 8'h10 ;
			data[75208] <= 8'h10 ;
			data[75209] <= 8'h10 ;
			data[75210] <= 8'h10 ;
			data[75211] <= 8'h10 ;
			data[75212] <= 8'h10 ;
			data[75213] <= 8'h10 ;
			data[75214] <= 8'h10 ;
			data[75215] <= 8'h10 ;
			data[75216] <= 8'h10 ;
			data[75217] <= 8'h10 ;
			data[75218] <= 8'h10 ;
			data[75219] <= 8'h10 ;
			data[75220] <= 8'h10 ;
			data[75221] <= 8'h10 ;
			data[75222] <= 8'h10 ;
			data[75223] <= 8'h10 ;
			data[75224] <= 8'h10 ;
			data[75225] <= 8'h10 ;
			data[75226] <= 8'h10 ;
			data[75227] <= 8'h10 ;
			data[75228] <= 8'h10 ;
			data[75229] <= 8'h10 ;
			data[75230] <= 8'h10 ;
			data[75231] <= 8'h10 ;
			data[75232] <= 8'h10 ;
			data[75233] <= 8'h10 ;
			data[75234] <= 8'h10 ;
			data[75235] <= 8'h10 ;
			data[75236] <= 8'h10 ;
			data[75237] <= 8'h10 ;
			data[75238] <= 8'h10 ;
			data[75239] <= 8'h10 ;
			data[75240] <= 8'h10 ;
			data[75241] <= 8'h10 ;
			data[75242] <= 8'h10 ;
			data[75243] <= 8'h10 ;
			data[75244] <= 8'h10 ;
			data[75245] <= 8'h10 ;
			data[75246] <= 8'h10 ;
			data[75247] <= 8'h10 ;
			data[75248] <= 8'h10 ;
			data[75249] <= 8'h10 ;
			data[75250] <= 8'h10 ;
			data[75251] <= 8'h10 ;
			data[75252] <= 8'h10 ;
			data[75253] <= 8'h10 ;
			data[75254] <= 8'h10 ;
			data[75255] <= 8'h10 ;
			data[75256] <= 8'h10 ;
			data[75257] <= 8'h10 ;
			data[75258] <= 8'h10 ;
			data[75259] <= 8'h10 ;
			data[75260] <= 8'h10 ;
			data[75261] <= 8'h10 ;
			data[75262] <= 8'h10 ;
			data[75263] <= 8'h10 ;
			data[75264] <= 8'h10 ;
			data[75265] <= 8'h10 ;
			data[75266] <= 8'h10 ;
			data[75267] <= 8'h10 ;
			data[75268] <= 8'h10 ;
			data[75269] <= 8'h10 ;
			data[75270] <= 8'h10 ;
			data[75271] <= 8'h10 ;
			data[75272] <= 8'h10 ;
			data[75273] <= 8'h10 ;
			data[75274] <= 8'h10 ;
			data[75275] <= 8'h10 ;
			data[75276] <= 8'h10 ;
			data[75277] <= 8'h10 ;
			data[75278] <= 8'h10 ;
			data[75279] <= 8'h10 ;
			data[75280] <= 8'h10 ;
			data[75281] <= 8'h10 ;
			data[75282] <= 8'h10 ;
			data[75283] <= 8'h10 ;
			data[75284] <= 8'h10 ;
			data[75285] <= 8'h10 ;
			data[75286] <= 8'h10 ;
			data[75287] <= 8'h10 ;
			data[75288] <= 8'h10 ;
			data[75289] <= 8'h10 ;
			data[75290] <= 8'h10 ;
			data[75291] <= 8'h10 ;
			data[75292] <= 8'h10 ;
			data[75293] <= 8'h10 ;
			data[75294] <= 8'h10 ;
			data[75295] <= 8'h10 ;
			data[75296] <= 8'h10 ;
			data[75297] <= 8'h10 ;
			data[75298] <= 8'h10 ;
			data[75299] <= 8'h10 ;
			data[75300] <= 8'h10 ;
			data[75301] <= 8'h10 ;
			data[75302] <= 8'h10 ;
			data[75303] <= 8'h10 ;
			data[75304] <= 8'h10 ;
			data[75305] <= 8'h10 ;
			data[75306] <= 8'h10 ;
			data[75307] <= 8'h10 ;
			data[75308] <= 8'h10 ;
			data[75309] <= 8'h10 ;
			data[75310] <= 8'h10 ;
			data[75311] <= 8'h10 ;
			data[75312] <= 8'h10 ;
			data[75313] <= 8'h10 ;
			data[75314] <= 8'h10 ;
			data[75315] <= 8'h10 ;
			data[75316] <= 8'h10 ;
			data[75317] <= 8'h10 ;
			data[75318] <= 8'h10 ;
			data[75319] <= 8'h10 ;
			data[75320] <= 8'h10 ;
			data[75321] <= 8'h10 ;
			data[75322] <= 8'h10 ;
			data[75323] <= 8'h10 ;
			data[75324] <= 8'h10 ;
			data[75325] <= 8'h10 ;
			data[75326] <= 8'h10 ;
			data[75327] <= 8'h10 ;
			data[75328] <= 8'h10 ;
			data[75329] <= 8'h10 ;
			data[75330] <= 8'h10 ;
			data[75331] <= 8'h10 ;
			data[75332] <= 8'h10 ;
			data[75333] <= 8'h10 ;
			data[75334] <= 8'h10 ;
			data[75335] <= 8'h10 ;
			data[75336] <= 8'h10 ;
			data[75337] <= 8'h10 ;
			data[75338] <= 8'h10 ;
			data[75339] <= 8'h10 ;
			data[75340] <= 8'h10 ;
			data[75341] <= 8'h10 ;
			data[75342] <= 8'h10 ;
			data[75343] <= 8'h10 ;
			data[75344] <= 8'h10 ;
			data[75345] <= 8'h10 ;
			data[75346] <= 8'h10 ;
			data[75347] <= 8'h10 ;
			data[75348] <= 8'h10 ;
			data[75349] <= 8'h10 ;
			data[75350] <= 8'h10 ;
			data[75351] <= 8'h10 ;
			data[75352] <= 8'h10 ;
			data[75353] <= 8'h10 ;
			data[75354] <= 8'h10 ;
			data[75355] <= 8'h10 ;
			data[75356] <= 8'h10 ;
			data[75357] <= 8'h10 ;
			data[75358] <= 8'h10 ;
			data[75359] <= 8'h10 ;
			data[75360] <= 8'h10 ;
			data[75361] <= 8'h10 ;
			data[75362] <= 8'h10 ;
			data[75363] <= 8'h10 ;
			data[75364] <= 8'h10 ;
			data[75365] <= 8'h10 ;
			data[75366] <= 8'h10 ;
			data[75367] <= 8'h10 ;
			data[75368] <= 8'h10 ;
			data[75369] <= 8'h10 ;
			data[75370] <= 8'h10 ;
			data[75371] <= 8'h10 ;
			data[75372] <= 8'h10 ;
			data[75373] <= 8'h10 ;
			data[75374] <= 8'h10 ;
			data[75375] <= 8'h10 ;
			data[75376] <= 8'h10 ;
			data[75377] <= 8'h10 ;
			data[75378] <= 8'h10 ;
			data[75379] <= 8'h10 ;
			data[75380] <= 8'h10 ;
			data[75381] <= 8'h10 ;
			data[75382] <= 8'h10 ;
			data[75383] <= 8'h10 ;
			data[75384] <= 8'h10 ;
			data[75385] <= 8'h10 ;
			data[75386] <= 8'h10 ;
			data[75387] <= 8'h10 ;
			data[75388] <= 8'h10 ;
			data[75389] <= 8'h10 ;
			data[75390] <= 8'h10 ;
			data[75391] <= 8'h10 ;
			data[75392] <= 8'h10 ;
			data[75393] <= 8'h10 ;
			data[75394] <= 8'h10 ;
			data[75395] <= 8'h10 ;
			data[75396] <= 8'h10 ;
			data[75397] <= 8'h10 ;
			data[75398] <= 8'h10 ;
			data[75399] <= 8'h10 ;
			data[75400] <= 8'h10 ;
			data[75401] <= 8'h10 ;
			data[75402] <= 8'h10 ;
			data[75403] <= 8'h10 ;
			data[75404] <= 8'h10 ;
			data[75405] <= 8'h10 ;
			data[75406] <= 8'h10 ;
			data[75407] <= 8'h10 ;
			data[75408] <= 8'h10 ;
			data[75409] <= 8'h10 ;
			data[75410] <= 8'h10 ;
			data[75411] <= 8'h10 ;
			data[75412] <= 8'h10 ;
			data[75413] <= 8'h10 ;
			data[75414] <= 8'h10 ;
			data[75415] <= 8'h10 ;
			data[75416] <= 8'h10 ;
			data[75417] <= 8'h10 ;
			data[75418] <= 8'h10 ;
			data[75419] <= 8'h10 ;
			data[75420] <= 8'h10 ;
			data[75421] <= 8'h10 ;
			data[75422] <= 8'h10 ;
			data[75423] <= 8'h10 ;
			data[75424] <= 8'h10 ;
			data[75425] <= 8'h10 ;
			data[75426] <= 8'h10 ;
			data[75427] <= 8'h10 ;
			data[75428] <= 8'h10 ;
			data[75429] <= 8'h10 ;
			data[75430] <= 8'h10 ;
			data[75431] <= 8'h10 ;
			data[75432] <= 8'h10 ;
			data[75433] <= 8'h10 ;
			data[75434] <= 8'h10 ;
			data[75435] <= 8'h10 ;
			data[75436] <= 8'h10 ;
			data[75437] <= 8'h10 ;
			data[75438] <= 8'h10 ;
			data[75439] <= 8'h10 ;
			data[75440] <= 8'h10 ;
			data[75441] <= 8'h10 ;
			data[75442] <= 8'h10 ;
			data[75443] <= 8'h10 ;
			data[75444] <= 8'h10 ;
			data[75445] <= 8'h10 ;
			data[75446] <= 8'h10 ;
			data[75447] <= 8'h10 ;
			data[75448] <= 8'h10 ;
			data[75449] <= 8'h10 ;
			data[75450] <= 8'h10 ;
			data[75451] <= 8'h10 ;
			data[75452] <= 8'h10 ;
			data[75453] <= 8'h10 ;
			data[75454] <= 8'h10 ;
			data[75455] <= 8'h10 ;
			data[75456] <= 8'h10 ;
			data[75457] <= 8'h10 ;
			data[75458] <= 8'h10 ;
			data[75459] <= 8'h10 ;
			data[75460] <= 8'h10 ;
			data[75461] <= 8'h10 ;
			data[75462] <= 8'h10 ;
			data[75463] <= 8'h10 ;
			data[75464] <= 8'h10 ;
			data[75465] <= 8'h10 ;
			data[75466] <= 8'h10 ;
			data[75467] <= 8'h10 ;
			data[75468] <= 8'h10 ;
			data[75469] <= 8'h10 ;
			data[75470] <= 8'h10 ;
			data[75471] <= 8'h10 ;
			data[75472] <= 8'h10 ;
			data[75473] <= 8'h10 ;
			data[75474] <= 8'h10 ;
			data[75475] <= 8'h10 ;
			data[75476] <= 8'h10 ;
			data[75477] <= 8'h10 ;
			data[75478] <= 8'h10 ;
			data[75479] <= 8'h10 ;
			data[75480] <= 8'h10 ;
			data[75481] <= 8'h10 ;
			data[75482] <= 8'h10 ;
			data[75483] <= 8'h10 ;
			data[75484] <= 8'h10 ;
			data[75485] <= 8'h10 ;
			data[75486] <= 8'h10 ;
			data[75487] <= 8'h10 ;
			data[75488] <= 8'h10 ;
			data[75489] <= 8'h10 ;
			data[75490] <= 8'h10 ;
			data[75491] <= 8'h10 ;
			data[75492] <= 8'h10 ;
			data[75493] <= 8'h10 ;
			data[75494] <= 8'h10 ;
			data[75495] <= 8'h10 ;
			data[75496] <= 8'h10 ;
			data[75497] <= 8'h10 ;
			data[75498] <= 8'h10 ;
			data[75499] <= 8'h10 ;
			data[75500] <= 8'h10 ;
			data[75501] <= 8'h10 ;
			data[75502] <= 8'h10 ;
			data[75503] <= 8'h10 ;
			data[75504] <= 8'h10 ;
			data[75505] <= 8'h10 ;
			data[75506] <= 8'h10 ;
			data[75507] <= 8'h10 ;
			data[75508] <= 8'h10 ;
			data[75509] <= 8'h10 ;
			data[75510] <= 8'h10 ;
			data[75511] <= 8'h10 ;
			data[75512] <= 8'h10 ;
			data[75513] <= 8'h10 ;
			data[75514] <= 8'h10 ;
			data[75515] <= 8'h10 ;
			data[75516] <= 8'h10 ;
			data[75517] <= 8'h10 ;
			data[75518] <= 8'h10 ;
			data[75519] <= 8'h10 ;
			data[75520] <= 8'h10 ;
			data[75521] <= 8'h10 ;
			data[75522] <= 8'h10 ;
			data[75523] <= 8'h10 ;
			data[75524] <= 8'h10 ;
			data[75525] <= 8'h10 ;
			data[75526] <= 8'h10 ;
			data[75527] <= 8'h10 ;
			data[75528] <= 8'h10 ;
			data[75529] <= 8'h10 ;
			data[75530] <= 8'h10 ;
			data[75531] <= 8'h10 ;
			data[75532] <= 8'h10 ;
			data[75533] <= 8'h10 ;
			data[75534] <= 8'h10 ;
			data[75535] <= 8'h10 ;
			data[75536] <= 8'h10 ;
			data[75537] <= 8'h10 ;
			data[75538] <= 8'h10 ;
			data[75539] <= 8'h10 ;
			data[75540] <= 8'h10 ;
			data[75541] <= 8'h10 ;
			data[75542] <= 8'h10 ;
			data[75543] <= 8'h10 ;
			data[75544] <= 8'h10 ;
			data[75545] <= 8'h10 ;
			data[75546] <= 8'h10 ;
			data[75547] <= 8'h10 ;
			data[75548] <= 8'h10 ;
			data[75549] <= 8'h10 ;
			data[75550] <= 8'h10 ;
			data[75551] <= 8'h10 ;
			data[75552] <= 8'h10 ;
			data[75553] <= 8'h10 ;
			data[75554] <= 8'h10 ;
			data[75555] <= 8'h10 ;
			data[75556] <= 8'h10 ;
			data[75557] <= 8'h10 ;
			data[75558] <= 8'h10 ;
			data[75559] <= 8'h10 ;
			data[75560] <= 8'h10 ;
			data[75561] <= 8'h10 ;
			data[75562] <= 8'h10 ;
			data[75563] <= 8'h10 ;
			data[75564] <= 8'h10 ;
			data[75565] <= 8'h10 ;
			data[75566] <= 8'h10 ;
			data[75567] <= 8'h10 ;
			data[75568] <= 8'h10 ;
			data[75569] <= 8'h10 ;
			data[75570] <= 8'h10 ;
			data[75571] <= 8'h10 ;
			data[75572] <= 8'h10 ;
			data[75573] <= 8'h10 ;
			data[75574] <= 8'h10 ;
			data[75575] <= 8'h10 ;
			data[75576] <= 8'h10 ;
			data[75577] <= 8'h10 ;
			data[75578] <= 8'h10 ;
			data[75579] <= 8'h10 ;
			data[75580] <= 8'h10 ;
			data[75581] <= 8'h10 ;
			data[75582] <= 8'h10 ;
			data[75583] <= 8'h10 ;
			data[75584] <= 8'h10 ;
			data[75585] <= 8'h10 ;
			data[75586] <= 8'h10 ;
			data[75587] <= 8'h10 ;
			data[75588] <= 8'h10 ;
			data[75589] <= 8'h10 ;
			data[75590] <= 8'h10 ;
			data[75591] <= 8'h10 ;
			data[75592] <= 8'h10 ;
			data[75593] <= 8'h10 ;
			data[75594] <= 8'h10 ;
			data[75595] <= 8'h10 ;
			data[75596] <= 8'h10 ;
			data[75597] <= 8'h10 ;
			data[75598] <= 8'h10 ;
			data[75599] <= 8'h10 ;
			data[75600] <= 8'h10 ;
			data[75601] <= 8'h10 ;
			data[75602] <= 8'h10 ;
			data[75603] <= 8'h10 ;
			data[75604] <= 8'h10 ;
			data[75605] <= 8'h10 ;
			data[75606] <= 8'h10 ;
			data[75607] <= 8'h10 ;
			data[75608] <= 8'h10 ;
			data[75609] <= 8'h10 ;
			data[75610] <= 8'h10 ;
			data[75611] <= 8'h10 ;
			data[75612] <= 8'h10 ;
			data[75613] <= 8'h10 ;
			data[75614] <= 8'h10 ;
			data[75615] <= 8'h10 ;
			data[75616] <= 8'h10 ;
			data[75617] <= 8'h10 ;
			data[75618] <= 8'h10 ;
			data[75619] <= 8'h10 ;
			data[75620] <= 8'h10 ;
			data[75621] <= 8'h10 ;
			data[75622] <= 8'h10 ;
			data[75623] <= 8'h10 ;
			data[75624] <= 8'h10 ;
			data[75625] <= 8'h10 ;
			data[75626] <= 8'h10 ;
			data[75627] <= 8'h10 ;
			data[75628] <= 8'h10 ;
			data[75629] <= 8'h10 ;
			data[75630] <= 8'h10 ;
			data[75631] <= 8'h10 ;
			data[75632] <= 8'h10 ;
			data[75633] <= 8'h10 ;
			data[75634] <= 8'h10 ;
			data[75635] <= 8'h10 ;
			data[75636] <= 8'h10 ;
			data[75637] <= 8'h10 ;
			data[75638] <= 8'h10 ;
			data[75639] <= 8'h10 ;
			data[75640] <= 8'h10 ;
			data[75641] <= 8'h10 ;
			data[75642] <= 8'h10 ;
			data[75643] <= 8'h10 ;
			data[75644] <= 8'h10 ;
			data[75645] <= 8'h10 ;
			data[75646] <= 8'h10 ;
			data[75647] <= 8'h10 ;
			data[75648] <= 8'h10 ;
			data[75649] <= 8'h10 ;
			data[75650] <= 8'h10 ;
			data[75651] <= 8'h10 ;
			data[75652] <= 8'h10 ;
			data[75653] <= 8'h10 ;
			data[75654] <= 8'h10 ;
			data[75655] <= 8'h10 ;
			data[75656] <= 8'h10 ;
			data[75657] <= 8'h10 ;
			data[75658] <= 8'h10 ;
			data[75659] <= 8'h10 ;
			data[75660] <= 8'h10 ;
			data[75661] <= 8'h10 ;
			data[75662] <= 8'h10 ;
			data[75663] <= 8'h10 ;
			data[75664] <= 8'h10 ;
			data[75665] <= 8'h10 ;
			data[75666] <= 8'h10 ;
			data[75667] <= 8'h10 ;
			data[75668] <= 8'h10 ;
			data[75669] <= 8'h10 ;
			data[75670] <= 8'h10 ;
			data[75671] <= 8'h10 ;
			data[75672] <= 8'h10 ;
			data[75673] <= 8'h10 ;
			data[75674] <= 8'h10 ;
			data[75675] <= 8'h10 ;
			data[75676] <= 8'h10 ;
			data[75677] <= 8'h10 ;
			data[75678] <= 8'h10 ;
			data[75679] <= 8'h10 ;
			data[75680] <= 8'h10 ;
			data[75681] <= 8'h10 ;
			data[75682] <= 8'h10 ;
			data[75683] <= 8'h10 ;
			data[75684] <= 8'h10 ;
			data[75685] <= 8'h10 ;
			data[75686] <= 8'h10 ;
			data[75687] <= 8'h10 ;
			data[75688] <= 8'h10 ;
			data[75689] <= 8'h10 ;
			data[75690] <= 8'h10 ;
			data[75691] <= 8'h10 ;
			data[75692] <= 8'h10 ;
			data[75693] <= 8'h10 ;
			data[75694] <= 8'h10 ;
			data[75695] <= 8'h10 ;
			data[75696] <= 8'h10 ;
			data[75697] <= 8'h10 ;
			data[75698] <= 8'h10 ;
			data[75699] <= 8'h10 ;
			data[75700] <= 8'h10 ;
			data[75701] <= 8'h10 ;
			data[75702] <= 8'h10 ;
			data[75703] <= 8'h10 ;
			data[75704] <= 8'h10 ;
			data[75705] <= 8'h10 ;
			data[75706] <= 8'h10 ;
			data[75707] <= 8'h10 ;
			data[75708] <= 8'h10 ;
			data[75709] <= 8'h10 ;
			data[75710] <= 8'h10 ;
			data[75711] <= 8'h10 ;
			data[75712] <= 8'h10 ;
			data[75713] <= 8'h10 ;
			data[75714] <= 8'h10 ;
			data[75715] <= 8'h10 ;
			data[75716] <= 8'h10 ;
			data[75717] <= 8'h10 ;
			data[75718] <= 8'h10 ;
			data[75719] <= 8'h10 ;
			data[75720] <= 8'h10 ;
			data[75721] <= 8'h10 ;
			data[75722] <= 8'h10 ;
			data[75723] <= 8'h10 ;
			data[75724] <= 8'h10 ;
			data[75725] <= 8'h10 ;
			data[75726] <= 8'h10 ;
			data[75727] <= 8'h10 ;
			data[75728] <= 8'h10 ;
			data[75729] <= 8'h10 ;
			data[75730] <= 8'h10 ;
			data[75731] <= 8'h10 ;
			data[75732] <= 8'h10 ;
			data[75733] <= 8'h10 ;
			data[75734] <= 8'h10 ;
			data[75735] <= 8'h10 ;
			data[75736] <= 8'h10 ;
			data[75737] <= 8'h10 ;
			data[75738] <= 8'h10 ;
			data[75739] <= 8'h10 ;
			data[75740] <= 8'h10 ;
			data[75741] <= 8'h10 ;
			data[75742] <= 8'h10 ;
			data[75743] <= 8'h10 ;
			data[75744] <= 8'h10 ;
			data[75745] <= 8'h10 ;
			data[75746] <= 8'h10 ;
			data[75747] <= 8'h10 ;
			data[75748] <= 8'h10 ;
			data[75749] <= 8'h10 ;
			data[75750] <= 8'h10 ;
			data[75751] <= 8'h10 ;
			data[75752] <= 8'h10 ;
			data[75753] <= 8'h10 ;
			data[75754] <= 8'h10 ;
			data[75755] <= 8'h10 ;
			data[75756] <= 8'h10 ;
			data[75757] <= 8'h10 ;
			data[75758] <= 8'h10 ;
			data[75759] <= 8'h10 ;
			data[75760] <= 8'h10 ;
			data[75761] <= 8'h10 ;
			data[75762] <= 8'h10 ;
			data[75763] <= 8'h10 ;
			data[75764] <= 8'h10 ;
			data[75765] <= 8'h10 ;
			data[75766] <= 8'h10 ;
			data[75767] <= 8'h10 ;
			data[75768] <= 8'h10 ;
			data[75769] <= 8'h10 ;
			data[75770] <= 8'h10 ;
			data[75771] <= 8'h10 ;
			data[75772] <= 8'h10 ;
			data[75773] <= 8'h10 ;
			data[75774] <= 8'h10 ;
			data[75775] <= 8'h10 ;
			data[75776] <= 8'h10 ;
			data[75777] <= 8'h10 ;
			data[75778] <= 8'h10 ;
			data[75779] <= 8'h10 ;
			data[75780] <= 8'h10 ;
			data[75781] <= 8'h10 ;
			data[75782] <= 8'h10 ;
			data[75783] <= 8'h10 ;
			data[75784] <= 8'h10 ;
			data[75785] <= 8'h10 ;
			data[75786] <= 8'h10 ;
			data[75787] <= 8'h10 ;
			data[75788] <= 8'h10 ;
			data[75789] <= 8'h10 ;
			data[75790] <= 8'h10 ;
			data[75791] <= 8'h10 ;
			data[75792] <= 8'h10 ;
			data[75793] <= 8'h10 ;
			data[75794] <= 8'h10 ;
			data[75795] <= 8'h10 ;
			data[75796] <= 8'h10 ;
			data[75797] <= 8'h10 ;
			data[75798] <= 8'h10 ;
			data[75799] <= 8'h10 ;
			data[75800] <= 8'h10 ;
			data[75801] <= 8'h10 ;
			data[75802] <= 8'h10 ;
			data[75803] <= 8'h10 ;
			data[75804] <= 8'h10 ;
			data[75805] <= 8'h10 ;
			data[75806] <= 8'h10 ;
			data[75807] <= 8'h10 ;
			data[75808] <= 8'h10 ;
			data[75809] <= 8'h10 ;
			data[75810] <= 8'h10 ;
			data[75811] <= 8'h10 ;
			data[75812] <= 8'h10 ;
			data[75813] <= 8'h10 ;
			data[75814] <= 8'h10 ;
			data[75815] <= 8'h10 ;
			data[75816] <= 8'h10 ;
			data[75817] <= 8'h10 ;
			data[75818] <= 8'h10 ;
			data[75819] <= 8'h10 ;
			data[75820] <= 8'h10 ;
			data[75821] <= 8'h10 ;
			data[75822] <= 8'h10 ;
			data[75823] <= 8'h10 ;
			data[75824] <= 8'h10 ;
			data[75825] <= 8'h10 ;
			data[75826] <= 8'h10 ;
			data[75827] <= 8'h10 ;
			data[75828] <= 8'h10 ;
			data[75829] <= 8'h10 ;
			data[75830] <= 8'h10 ;
			data[75831] <= 8'h10 ;
			data[75832] <= 8'h10 ;
			data[75833] <= 8'h10 ;
			data[75834] <= 8'h10 ;
			data[75835] <= 8'h10 ;
			data[75836] <= 8'h10 ;
			data[75837] <= 8'h10 ;
			data[75838] <= 8'h10 ;
			data[75839] <= 8'h10 ;
			data[75840] <= 8'h10 ;
			data[75841] <= 8'h10 ;
			data[75842] <= 8'h10 ;
			data[75843] <= 8'h10 ;
			data[75844] <= 8'h10 ;
			data[75845] <= 8'h10 ;
			data[75846] <= 8'h10 ;
			data[75847] <= 8'h10 ;
			data[75848] <= 8'h10 ;
			data[75849] <= 8'h10 ;
			data[75850] <= 8'h10 ;
			data[75851] <= 8'h10 ;
			data[75852] <= 8'h10 ;
			data[75853] <= 8'h10 ;
			data[75854] <= 8'h10 ;
			data[75855] <= 8'h10 ;
			data[75856] <= 8'h10 ;
			data[75857] <= 8'h10 ;
			data[75858] <= 8'h10 ;
			data[75859] <= 8'h10 ;
			data[75860] <= 8'h10 ;
			data[75861] <= 8'h10 ;
			data[75862] <= 8'h10 ;
			data[75863] <= 8'h10 ;
			data[75864] <= 8'h10 ;
			data[75865] <= 8'h10 ;
			data[75866] <= 8'h10 ;
			data[75867] <= 8'h10 ;
			data[75868] <= 8'h10 ;
			data[75869] <= 8'h10 ;
			data[75870] <= 8'h10 ;
			data[75871] <= 8'h10 ;
			data[75872] <= 8'h10 ;
			data[75873] <= 8'h10 ;
			data[75874] <= 8'h10 ;
			data[75875] <= 8'h10 ;
			data[75876] <= 8'h10 ;
			data[75877] <= 8'h10 ;
			data[75878] <= 8'h10 ;
			data[75879] <= 8'h10 ;
			data[75880] <= 8'h10 ;
			data[75881] <= 8'h10 ;
			data[75882] <= 8'h10 ;
			data[75883] <= 8'h10 ;
			data[75884] <= 8'h10 ;
			data[75885] <= 8'h10 ;
			data[75886] <= 8'h10 ;
			data[75887] <= 8'h10 ;
			data[75888] <= 8'h10 ;
			data[75889] <= 8'h10 ;
			data[75890] <= 8'h10 ;
			data[75891] <= 8'h10 ;
			data[75892] <= 8'h10 ;
			data[75893] <= 8'h10 ;
			data[75894] <= 8'h10 ;
			data[75895] <= 8'h10 ;
			data[75896] <= 8'h10 ;
			data[75897] <= 8'h10 ;
			data[75898] <= 8'h10 ;
			data[75899] <= 8'h10 ;
			data[75900] <= 8'h10 ;
			data[75901] <= 8'h10 ;
			data[75902] <= 8'h10 ;
			data[75903] <= 8'h10 ;
			data[75904] <= 8'h10 ;
			data[75905] <= 8'h10 ;
			data[75906] <= 8'h10 ;
			data[75907] <= 8'h10 ;
			data[75908] <= 8'h10 ;
			data[75909] <= 8'h10 ;
			data[75910] <= 8'h10 ;
			data[75911] <= 8'h10 ;
			data[75912] <= 8'h10 ;
			data[75913] <= 8'h10 ;
			data[75914] <= 8'h10 ;
			data[75915] <= 8'h10 ;
			data[75916] <= 8'h10 ;
			data[75917] <= 8'h10 ;
			data[75918] <= 8'h10 ;
			data[75919] <= 8'h10 ;
			data[75920] <= 8'h10 ;
			data[75921] <= 8'h10 ;
			data[75922] <= 8'h10 ;
			data[75923] <= 8'h10 ;
			data[75924] <= 8'h10 ;
			data[75925] <= 8'h10 ;
			data[75926] <= 8'h10 ;
			data[75927] <= 8'h10 ;
			data[75928] <= 8'h10 ;
			data[75929] <= 8'h10 ;
			data[75930] <= 8'h10 ;
			data[75931] <= 8'h10 ;
			data[75932] <= 8'h10 ;
			data[75933] <= 8'h10 ;
			data[75934] <= 8'h10 ;
			data[75935] <= 8'h10 ;
			data[75936] <= 8'h10 ;
			data[75937] <= 8'h10 ;
			data[75938] <= 8'h10 ;
			data[75939] <= 8'h10 ;
			data[75940] <= 8'h10 ;
			data[75941] <= 8'h10 ;
			data[75942] <= 8'h10 ;
			data[75943] <= 8'h10 ;
			data[75944] <= 8'h10 ;
			data[75945] <= 8'h10 ;
			data[75946] <= 8'h10 ;
			data[75947] <= 8'h10 ;
			data[75948] <= 8'h10 ;
			data[75949] <= 8'h10 ;
			data[75950] <= 8'h10 ;
			data[75951] <= 8'h10 ;
			data[75952] <= 8'h10 ;
			data[75953] <= 8'h10 ;
			data[75954] <= 8'h10 ;
			data[75955] <= 8'h10 ;
			data[75956] <= 8'h10 ;
			data[75957] <= 8'h10 ;
			data[75958] <= 8'h10 ;
			data[75959] <= 8'h10 ;
			data[75960] <= 8'h10 ;
			data[75961] <= 8'h10 ;
			data[75962] <= 8'h10 ;
			data[75963] <= 8'h10 ;
			data[75964] <= 8'h10 ;
			data[75965] <= 8'h10 ;
			data[75966] <= 8'h10 ;
			data[75967] <= 8'h10 ;
			data[75968] <= 8'h10 ;
			data[75969] <= 8'h10 ;
			data[75970] <= 8'h10 ;
			data[75971] <= 8'h10 ;
			data[75972] <= 8'h10 ;
			data[75973] <= 8'h10 ;
			data[75974] <= 8'h10 ;
			data[75975] <= 8'h10 ;
			data[75976] <= 8'h10 ;
			data[75977] <= 8'h10 ;
			data[75978] <= 8'h10 ;
			data[75979] <= 8'h10 ;
			data[75980] <= 8'h10 ;
			data[75981] <= 8'h10 ;
			data[75982] <= 8'h10 ;
			data[75983] <= 8'h10 ;
			data[75984] <= 8'h10 ;
			data[75985] <= 8'h10 ;
			data[75986] <= 8'h10 ;
			data[75987] <= 8'h10 ;
			data[75988] <= 8'h10 ;
			data[75989] <= 8'h10 ;
			data[75990] <= 8'h10 ;
			data[75991] <= 8'h10 ;
			data[75992] <= 8'h10 ;
			data[75993] <= 8'h10 ;
			data[75994] <= 8'h10 ;
			data[75995] <= 8'h10 ;
			data[75996] <= 8'h10 ;
			data[75997] <= 8'h10 ;
			data[75998] <= 8'h10 ;
			data[75999] <= 8'h10 ;
			data[76000] <= 8'h10 ;
			data[76001] <= 8'h10 ;
			data[76002] <= 8'h10 ;
			data[76003] <= 8'h10 ;
			data[76004] <= 8'h10 ;
			data[76005] <= 8'h10 ;
			data[76006] <= 8'h10 ;
			data[76007] <= 8'h10 ;
			data[76008] <= 8'h10 ;
			data[76009] <= 8'h10 ;
			data[76010] <= 8'h10 ;
			data[76011] <= 8'h10 ;
			data[76012] <= 8'h10 ;
			data[76013] <= 8'h10 ;
			data[76014] <= 8'h10 ;
			data[76015] <= 8'h10 ;
			data[76016] <= 8'h10 ;
			data[76017] <= 8'h10 ;
			data[76018] <= 8'h10 ;
			data[76019] <= 8'h10 ;
			data[76020] <= 8'h10 ;
			data[76021] <= 8'h10 ;
			data[76022] <= 8'h10 ;
			data[76023] <= 8'h10 ;
			data[76024] <= 8'h10 ;
			data[76025] <= 8'h10 ;
			data[76026] <= 8'h10 ;
			data[76027] <= 8'h10 ;
			data[76028] <= 8'h10 ;
			data[76029] <= 8'h10 ;
			data[76030] <= 8'h10 ;
			data[76031] <= 8'h10 ;
			data[76032] <= 8'h10 ;
			data[76033] <= 8'h10 ;
			data[76034] <= 8'h10 ;
			data[76035] <= 8'h10 ;
			data[76036] <= 8'h10 ;
			data[76037] <= 8'h10 ;
			data[76038] <= 8'h10 ;
			data[76039] <= 8'h10 ;
			data[76040] <= 8'h10 ;
			data[76041] <= 8'h10 ;
			data[76042] <= 8'h10 ;
			data[76043] <= 8'h10 ;
			data[76044] <= 8'h10 ;
			data[76045] <= 8'h10 ;
			data[76046] <= 8'h10 ;
			data[76047] <= 8'h10 ;
			data[76048] <= 8'h10 ;
			data[76049] <= 8'h10 ;
			data[76050] <= 8'h10 ;
			data[76051] <= 8'h10 ;
			data[76052] <= 8'h10 ;
			data[76053] <= 8'h10 ;
			data[76054] <= 8'h10 ;
			data[76055] <= 8'h10 ;
			data[76056] <= 8'h10 ;
			data[76057] <= 8'h10 ;
			data[76058] <= 8'h10 ;
			data[76059] <= 8'h10 ;
			data[76060] <= 8'h10 ;
			data[76061] <= 8'h10 ;
			data[76062] <= 8'h10 ;
			data[76063] <= 8'h10 ;
			data[76064] <= 8'h10 ;
			data[76065] <= 8'h10 ;
			data[76066] <= 8'h10 ;
			data[76067] <= 8'h10 ;
			data[76068] <= 8'h10 ;
			data[76069] <= 8'h10 ;
			data[76070] <= 8'h10 ;
			data[76071] <= 8'h10 ;
			data[76072] <= 8'h10 ;
			data[76073] <= 8'h10 ;
			data[76074] <= 8'h10 ;
			data[76075] <= 8'h10 ;
			data[76076] <= 8'h10 ;
			data[76077] <= 8'h10 ;
			data[76078] <= 8'h10 ;
			data[76079] <= 8'h10 ;
			data[76080] <= 8'h10 ;
			data[76081] <= 8'h10 ;
			data[76082] <= 8'h10 ;
			data[76083] <= 8'h10 ;
			data[76084] <= 8'h10 ;
			data[76085] <= 8'h10 ;
			data[76086] <= 8'h10 ;
			data[76087] <= 8'h10 ;
			data[76088] <= 8'h10 ;
			data[76089] <= 8'h10 ;
			data[76090] <= 8'h10 ;
			data[76091] <= 8'h10 ;
			data[76092] <= 8'h10 ;
			data[76093] <= 8'h10 ;
			data[76094] <= 8'h10 ;
			data[76095] <= 8'h10 ;
			data[76096] <= 8'h10 ;
			data[76097] <= 8'h10 ;
			data[76098] <= 8'h10 ;
			data[76099] <= 8'h10 ;
			data[76100] <= 8'h10 ;
			data[76101] <= 8'h10 ;
			data[76102] <= 8'h10 ;
			data[76103] <= 8'h10 ;
			data[76104] <= 8'h10 ;
			data[76105] <= 8'h10 ;
			data[76106] <= 8'h10 ;
			data[76107] <= 8'h10 ;
			data[76108] <= 8'h10 ;
			data[76109] <= 8'h10 ;
			data[76110] <= 8'h10 ;
			data[76111] <= 8'h10 ;
			data[76112] <= 8'h10 ;
			data[76113] <= 8'h10 ;
			data[76114] <= 8'h10 ;
			data[76115] <= 8'h10 ;
			data[76116] <= 8'h10 ;
			data[76117] <= 8'h10 ;
			data[76118] <= 8'h10 ;
			data[76119] <= 8'h10 ;
			data[76120] <= 8'h10 ;
			data[76121] <= 8'h10 ;
			data[76122] <= 8'h10 ;
			data[76123] <= 8'h10 ;
			data[76124] <= 8'h10 ;
			data[76125] <= 8'h10 ;
			data[76126] <= 8'h10 ;
			data[76127] <= 8'h10 ;
			data[76128] <= 8'h10 ;
			data[76129] <= 8'h10 ;
			data[76130] <= 8'h10 ;
			data[76131] <= 8'h10 ;
			data[76132] <= 8'h10 ;
			data[76133] <= 8'h10 ;
			data[76134] <= 8'h10 ;
			data[76135] <= 8'h10 ;
			data[76136] <= 8'h10 ;
			data[76137] <= 8'h10 ;
			data[76138] <= 8'h10 ;
			data[76139] <= 8'h10 ;
			data[76140] <= 8'h10 ;
			data[76141] <= 8'h10 ;
			data[76142] <= 8'h10 ;
			data[76143] <= 8'h10 ;
			data[76144] <= 8'h10 ;
			data[76145] <= 8'h10 ;
			data[76146] <= 8'h10 ;
			data[76147] <= 8'h10 ;
			data[76148] <= 8'h10 ;
			data[76149] <= 8'h10 ;
			data[76150] <= 8'h10 ;
			data[76151] <= 8'h10 ;
			data[76152] <= 8'h10 ;
			data[76153] <= 8'h10 ;
			data[76154] <= 8'h10 ;
			data[76155] <= 8'h10 ;
			data[76156] <= 8'h10 ;
			data[76157] <= 8'h10 ;
			data[76158] <= 8'h10 ;
			data[76159] <= 8'h10 ;
			data[76160] <= 8'h10 ;
			data[76161] <= 8'h10 ;
			data[76162] <= 8'h10 ;
			data[76163] <= 8'h10 ;
			data[76164] <= 8'h10 ;
			data[76165] <= 8'h10 ;
			data[76166] <= 8'h10 ;
			data[76167] <= 8'h10 ;
			data[76168] <= 8'h10 ;
			data[76169] <= 8'h10 ;
			data[76170] <= 8'h10 ;
			data[76171] <= 8'h10 ;
			data[76172] <= 8'h10 ;
			data[76173] <= 8'h10 ;
			data[76174] <= 8'h10 ;
			data[76175] <= 8'h10 ;
			data[76176] <= 8'h10 ;
			data[76177] <= 8'h10 ;
			data[76178] <= 8'h10 ;
			data[76179] <= 8'h10 ;
			data[76180] <= 8'h10 ;
			data[76181] <= 8'h10 ;
			data[76182] <= 8'h10 ;
			data[76183] <= 8'h10 ;
			data[76184] <= 8'h10 ;
			data[76185] <= 8'h10 ;
			data[76186] <= 8'h10 ;
			data[76187] <= 8'h10 ;
			data[76188] <= 8'h10 ;
			data[76189] <= 8'h10 ;
			data[76190] <= 8'h10 ;
			data[76191] <= 8'h10 ;
			data[76192] <= 8'h10 ;
			data[76193] <= 8'h10 ;
			data[76194] <= 8'h10 ;
			data[76195] <= 8'h10 ;
			data[76196] <= 8'h10 ;
			data[76197] <= 8'h10 ;
			data[76198] <= 8'h10 ;
			data[76199] <= 8'h10 ;
			data[76200] <= 8'h10 ;
			data[76201] <= 8'h10 ;
			data[76202] <= 8'h10 ;
			data[76203] <= 8'h10 ;
			data[76204] <= 8'h10 ;
			data[76205] <= 8'h10 ;
			data[76206] <= 8'h10 ;
			data[76207] <= 8'h10 ;
			data[76208] <= 8'h10 ;
			data[76209] <= 8'h10 ;
			data[76210] <= 8'h10 ;
			data[76211] <= 8'h10 ;
			data[76212] <= 8'h10 ;
			data[76213] <= 8'h10 ;
			data[76214] <= 8'h10 ;
			data[76215] <= 8'h10 ;
			data[76216] <= 8'h10 ;
			data[76217] <= 8'h10 ;
			data[76218] <= 8'h10 ;
			data[76219] <= 8'h10 ;
			data[76220] <= 8'h10 ;
			data[76221] <= 8'h10 ;
			data[76222] <= 8'h10 ;
			data[76223] <= 8'h10 ;
			data[76224] <= 8'h10 ;
			data[76225] <= 8'h10 ;
			data[76226] <= 8'h10 ;
			data[76227] <= 8'h10 ;
			data[76228] <= 8'h10 ;
			data[76229] <= 8'h10 ;
			data[76230] <= 8'h10 ;
			data[76231] <= 8'h10 ;
			data[76232] <= 8'h10 ;
			data[76233] <= 8'h10 ;
			data[76234] <= 8'h10 ;
			data[76235] <= 8'h10 ;
			data[76236] <= 8'h10 ;
			data[76237] <= 8'h10 ;
			data[76238] <= 8'h10 ;
			data[76239] <= 8'h10 ;
			data[76240] <= 8'h10 ;
			data[76241] <= 8'h10 ;
			data[76242] <= 8'h10 ;
			data[76243] <= 8'h10 ;
			data[76244] <= 8'h10 ;
			data[76245] <= 8'h10 ;
			data[76246] <= 8'h10 ;
			data[76247] <= 8'h10 ;
			data[76248] <= 8'h10 ;
			data[76249] <= 8'h10 ;
			data[76250] <= 8'h10 ;
			data[76251] <= 8'h10 ;
			data[76252] <= 8'h10 ;
			data[76253] <= 8'h10 ;
			data[76254] <= 8'h10 ;
			data[76255] <= 8'h10 ;
			data[76256] <= 8'h10 ;
			data[76257] <= 8'h10 ;
			data[76258] <= 8'h10 ;
			data[76259] <= 8'h10 ;
			data[76260] <= 8'h10 ;
			data[76261] <= 8'h10 ;
			data[76262] <= 8'h10 ;
			data[76263] <= 8'h10 ;
			data[76264] <= 8'h10 ;
			data[76265] <= 8'h10 ;
			data[76266] <= 8'h10 ;
			data[76267] <= 8'h10 ;
			data[76268] <= 8'h10 ;
			data[76269] <= 8'h10 ;
			data[76270] <= 8'h10 ;
			data[76271] <= 8'h10 ;
			data[76272] <= 8'h10 ;
			data[76273] <= 8'h10 ;
			data[76274] <= 8'h10 ;
			data[76275] <= 8'h10 ;
			data[76276] <= 8'h10 ;
			data[76277] <= 8'h10 ;
			data[76278] <= 8'h10 ;
			data[76279] <= 8'h10 ;
			data[76280] <= 8'h10 ;
			data[76281] <= 8'h10 ;
			data[76282] <= 8'h10 ;
			data[76283] <= 8'h10 ;
			data[76284] <= 8'h10 ;
			data[76285] <= 8'h10 ;
			data[76286] <= 8'h10 ;
			data[76287] <= 8'h10 ;
			data[76288] <= 8'h10 ;
			data[76289] <= 8'h10 ;
			data[76290] <= 8'h10 ;
			data[76291] <= 8'h10 ;
			data[76292] <= 8'h10 ;
			data[76293] <= 8'h10 ;
			data[76294] <= 8'h10 ;
			data[76295] <= 8'h10 ;
			data[76296] <= 8'h10 ;
			data[76297] <= 8'h10 ;
			data[76298] <= 8'h10 ;
			data[76299] <= 8'h10 ;
			data[76300] <= 8'h10 ;
			data[76301] <= 8'h10 ;
			data[76302] <= 8'h10 ;
			data[76303] <= 8'h10 ;
			data[76304] <= 8'h10 ;
			data[76305] <= 8'h10 ;
			data[76306] <= 8'h10 ;
			data[76307] <= 8'h10 ;
			data[76308] <= 8'h10 ;
			data[76309] <= 8'h10 ;
			data[76310] <= 8'h10 ;
			data[76311] <= 8'h10 ;
			data[76312] <= 8'h10 ;
			data[76313] <= 8'h10 ;
			data[76314] <= 8'h10 ;
			data[76315] <= 8'h10 ;
			data[76316] <= 8'h10 ;
			data[76317] <= 8'h10 ;
			data[76318] <= 8'h10 ;
			data[76319] <= 8'h10 ;
			data[76320] <= 8'h10 ;
			data[76321] <= 8'h10 ;
			data[76322] <= 8'h10 ;
			data[76323] <= 8'h10 ;
			data[76324] <= 8'h10 ;
			data[76325] <= 8'h10 ;
			data[76326] <= 8'h10 ;
			data[76327] <= 8'h10 ;
			data[76328] <= 8'h10 ;
			data[76329] <= 8'h10 ;
			data[76330] <= 8'h10 ;
			data[76331] <= 8'h10 ;
			data[76332] <= 8'h10 ;
			data[76333] <= 8'h10 ;
			data[76334] <= 8'h10 ;
			data[76335] <= 8'h10 ;
			data[76336] <= 8'h10 ;
			data[76337] <= 8'h10 ;
			data[76338] <= 8'h10 ;
			data[76339] <= 8'h10 ;
			data[76340] <= 8'h10 ;
			data[76341] <= 8'h10 ;
			data[76342] <= 8'h10 ;
			data[76343] <= 8'h10 ;
			data[76344] <= 8'h10 ;
			data[76345] <= 8'h10 ;
			data[76346] <= 8'h10 ;
			data[76347] <= 8'h10 ;
			data[76348] <= 8'h10 ;
			data[76349] <= 8'h10 ;
			data[76350] <= 8'h10 ;
			data[76351] <= 8'h10 ;
			data[76352] <= 8'h10 ;
			data[76353] <= 8'h10 ;
			data[76354] <= 8'h10 ;
			data[76355] <= 8'h10 ;
			data[76356] <= 8'h10 ;
			data[76357] <= 8'h10 ;
			data[76358] <= 8'h10 ;
			data[76359] <= 8'h10 ;
			data[76360] <= 8'h10 ;
			data[76361] <= 8'h10 ;
			data[76362] <= 8'h10 ;
			data[76363] <= 8'h10 ;
			data[76364] <= 8'h10 ;
			data[76365] <= 8'h10 ;
			data[76366] <= 8'h10 ;
			data[76367] <= 8'h10 ;
			data[76368] <= 8'h10 ;
			data[76369] <= 8'h10 ;
			data[76370] <= 8'h10 ;
			data[76371] <= 8'h10 ;
			data[76372] <= 8'h10 ;
			data[76373] <= 8'h10 ;
			data[76374] <= 8'h10 ;
			data[76375] <= 8'h10 ;
			data[76376] <= 8'h10 ;
			data[76377] <= 8'h10 ;
			data[76378] <= 8'h10 ;
			data[76379] <= 8'h10 ;
			data[76380] <= 8'h10 ;
			data[76381] <= 8'h10 ;
			data[76382] <= 8'h10 ;
			data[76383] <= 8'h10 ;
			data[76384] <= 8'h10 ;
			data[76385] <= 8'h10 ;
			data[76386] <= 8'h10 ;
			data[76387] <= 8'h10 ;
			data[76388] <= 8'h10 ;
			data[76389] <= 8'h10 ;
			data[76390] <= 8'h10 ;
			data[76391] <= 8'h10 ;
			data[76392] <= 8'h10 ;
			data[76393] <= 8'h10 ;
			data[76394] <= 8'h10 ;
			data[76395] <= 8'h10 ;
			data[76396] <= 8'h10 ;
			data[76397] <= 8'h10 ;
			data[76398] <= 8'h10 ;
			data[76399] <= 8'h10 ;
			data[76400] <= 8'h10 ;
			data[76401] <= 8'h10 ;
			data[76402] <= 8'h10 ;
			data[76403] <= 8'h10 ;
			data[76404] <= 8'h10 ;
			data[76405] <= 8'h10 ;
			data[76406] <= 8'h10 ;
			data[76407] <= 8'h10 ;
			data[76408] <= 8'h10 ;
			data[76409] <= 8'h10 ;
			data[76410] <= 8'h10 ;
			data[76411] <= 8'h10 ;
			data[76412] <= 8'h10 ;
			data[76413] <= 8'h10 ;
			data[76414] <= 8'h10 ;
			data[76415] <= 8'h10 ;
			data[76416] <= 8'h10 ;
			data[76417] <= 8'h10 ;
			data[76418] <= 8'h10 ;
			data[76419] <= 8'h10 ;
			data[76420] <= 8'h10 ;
			data[76421] <= 8'h10 ;
			data[76422] <= 8'h10 ;
			data[76423] <= 8'h10 ;
			data[76424] <= 8'h10 ;
			data[76425] <= 8'h10 ;
			data[76426] <= 8'h10 ;
			data[76427] <= 8'h10 ;
			data[76428] <= 8'h10 ;
			data[76429] <= 8'h10 ;
			data[76430] <= 8'h10 ;
			data[76431] <= 8'h10 ;
			data[76432] <= 8'h10 ;
			data[76433] <= 8'h10 ;
			data[76434] <= 8'h10 ;
			data[76435] <= 8'h10 ;
			data[76436] <= 8'h10 ;
			data[76437] <= 8'h10 ;
			data[76438] <= 8'h10 ;
			data[76439] <= 8'h10 ;
			data[76440] <= 8'h10 ;
			data[76441] <= 8'h10 ;
			data[76442] <= 8'h10 ;
			data[76443] <= 8'h10 ;
			data[76444] <= 8'h10 ;
			data[76445] <= 8'h10 ;
			data[76446] <= 8'h10 ;
			data[76447] <= 8'h10 ;
			data[76448] <= 8'h10 ;
			data[76449] <= 8'h10 ;
			data[76450] <= 8'h10 ;
			data[76451] <= 8'h10 ;
			data[76452] <= 8'h10 ;
			data[76453] <= 8'h10 ;
			data[76454] <= 8'h10 ;
			data[76455] <= 8'h10 ;
			data[76456] <= 8'h10 ;
			data[76457] <= 8'h10 ;
			data[76458] <= 8'h10 ;
			data[76459] <= 8'h10 ;
			data[76460] <= 8'h10 ;
			data[76461] <= 8'h10 ;
			data[76462] <= 8'h10 ;
			data[76463] <= 8'h10 ;
			data[76464] <= 8'h10 ;
			data[76465] <= 8'h10 ;
			data[76466] <= 8'h10 ;
			data[76467] <= 8'h10 ;
			data[76468] <= 8'h10 ;
			data[76469] <= 8'h10 ;
			data[76470] <= 8'h10 ;
			data[76471] <= 8'h10 ;
			data[76472] <= 8'h10 ;
			data[76473] <= 8'h10 ;
			data[76474] <= 8'h10 ;
			data[76475] <= 8'h10 ;
			data[76476] <= 8'h10 ;
			data[76477] <= 8'h10 ;
			data[76478] <= 8'h10 ;
			data[76479] <= 8'h10 ;
			data[76480] <= 8'h10 ;
			data[76481] <= 8'h10 ;
			data[76482] <= 8'h10 ;
			data[76483] <= 8'h10 ;
			data[76484] <= 8'h10 ;
			data[76485] <= 8'h10 ;
			data[76486] <= 8'h10 ;
			data[76487] <= 8'h10 ;
			data[76488] <= 8'h10 ;
			data[76489] <= 8'h10 ;
			data[76490] <= 8'h10 ;
			data[76491] <= 8'h10 ;
			data[76492] <= 8'h10 ;
			data[76493] <= 8'h10 ;
			data[76494] <= 8'h10 ;
			data[76495] <= 8'h10 ;
			data[76496] <= 8'h10 ;
			data[76497] <= 8'h10 ;
			data[76498] <= 8'h10 ;
			data[76499] <= 8'h10 ;
			data[76500] <= 8'h10 ;
			data[76501] <= 8'h10 ;
			data[76502] <= 8'h10 ;
			data[76503] <= 8'h10 ;
			data[76504] <= 8'h10 ;
			data[76505] <= 8'h10 ;
			data[76506] <= 8'h10 ;
			data[76507] <= 8'h10 ;
			data[76508] <= 8'h10 ;
			data[76509] <= 8'h10 ;
			data[76510] <= 8'h10 ;
			data[76511] <= 8'h10 ;
			data[76512] <= 8'h10 ;
			data[76513] <= 8'h10 ;
			data[76514] <= 8'h10 ;
			data[76515] <= 8'h10 ;
			data[76516] <= 8'h10 ;
			data[76517] <= 8'h10 ;
			data[76518] <= 8'h10 ;
			data[76519] <= 8'h10 ;
			data[76520] <= 8'h10 ;
			data[76521] <= 8'h10 ;
			data[76522] <= 8'h10 ;
			data[76523] <= 8'h10 ;
			data[76524] <= 8'h10 ;
			data[76525] <= 8'h10 ;
			data[76526] <= 8'h10 ;
			data[76527] <= 8'h10 ;
			data[76528] <= 8'h10 ;
			data[76529] <= 8'h10 ;
			data[76530] <= 8'h10 ;
			data[76531] <= 8'h10 ;
			data[76532] <= 8'h10 ;
			data[76533] <= 8'h10 ;
			data[76534] <= 8'h10 ;
			data[76535] <= 8'h10 ;
			data[76536] <= 8'h10 ;
			data[76537] <= 8'h10 ;
			data[76538] <= 8'h10 ;
			data[76539] <= 8'h10 ;
			data[76540] <= 8'h10 ;
			data[76541] <= 8'h10 ;
			data[76542] <= 8'h10 ;
			data[76543] <= 8'h10 ;
			data[76544] <= 8'h10 ;
			data[76545] <= 8'h10 ;
			data[76546] <= 8'h10 ;
			data[76547] <= 8'h10 ;
			data[76548] <= 8'h10 ;
			data[76549] <= 8'h10 ;
			data[76550] <= 8'h10 ;
			data[76551] <= 8'h10 ;
			data[76552] <= 8'h10 ;
			data[76553] <= 8'h10 ;
			data[76554] <= 8'h10 ;
			data[76555] <= 8'h10 ;
			data[76556] <= 8'h10 ;
			data[76557] <= 8'h10 ;
			data[76558] <= 8'h10 ;
			data[76559] <= 8'h10 ;
			data[76560] <= 8'h10 ;
			data[76561] <= 8'h10 ;
			data[76562] <= 8'h10 ;
			data[76563] <= 8'h10 ;
			data[76564] <= 8'h10 ;
			data[76565] <= 8'h10 ;
			data[76566] <= 8'h10 ;
			data[76567] <= 8'h10 ;
			data[76568] <= 8'h10 ;
			data[76569] <= 8'h10 ;
			data[76570] <= 8'h10 ;
			data[76571] <= 8'h10 ;
			data[76572] <= 8'h10 ;
			data[76573] <= 8'h10 ;
			data[76574] <= 8'h10 ;
			data[76575] <= 8'h10 ;
			data[76576] <= 8'h10 ;
			data[76577] <= 8'h10 ;
			data[76578] <= 8'h10 ;
			data[76579] <= 8'h10 ;
			data[76580] <= 8'h10 ;
			data[76581] <= 8'h10 ;
			data[76582] <= 8'h10 ;
			data[76583] <= 8'h10 ;
			data[76584] <= 8'h10 ;
			data[76585] <= 8'h10 ;
			data[76586] <= 8'h10 ;
			data[76587] <= 8'h10 ;
			data[76588] <= 8'h10 ;
			data[76589] <= 8'h10 ;
			data[76590] <= 8'h10 ;
			data[76591] <= 8'h10 ;
			data[76592] <= 8'h10 ;
			data[76593] <= 8'h10 ;
			data[76594] <= 8'h10 ;
			data[76595] <= 8'h10 ;
			data[76596] <= 8'h10 ;
			data[76597] <= 8'h10 ;
			data[76598] <= 8'h10 ;
			data[76599] <= 8'h10 ;
			data[76600] <= 8'h10 ;
			data[76601] <= 8'h10 ;
			data[76602] <= 8'h10 ;
			data[76603] <= 8'h10 ;
			data[76604] <= 8'h10 ;
			data[76605] <= 8'h10 ;
			data[76606] <= 8'h10 ;
			data[76607] <= 8'h10 ;
			data[76608] <= 8'h10 ;
			data[76609] <= 8'h10 ;
			data[76610] <= 8'h10 ;
			data[76611] <= 8'h10 ;
			data[76612] <= 8'h10 ;
			data[76613] <= 8'h10 ;
			data[76614] <= 8'h10 ;
			data[76615] <= 8'h10 ;
			data[76616] <= 8'h10 ;
			data[76617] <= 8'h10 ;
			data[76618] <= 8'h10 ;
			data[76619] <= 8'h10 ;
			data[76620] <= 8'h10 ;
			data[76621] <= 8'h10 ;
			data[76622] <= 8'h10 ;
			data[76623] <= 8'h10 ;
			data[76624] <= 8'h10 ;
			data[76625] <= 8'h10 ;
			data[76626] <= 8'h10 ;
			data[76627] <= 8'h10 ;
			data[76628] <= 8'h10 ;
			data[76629] <= 8'h10 ;
			data[76630] <= 8'h10 ;
			data[76631] <= 8'h10 ;
			data[76632] <= 8'h10 ;
			data[76633] <= 8'h10 ;
			data[76634] <= 8'h10 ;
			data[76635] <= 8'h10 ;
			data[76636] <= 8'h10 ;
			data[76637] <= 8'h10 ;
			data[76638] <= 8'h10 ;
			data[76639] <= 8'h10 ;
			data[76640] <= 8'h10 ;
			data[76641] <= 8'h10 ;
			data[76642] <= 8'h10 ;
			data[76643] <= 8'h10 ;
			data[76644] <= 8'h10 ;
			data[76645] <= 8'h10 ;
			data[76646] <= 8'h10 ;
			data[76647] <= 8'h10 ;
			data[76648] <= 8'h10 ;
			data[76649] <= 8'h10 ;
			data[76650] <= 8'h10 ;
			data[76651] <= 8'h10 ;
			data[76652] <= 8'h10 ;
			data[76653] <= 8'h10 ;
			data[76654] <= 8'h10 ;
			data[76655] <= 8'h10 ;
			data[76656] <= 8'h10 ;
			data[76657] <= 8'h10 ;
			data[76658] <= 8'h10 ;
			data[76659] <= 8'h10 ;
			data[76660] <= 8'h10 ;
			data[76661] <= 8'h10 ;
			data[76662] <= 8'h10 ;
			data[76663] <= 8'h10 ;
			data[76664] <= 8'h10 ;
			data[76665] <= 8'h10 ;
			data[76666] <= 8'h10 ;
			data[76667] <= 8'h10 ;
			data[76668] <= 8'h10 ;
			data[76669] <= 8'h10 ;
			data[76670] <= 8'h10 ;
			data[76671] <= 8'h10 ;
			data[76672] <= 8'h10 ;
			data[76673] <= 8'h10 ;
			data[76674] <= 8'h10 ;
			data[76675] <= 8'h10 ;
			data[76676] <= 8'h10 ;
			data[76677] <= 8'h10 ;
			data[76678] <= 8'h10 ;
			data[76679] <= 8'h10 ;
			data[76680] <= 8'h10 ;
			data[76681] <= 8'h10 ;
			data[76682] <= 8'h10 ;
			data[76683] <= 8'h10 ;
			data[76684] <= 8'h10 ;
			data[76685] <= 8'h10 ;
			data[76686] <= 8'h10 ;
			data[76687] <= 8'h10 ;
			data[76688] <= 8'h10 ;
			data[76689] <= 8'h10 ;
			data[76690] <= 8'h10 ;
			data[76691] <= 8'h10 ;
			data[76692] <= 8'h10 ;
			data[76693] <= 8'h10 ;
			data[76694] <= 8'h10 ;
			data[76695] <= 8'h10 ;
			data[76696] <= 8'h10 ;
			data[76697] <= 8'h10 ;
			data[76698] <= 8'h10 ;
			data[76699] <= 8'h10 ;
			data[76700] <= 8'h10 ;
			data[76701] <= 8'h10 ;
			data[76702] <= 8'h10 ;
			data[76703] <= 8'h10 ;
			data[76704] <= 8'h10 ;
			data[76705] <= 8'h10 ;
			data[76706] <= 8'h10 ;
			data[76707] <= 8'h10 ;
			data[76708] <= 8'h10 ;
			data[76709] <= 8'h10 ;
			data[76710] <= 8'h10 ;
			data[76711] <= 8'h10 ;
			data[76712] <= 8'h10 ;
			data[76713] <= 8'h10 ;
			data[76714] <= 8'h10 ;
			data[76715] <= 8'h10 ;
			data[76716] <= 8'h10 ;
			data[76717] <= 8'h10 ;
			data[76718] <= 8'h10 ;
			data[76719] <= 8'h10 ;
			data[76720] <= 8'h10 ;
			data[76721] <= 8'h10 ;
			data[76722] <= 8'h10 ;
			data[76723] <= 8'h10 ;
			data[76724] <= 8'h10 ;
			data[76725] <= 8'h10 ;
			data[76726] <= 8'h10 ;
			data[76727] <= 8'h10 ;
			data[76728] <= 8'h10 ;
			data[76729] <= 8'h10 ;
			data[76730] <= 8'h10 ;
			data[76731] <= 8'h10 ;
			data[76732] <= 8'h10 ;
			data[76733] <= 8'h10 ;
			data[76734] <= 8'h10 ;
			data[76735] <= 8'h10 ;
			data[76736] <= 8'h10 ;
			data[76737] <= 8'h10 ;
			data[76738] <= 8'h10 ;
			data[76739] <= 8'h10 ;
			data[76740] <= 8'h10 ;
			data[76741] <= 8'h10 ;
			data[76742] <= 8'h10 ;
			data[76743] <= 8'h10 ;
			data[76744] <= 8'h10 ;
			data[76745] <= 8'h10 ;
			data[76746] <= 8'h10 ;
			data[76747] <= 8'h10 ;
			data[76748] <= 8'h10 ;
			data[76749] <= 8'h10 ;
			data[76750] <= 8'h10 ;
			data[76751] <= 8'h10 ;
			data[76752] <= 8'h10 ;
			data[76753] <= 8'h10 ;
			data[76754] <= 8'h10 ;
			data[76755] <= 8'h10 ;
			data[76756] <= 8'h10 ;
			data[76757] <= 8'h10 ;
			data[76758] <= 8'h10 ;
			data[76759] <= 8'h10 ;
			data[76760] <= 8'h10 ;
			data[76761] <= 8'h10 ;
			data[76762] <= 8'h10 ;
			data[76763] <= 8'h10 ;
			data[76764] <= 8'h10 ;
			data[76765] <= 8'h10 ;
			data[76766] <= 8'h10 ;
			data[76767] <= 8'h10 ;
			data[76768] <= 8'h10 ;
			data[76769] <= 8'h10 ;
			data[76770] <= 8'h10 ;
			data[76771] <= 8'h10 ;
			data[76772] <= 8'h10 ;
			data[76773] <= 8'h10 ;
			data[76774] <= 8'h10 ;
			data[76775] <= 8'h10 ;
			data[76776] <= 8'h10 ;
			data[76777] <= 8'h10 ;
			data[76778] <= 8'h10 ;
			data[76779] <= 8'h10 ;
			data[76780] <= 8'h10 ;
			data[76781] <= 8'h10 ;
			data[76782] <= 8'h10 ;
			data[76783] <= 8'h10 ;
			data[76784] <= 8'h10 ;
			data[76785] <= 8'h10 ;
			data[76786] <= 8'h10 ;
			data[76787] <= 8'h10 ;
			data[76788] <= 8'h10 ;
			data[76789] <= 8'h10 ;
			data[76790] <= 8'h10 ;
			data[76791] <= 8'h10 ;
			data[76792] <= 8'h10 ;
			data[76793] <= 8'h10 ;
			data[76794] <= 8'h10 ;
			data[76795] <= 8'h10 ;
			data[76796] <= 8'h10 ;
			data[76797] <= 8'h10 ;
			data[76798] <= 8'h10 ;
			data[76799] <= 8'h10 ;
			data[76800] <= 8'h10 ;
			data[76801] <= 8'h10 ;
			data[76802] <= 8'h10 ;
			data[76803] <= 8'h10 ;
			data[76804] <= 8'h10 ;
			data[76805] <= 8'h10 ;
			data[76806] <= 8'h10 ;
			data[76807] <= 8'h10 ;
			data[76808] <= 8'h10 ;
			data[76809] <= 8'h10 ;
			data[76810] <= 8'h10 ;
			data[76811] <= 8'h10 ;
			data[76812] <= 8'h10 ;
			data[76813] <= 8'h10 ;
			data[76814] <= 8'h10 ;
			data[76815] <= 8'h10 ;
			data[76816] <= 8'h10 ;
			data[76817] <= 8'h10 ;
			data[76818] <= 8'h10 ;
			data[76819] <= 8'h10 ;
			data[76820] <= 8'h10 ;
			data[76821] <= 8'h10 ;
			data[76822] <= 8'h10 ;
			data[76823] <= 8'h10 ;
			data[76824] <= 8'h10 ;
			data[76825] <= 8'h10 ;
			data[76826] <= 8'h10 ;
			data[76827] <= 8'h10 ;
			data[76828] <= 8'h10 ;
			data[76829] <= 8'h10 ;
			data[76830] <= 8'h10 ;
			data[76831] <= 8'h10 ;
			data[76832] <= 8'h10 ;
			data[76833] <= 8'h10 ;
			data[76834] <= 8'h10 ;
			data[76835] <= 8'h10 ;
			data[76836] <= 8'h10 ;
			data[76837] <= 8'h10 ;
			data[76838] <= 8'h10 ;
			data[76839] <= 8'h10 ;
			data[76840] <= 8'h10 ;
			data[76841] <= 8'h10 ;
			data[76842] <= 8'h10 ;
			data[76843] <= 8'h10 ;
			data[76844] <= 8'h10 ;
			data[76845] <= 8'h10 ;
			data[76846] <= 8'h10 ;
			data[76847] <= 8'h10 ;
			data[76848] <= 8'h10 ;
			data[76849] <= 8'h10 ;
			data[76850] <= 8'h10 ;
			data[76851] <= 8'h10 ;
			data[76852] <= 8'h10 ;
			data[76853] <= 8'h10 ;
			data[76854] <= 8'h10 ;
			data[76855] <= 8'h10 ;
			data[76856] <= 8'h10 ;
			data[76857] <= 8'h10 ;
			data[76858] <= 8'h10 ;
			data[76859] <= 8'h10 ;
			data[76860] <= 8'h10 ;
			data[76861] <= 8'h10 ;
			data[76862] <= 8'h10 ;
			data[76863] <= 8'h10 ;
			data[76864] <= 8'h10 ;
			data[76865] <= 8'h10 ;
			data[76866] <= 8'h10 ;
			data[76867] <= 8'h10 ;
			data[76868] <= 8'h10 ;
			data[76869] <= 8'h10 ;
			data[76870] <= 8'h10 ;
			data[76871] <= 8'h10 ;
			data[76872] <= 8'h10 ;
			data[76873] <= 8'h10 ;
			data[76874] <= 8'h10 ;
			data[76875] <= 8'h10 ;
			data[76876] <= 8'h10 ;
			data[76877] <= 8'h10 ;
			data[76878] <= 8'h10 ;
			data[76879] <= 8'h10 ;
			data[76880] <= 8'h10 ;
			data[76881] <= 8'h10 ;
			data[76882] <= 8'h10 ;
			data[76883] <= 8'h10 ;
			data[76884] <= 8'h10 ;
			data[76885] <= 8'h10 ;
			data[76886] <= 8'h10 ;
			data[76887] <= 8'h10 ;
			data[76888] <= 8'h10 ;
			data[76889] <= 8'h10 ;
			data[76890] <= 8'h10 ;
			data[76891] <= 8'h10 ;
			data[76892] <= 8'h10 ;
			data[76893] <= 8'h10 ;
			data[76894] <= 8'h10 ;
			data[76895] <= 8'h10 ;
			data[76896] <= 8'h10 ;
			data[76897] <= 8'h10 ;
			data[76898] <= 8'h10 ;
			data[76899] <= 8'h10 ;
			data[76900] <= 8'h10 ;
			data[76901] <= 8'h10 ;
			data[76902] <= 8'h10 ;
			data[76903] <= 8'h10 ;
			data[76904] <= 8'h10 ;
			data[76905] <= 8'h10 ;
			data[76906] <= 8'h10 ;
			data[76907] <= 8'h10 ;
			data[76908] <= 8'h10 ;
			data[76909] <= 8'h10 ;
			data[76910] <= 8'h10 ;
			data[76911] <= 8'h10 ;
			data[76912] <= 8'h10 ;
			data[76913] <= 8'h10 ;
			data[76914] <= 8'h10 ;
			data[76915] <= 8'h10 ;
			data[76916] <= 8'h10 ;
			data[76917] <= 8'h10 ;
			data[76918] <= 8'h10 ;
			data[76919] <= 8'h10 ;
			data[76920] <= 8'h10 ;
			data[76921] <= 8'h10 ;
			data[76922] <= 8'h10 ;
			data[76923] <= 8'h10 ;
			data[76924] <= 8'h10 ;
			data[76925] <= 8'h10 ;
			data[76926] <= 8'h10 ;
			data[76927] <= 8'h10 ;
			data[76928] <= 8'h10 ;
			data[76929] <= 8'h10 ;
			data[76930] <= 8'h10 ;
			data[76931] <= 8'h10 ;
			data[76932] <= 8'h10 ;
			data[76933] <= 8'h10 ;
			data[76934] <= 8'h10 ;
			data[76935] <= 8'h10 ;
			data[76936] <= 8'h10 ;
			data[76937] <= 8'h10 ;
			data[76938] <= 8'h10 ;
			data[76939] <= 8'h10 ;
			data[76940] <= 8'h10 ;
			data[76941] <= 8'h10 ;
			data[76942] <= 8'h10 ;
			data[76943] <= 8'h10 ;
			data[76944] <= 8'h10 ;
			data[76945] <= 8'h10 ;
			data[76946] <= 8'h10 ;
			data[76947] <= 8'h10 ;
			data[76948] <= 8'h10 ;
			data[76949] <= 8'h10 ;
			data[76950] <= 8'h10 ;
			data[76951] <= 8'h10 ;
			data[76952] <= 8'h10 ;
			data[76953] <= 8'h10 ;
			data[76954] <= 8'h10 ;
			data[76955] <= 8'h10 ;
			data[76956] <= 8'h10 ;
			data[76957] <= 8'h10 ;
			data[76958] <= 8'h10 ;
			data[76959] <= 8'h10 ;
			data[76960] <= 8'h10 ;
			data[76961] <= 8'h10 ;
			data[76962] <= 8'h10 ;
			data[76963] <= 8'h10 ;
			data[76964] <= 8'h10 ;
			data[76965] <= 8'h10 ;
			data[76966] <= 8'h10 ;
			data[76967] <= 8'h10 ;
			data[76968] <= 8'h10 ;
			data[76969] <= 8'h10 ;
			data[76970] <= 8'h10 ;
			data[76971] <= 8'h10 ;
			data[76972] <= 8'h10 ;
			data[76973] <= 8'h10 ;
			data[76974] <= 8'h10 ;
			data[76975] <= 8'h10 ;
			data[76976] <= 8'h10 ;
			data[76977] <= 8'h10 ;
			data[76978] <= 8'h10 ;
			data[76979] <= 8'h10 ;
			data[76980] <= 8'h10 ;
			data[76981] <= 8'h10 ;
			data[76982] <= 8'h10 ;
			data[76983] <= 8'h10 ;
			data[76984] <= 8'h10 ;
			data[76985] <= 8'h10 ;
			data[76986] <= 8'h10 ;
			data[76987] <= 8'h10 ;
			data[76988] <= 8'h10 ;
			data[76989] <= 8'h10 ;
			data[76990] <= 8'h10 ;
			data[76991] <= 8'h10 ;
			data[76992] <= 8'h10 ;
			data[76993] <= 8'h10 ;
			data[76994] <= 8'h10 ;
			data[76995] <= 8'h10 ;
			data[76996] <= 8'h10 ;
			data[76997] <= 8'h10 ;
			data[76998] <= 8'h10 ;
			data[76999] <= 8'h10 ;
			data[77000] <= 8'h10 ;
			data[77001] <= 8'h10 ;
			data[77002] <= 8'h10 ;
			data[77003] <= 8'h10 ;
			data[77004] <= 8'h10 ;
			data[77005] <= 8'h10 ;
			data[77006] <= 8'h10 ;
			data[77007] <= 8'h10 ;
			data[77008] <= 8'h10 ;
			data[77009] <= 8'h10 ;
			data[77010] <= 8'h10 ;
			data[77011] <= 8'h10 ;
			data[77012] <= 8'h10 ;
			data[77013] <= 8'h10 ;
			data[77014] <= 8'h10 ;
			data[77015] <= 8'h10 ;
			data[77016] <= 8'h10 ;
			data[77017] <= 8'h10 ;
			data[77018] <= 8'h10 ;
			data[77019] <= 8'h10 ;
			data[77020] <= 8'h10 ;
			data[77021] <= 8'h10 ;
			data[77022] <= 8'h10 ;
			data[77023] <= 8'h10 ;
			data[77024] <= 8'h10 ;
			data[77025] <= 8'h10 ;
			data[77026] <= 8'h10 ;
			data[77027] <= 8'h10 ;
			data[77028] <= 8'h10 ;
			data[77029] <= 8'h10 ;
			data[77030] <= 8'h10 ;
			data[77031] <= 8'h10 ;
			data[77032] <= 8'h10 ;
			data[77033] <= 8'h10 ;
			data[77034] <= 8'h10 ;
			data[77035] <= 8'h10 ;
			data[77036] <= 8'h10 ;
			data[77037] <= 8'h10 ;
			data[77038] <= 8'h10 ;
			data[77039] <= 8'h10 ;
			data[77040] <= 8'h10 ;
			data[77041] <= 8'h10 ;
			data[77042] <= 8'h10 ;
			data[77043] <= 8'h10 ;
			data[77044] <= 8'h10 ;
			data[77045] <= 8'h10 ;
			data[77046] <= 8'h10 ;
			data[77047] <= 8'h10 ;
			data[77048] <= 8'h10 ;
			data[77049] <= 8'h10 ;
			data[77050] <= 8'h10 ;
			data[77051] <= 8'h10 ;
			data[77052] <= 8'h10 ;
			data[77053] <= 8'h10 ;
			data[77054] <= 8'h10 ;
			data[77055] <= 8'h10 ;
			data[77056] <= 8'h10 ;
			data[77057] <= 8'h10 ;
			data[77058] <= 8'h10 ;
			data[77059] <= 8'h10 ;
			data[77060] <= 8'h10 ;
			data[77061] <= 8'h10 ;
			data[77062] <= 8'h10 ;
			data[77063] <= 8'h10 ;
			data[77064] <= 8'h10 ;
			data[77065] <= 8'h10 ;
			data[77066] <= 8'h10 ;
			data[77067] <= 8'h10 ;
			data[77068] <= 8'h10 ;
			data[77069] <= 8'h10 ;
			data[77070] <= 8'h10 ;
			data[77071] <= 8'h10 ;
			data[77072] <= 8'h10 ;
			data[77073] <= 8'h10 ;
			data[77074] <= 8'h10 ;
			data[77075] <= 8'h10 ;
			data[77076] <= 8'h10 ;
			data[77077] <= 8'h10 ;
			data[77078] <= 8'h10 ;
			data[77079] <= 8'h10 ;
			data[77080] <= 8'h10 ;
			data[77081] <= 8'h10 ;
			data[77082] <= 8'h10 ;
			data[77083] <= 8'h10 ;
			data[77084] <= 8'h10 ;
			data[77085] <= 8'h10 ;
			data[77086] <= 8'h10 ;
			data[77087] <= 8'h10 ;
			data[77088] <= 8'h10 ;
			data[77089] <= 8'h10 ;
			data[77090] <= 8'h10 ;
			data[77091] <= 8'h10 ;
			data[77092] <= 8'h10 ;
			data[77093] <= 8'h10 ;
			data[77094] <= 8'h10 ;
			data[77095] <= 8'h10 ;
			data[77096] <= 8'h10 ;
			data[77097] <= 8'h10 ;
			data[77098] <= 8'h10 ;
			data[77099] <= 8'h10 ;
			data[77100] <= 8'h10 ;
			data[77101] <= 8'h10 ;
			data[77102] <= 8'h10 ;
			data[77103] <= 8'h10 ;
			data[77104] <= 8'h10 ;
			data[77105] <= 8'h10 ;
			data[77106] <= 8'h10 ;
			data[77107] <= 8'h10 ;
			data[77108] <= 8'h10 ;
			data[77109] <= 8'h10 ;
			data[77110] <= 8'h10 ;
			data[77111] <= 8'h10 ;
			data[77112] <= 8'h10 ;
			data[77113] <= 8'h10 ;
			data[77114] <= 8'h10 ;
			data[77115] <= 8'h10 ;
			data[77116] <= 8'h10 ;
			data[77117] <= 8'h10 ;
			data[77118] <= 8'h10 ;
			data[77119] <= 8'h10 ;
			data[77120] <= 8'h10 ;
			data[77121] <= 8'h10 ;
			data[77122] <= 8'h10 ;
			data[77123] <= 8'h10 ;
			data[77124] <= 8'h10 ;
			data[77125] <= 8'h10 ;
			data[77126] <= 8'h10 ;
			data[77127] <= 8'h10 ;
			data[77128] <= 8'h10 ;
			data[77129] <= 8'h10 ;
			data[77130] <= 8'h10 ;
			data[77131] <= 8'h10 ;
			data[77132] <= 8'h10 ;
			data[77133] <= 8'h10 ;
			data[77134] <= 8'h10 ;
			data[77135] <= 8'h10 ;
			data[77136] <= 8'h10 ;
			data[77137] <= 8'h10 ;
			data[77138] <= 8'h10 ;
			data[77139] <= 8'h10 ;
			data[77140] <= 8'h10 ;
			data[77141] <= 8'h10 ;
			data[77142] <= 8'h10 ;
			data[77143] <= 8'h10 ;
			data[77144] <= 8'h10 ;
			data[77145] <= 8'h10 ;
			data[77146] <= 8'h10 ;
			data[77147] <= 8'h10 ;
			data[77148] <= 8'h10 ;
			data[77149] <= 8'h10 ;
			data[77150] <= 8'h10 ;
			data[77151] <= 8'h10 ;
			data[77152] <= 8'h10 ;
			data[77153] <= 8'h10 ;
			data[77154] <= 8'h10 ;
			data[77155] <= 8'h10 ;
			data[77156] <= 8'h10 ;
			data[77157] <= 8'h10 ;
			data[77158] <= 8'h10 ;
			data[77159] <= 8'h10 ;
			data[77160] <= 8'h10 ;
			data[77161] <= 8'h10 ;
			data[77162] <= 8'h10 ;
			data[77163] <= 8'h10 ;
			data[77164] <= 8'h10 ;
			data[77165] <= 8'h10 ;
			data[77166] <= 8'h10 ;
			data[77167] <= 8'h10 ;
			data[77168] <= 8'h10 ;
			data[77169] <= 8'h10 ;
			data[77170] <= 8'h10 ;
			data[77171] <= 8'h10 ;
			data[77172] <= 8'h10 ;
			data[77173] <= 8'h10 ;
			data[77174] <= 8'h10 ;
			data[77175] <= 8'h10 ;
			data[77176] <= 8'h10 ;
			data[77177] <= 8'h10 ;
			data[77178] <= 8'h10 ;
			data[77179] <= 8'h10 ;
			data[77180] <= 8'h10 ;
			data[77181] <= 8'h10 ;
			data[77182] <= 8'h10 ;
			data[77183] <= 8'h10 ;
			data[77184] <= 8'h10 ;
			data[77185] <= 8'h10 ;
			data[77186] <= 8'h10 ;
			data[77187] <= 8'h10 ;
			data[77188] <= 8'h10 ;
			data[77189] <= 8'h10 ;
			data[77190] <= 8'h10 ;
			data[77191] <= 8'h10 ;
			data[77192] <= 8'h10 ;
			data[77193] <= 8'h10 ;
			data[77194] <= 8'h10 ;
			data[77195] <= 8'h10 ;
			data[77196] <= 8'h10 ;
			data[77197] <= 8'h10 ;
			data[77198] <= 8'h10 ;
			data[77199] <= 8'h10 ;
			data[77200] <= 8'h10 ;
			data[77201] <= 8'h10 ;
			data[77202] <= 8'h10 ;
			data[77203] <= 8'h10 ;
			data[77204] <= 8'h10 ;
			data[77205] <= 8'h10 ;
			data[77206] <= 8'h10 ;
			data[77207] <= 8'h10 ;
			data[77208] <= 8'h10 ;
			data[77209] <= 8'h10 ;
			data[77210] <= 8'h10 ;
			data[77211] <= 8'h10 ;
			data[77212] <= 8'h10 ;
			data[77213] <= 8'h10 ;
			data[77214] <= 8'h10 ;
			data[77215] <= 8'h10 ;
			data[77216] <= 8'h10 ;
			data[77217] <= 8'h10 ;
			data[77218] <= 8'h10 ;
			data[77219] <= 8'h10 ;
			data[77220] <= 8'h10 ;
			data[77221] <= 8'h10 ;
			data[77222] <= 8'h10 ;
			data[77223] <= 8'h10 ;
			data[77224] <= 8'h10 ;
			data[77225] <= 8'h10 ;
			data[77226] <= 8'h10 ;
			data[77227] <= 8'h10 ;
			data[77228] <= 8'h10 ;
			data[77229] <= 8'h10 ;
			data[77230] <= 8'h10 ;
			data[77231] <= 8'h10 ;
			data[77232] <= 8'h10 ;
			data[77233] <= 8'h10 ;
			data[77234] <= 8'h10 ;
			data[77235] <= 8'h10 ;
			data[77236] <= 8'h10 ;
			data[77237] <= 8'h10 ;
			data[77238] <= 8'h10 ;
			data[77239] <= 8'h10 ;
			data[77240] <= 8'h10 ;
			data[77241] <= 8'h10 ;
			data[77242] <= 8'h10 ;
			data[77243] <= 8'h10 ;
			data[77244] <= 8'h10 ;
			data[77245] <= 8'h10 ;
			data[77246] <= 8'h10 ;
			data[77247] <= 8'h10 ;
			data[77248] <= 8'h10 ;
			data[77249] <= 8'h10 ;
			data[77250] <= 8'h10 ;
			data[77251] <= 8'h10 ;
			data[77252] <= 8'h10 ;
			data[77253] <= 8'h10 ;
			data[77254] <= 8'h10 ;
			data[77255] <= 8'h10 ;
			data[77256] <= 8'h10 ;
			data[77257] <= 8'h10 ;
			data[77258] <= 8'h10 ;
			data[77259] <= 8'h10 ;
			data[77260] <= 8'h10 ;
			data[77261] <= 8'h10 ;
			data[77262] <= 8'h10 ;
			data[77263] <= 8'h10 ;
			data[77264] <= 8'h10 ;
			data[77265] <= 8'h10 ;
			data[77266] <= 8'h10 ;
			data[77267] <= 8'h10 ;
			data[77268] <= 8'h10 ;
			data[77269] <= 8'h10 ;
			data[77270] <= 8'h10 ;
			data[77271] <= 8'h10 ;
			data[77272] <= 8'h10 ;
			data[77273] <= 8'h10 ;
			data[77274] <= 8'h10 ;
			data[77275] <= 8'h10 ;
			data[77276] <= 8'h10 ;
			data[77277] <= 8'h10 ;
			data[77278] <= 8'h10 ;
			data[77279] <= 8'h10 ;
			data[77280] <= 8'h10 ;
			data[77281] <= 8'h10 ;
			data[77282] <= 8'h10 ;
			data[77283] <= 8'h10 ;
			data[77284] <= 8'h10 ;
			data[77285] <= 8'h10 ;
			data[77286] <= 8'h10 ;
			data[77287] <= 8'h10 ;
			data[77288] <= 8'h10 ;
			data[77289] <= 8'h10 ;
			data[77290] <= 8'h10 ;
			data[77291] <= 8'h10 ;
			data[77292] <= 8'h10 ;
			data[77293] <= 8'h10 ;
			data[77294] <= 8'h10 ;
			data[77295] <= 8'h10 ;
			data[77296] <= 8'h10 ;
			data[77297] <= 8'h10 ;
			data[77298] <= 8'h10 ;
			data[77299] <= 8'h10 ;
			data[77300] <= 8'h10 ;
			data[77301] <= 8'h10 ;
			data[77302] <= 8'h10 ;
			data[77303] <= 8'h10 ;
			data[77304] <= 8'h10 ;
			data[77305] <= 8'h10 ;
			data[77306] <= 8'h10 ;
			data[77307] <= 8'h10 ;
			data[77308] <= 8'h10 ;
			data[77309] <= 8'h10 ;
			data[77310] <= 8'h10 ;
			data[77311] <= 8'h10 ;
			data[77312] <= 8'h10 ;
			data[77313] <= 8'h10 ;
			data[77314] <= 8'h10 ;
			data[77315] <= 8'h10 ;
			data[77316] <= 8'h10 ;
			data[77317] <= 8'h10 ;
			data[77318] <= 8'h10 ;
			data[77319] <= 8'h10 ;
			data[77320] <= 8'h10 ;
			data[77321] <= 8'h10 ;
			data[77322] <= 8'h10 ;
			data[77323] <= 8'h10 ;
			data[77324] <= 8'h10 ;
			data[77325] <= 8'h10 ;
			data[77326] <= 8'h10 ;
			data[77327] <= 8'h10 ;
			data[77328] <= 8'h10 ;
			data[77329] <= 8'h10 ;
			data[77330] <= 8'h10 ;
			data[77331] <= 8'h10 ;
			data[77332] <= 8'h10 ;
			data[77333] <= 8'h10 ;
			data[77334] <= 8'h10 ;
			data[77335] <= 8'h10 ;
			data[77336] <= 8'h10 ;
			data[77337] <= 8'h10 ;
			data[77338] <= 8'h10 ;
			data[77339] <= 8'h10 ;
			data[77340] <= 8'h10 ;
			data[77341] <= 8'h10 ;
			data[77342] <= 8'h10 ;
			data[77343] <= 8'h10 ;
			data[77344] <= 8'h10 ;
			data[77345] <= 8'h10 ;
			data[77346] <= 8'h10 ;
			data[77347] <= 8'h10 ;
			data[77348] <= 8'h10 ;
			data[77349] <= 8'h10 ;
			data[77350] <= 8'h10 ;
			data[77351] <= 8'h10 ;
			data[77352] <= 8'h10 ;
			data[77353] <= 8'h10 ;
			data[77354] <= 8'h10 ;
			data[77355] <= 8'h10 ;
			data[77356] <= 8'h10 ;
			data[77357] <= 8'h10 ;
			data[77358] <= 8'h10 ;
			data[77359] <= 8'h10 ;
			data[77360] <= 8'h10 ;
			data[77361] <= 8'h10 ;
			data[77362] <= 8'h10 ;
			data[77363] <= 8'h10 ;
			data[77364] <= 8'h10 ;
			data[77365] <= 8'h10 ;
			data[77366] <= 8'h10 ;
			data[77367] <= 8'h10 ;
			data[77368] <= 8'h10 ;
			data[77369] <= 8'h10 ;
			data[77370] <= 8'h10 ;
			data[77371] <= 8'h10 ;
			data[77372] <= 8'h10 ;
			data[77373] <= 8'h10 ;
			data[77374] <= 8'h10 ;
			data[77375] <= 8'h10 ;
			data[77376] <= 8'h10 ;
			data[77377] <= 8'h10 ;
			data[77378] <= 8'h10 ;
			data[77379] <= 8'h10 ;
			data[77380] <= 8'h10 ;
			data[77381] <= 8'h10 ;
			data[77382] <= 8'h10 ;
			data[77383] <= 8'h10 ;
			data[77384] <= 8'h10 ;
			data[77385] <= 8'h10 ;
			data[77386] <= 8'h10 ;
			data[77387] <= 8'h10 ;
			data[77388] <= 8'h10 ;
			data[77389] <= 8'h10 ;
			data[77390] <= 8'h10 ;
			data[77391] <= 8'h10 ;
			data[77392] <= 8'h10 ;
			data[77393] <= 8'h10 ;
			data[77394] <= 8'h10 ;
			data[77395] <= 8'h10 ;
			data[77396] <= 8'h10 ;
			data[77397] <= 8'h10 ;
			data[77398] <= 8'h10 ;
			data[77399] <= 8'h10 ;
			data[77400] <= 8'h10 ;
			data[77401] <= 8'h10 ;
			data[77402] <= 8'h10 ;
			data[77403] <= 8'h10 ;
			data[77404] <= 8'h10 ;
			data[77405] <= 8'h10 ;
			data[77406] <= 8'h10 ;
			data[77407] <= 8'h10 ;
			data[77408] <= 8'h10 ;
			data[77409] <= 8'h10 ;
			data[77410] <= 8'h10 ;
			data[77411] <= 8'h10 ;
			data[77412] <= 8'h10 ;
			data[77413] <= 8'h10 ;
			data[77414] <= 8'h10 ;
			data[77415] <= 8'h10 ;
			data[77416] <= 8'h10 ;
			data[77417] <= 8'h10 ;
			data[77418] <= 8'h10 ;
			data[77419] <= 8'h10 ;
			data[77420] <= 8'h10 ;
			data[77421] <= 8'h10 ;
			data[77422] <= 8'h10 ;
			data[77423] <= 8'h10 ;
			data[77424] <= 8'h10 ;
			data[77425] <= 8'h10 ;
			data[77426] <= 8'h10 ;
			data[77427] <= 8'h10 ;
			data[77428] <= 8'h10 ;
			data[77429] <= 8'h10 ;
			data[77430] <= 8'h10 ;
			data[77431] <= 8'h10 ;
			data[77432] <= 8'h10 ;
			data[77433] <= 8'h10 ;
			data[77434] <= 8'h10 ;
			data[77435] <= 8'h10 ;
			data[77436] <= 8'h10 ;
			data[77437] <= 8'h10 ;
			data[77438] <= 8'h10 ;
			data[77439] <= 8'h10 ;
			data[77440] <= 8'h10 ;
			data[77441] <= 8'h10 ;
			data[77442] <= 8'h10 ;
			data[77443] <= 8'h10 ;
			data[77444] <= 8'h10 ;
			data[77445] <= 8'h10 ;
			data[77446] <= 8'h10 ;
			data[77447] <= 8'h10 ;
			data[77448] <= 8'h10 ;
			data[77449] <= 8'h10 ;
			data[77450] <= 8'h10 ;
			data[77451] <= 8'h10 ;
			data[77452] <= 8'h10 ;
			data[77453] <= 8'h10 ;
			data[77454] <= 8'h10 ;
			data[77455] <= 8'h10 ;
			data[77456] <= 8'h10 ;
			data[77457] <= 8'h10 ;
			data[77458] <= 8'h10 ;
			data[77459] <= 8'h10 ;
			data[77460] <= 8'h10 ;
			data[77461] <= 8'h10 ;
			data[77462] <= 8'h10 ;
			data[77463] <= 8'h10 ;
			data[77464] <= 8'h10 ;
			data[77465] <= 8'h10 ;
			data[77466] <= 8'h10 ;
			data[77467] <= 8'h10 ;
			data[77468] <= 8'h10 ;
			data[77469] <= 8'h10 ;
			data[77470] <= 8'h10 ;
			data[77471] <= 8'h10 ;
			data[77472] <= 8'h10 ;
			data[77473] <= 8'h10 ;
			data[77474] <= 8'h10 ;
			data[77475] <= 8'h10 ;
			data[77476] <= 8'h10 ;
			data[77477] <= 8'h10 ;
			data[77478] <= 8'h10 ;
			data[77479] <= 8'h10 ;
			data[77480] <= 8'h10 ;
			data[77481] <= 8'h10 ;
			data[77482] <= 8'h10 ;
			data[77483] <= 8'h10 ;
			data[77484] <= 8'h10 ;
			data[77485] <= 8'h10 ;
			data[77486] <= 8'h10 ;
			data[77487] <= 8'h10 ;
			data[77488] <= 8'h10 ;
			data[77489] <= 8'h10 ;
			data[77490] <= 8'h10 ;
			data[77491] <= 8'h10 ;
			data[77492] <= 8'h10 ;
			data[77493] <= 8'h10 ;
			data[77494] <= 8'h10 ;
			data[77495] <= 8'h10 ;
			data[77496] <= 8'h10 ;
			data[77497] <= 8'h10 ;
			data[77498] <= 8'h10 ;
			data[77499] <= 8'h10 ;
			data[77500] <= 8'h10 ;
			data[77501] <= 8'h10 ;
			data[77502] <= 8'h10 ;
			data[77503] <= 8'h10 ;
			data[77504] <= 8'h10 ;
			data[77505] <= 8'h10 ;
			data[77506] <= 8'h10 ;
			data[77507] <= 8'h10 ;
			data[77508] <= 8'h10 ;
			data[77509] <= 8'h10 ;
			data[77510] <= 8'h10 ;
			data[77511] <= 8'h10 ;
			data[77512] <= 8'h10 ;
			data[77513] <= 8'h10 ;
			data[77514] <= 8'h10 ;
			data[77515] <= 8'h10 ;
			data[77516] <= 8'h10 ;
			data[77517] <= 8'h10 ;
			data[77518] <= 8'h10 ;
			data[77519] <= 8'h10 ;
			data[77520] <= 8'h10 ;
			data[77521] <= 8'h10 ;
			data[77522] <= 8'h10 ;
			data[77523] <= 8'h10 ;
			data[77524] <= 8'h10 ;
			data[77525] <= 8'h10 ;
			data[77526] <= 8'h10 ;
			data[77527] <= 8'h10 ;
			data[77528] <= 8'h10 ;
			data[77529] <= 8'h10 ;
			data[77530] <= 8'h10 ;
			data[77531] <= 8'h10 ;
			data[77532] <= 8'h10 ;
			data[77533] <= 8'h10 ;
			data[77534] <= 8'h10 ;
			data[77535] <= 8'h10 ;
			data[77536] <= 8'h10 ;
			data[77537] <= 8'h10 ;
			data[77538] <= 8'h10 ;
			data[77539] <= 8'h10 ;
			data[77540] <= 8'h10 ;
			data[77541] <= 8'h10 ;
			data[77542] <= 8'h10 ;
			data[77543] <= 8'h10 ;
			data[77544] <= 8'h10 ;
			data[77545] <= 8'h10 ;
			data[77546] <= 8'h10 ;
			data[77547] <= 8'h10 ;
			data[77548] <= 8'h10 ;
			data[77549] <= 8'h10 ;
			data[77550] <= 8'h10 ;
			data[77551] <= 8'h10 ;
			data[77552] <= 8'h10 ;
			data[77553] <= 8'h10 ;
			data[77554] <= 8'h10 ;
			data[77555] <= 8'h10 ;
			data[77556] <= 8'h10 ;
			data[77557] <= 8'h10 ;
			data[77558] <= 8'h10 ;
			data[77559] <= 8'h10 ;
			data[77560] <= 8'h10 ;
			data[77561] <= 8'h10 ;
			data[77562] <= 8'h10 ;
			data[77563] <= 8'h10 ;
			data[77564] <= 8'h10 ;
			data[77565] <= 8'h10 ;
			data[77566] <= 8'h10 ;
			data[77567] <= 8'h10 ;
			data[77568] <= 8'h10 ;
			data[77569] <= 8'h10 ;
			data[77570] <= 8'h10 ;
			data[77571] <= 8'h10 ;
			data[77572] <= 8'h10 ;
			data[77573] <= 8'h10 ;
			data[77574] <= 8'h10 ;
			data[77575] <= 8'h10 ;
			data[77576] <= 8'h10 ;
			data[77577] <= 8'h10 ;
			data[77578] <= 8'h10 ;
			data[77579] <= 8'h10 ;
			data[77580] <= 8'h10 ;
			data[77581] <= 8'h10 ;
			data[77582] <= 8'h10 ;
			data[77583] <= 8'h10 ;
			data[77584] <= 8'h10 ;
			data[77585] <= 8'h10 ;
			data[77586] <= 8'h10 ;
			data[77587] <= 8'h10 ;
			data[77588] <= 8'h10 ;
			data[77589] <= 8'h10 ;
			data[77590] <= 8'h10 ;
			data[77591] <= 8'h10 ;
			data[77592] <= 8'h10 ;
			data[77593] <= 8'h10 ;
			data[77594] <= 8'h10 ;
			data[77595] <= 8'h10 ;
			data[77596] <= 8'h10 ;
			data[77597] <= 8'h10 ;
			data[77598] <= 8'h10 ;
			data[77599] <= 8'h10 ;
			data[77600] <= 8'h10 ;
			data[77601] <= 8'h10 ;
			data[77602] <= 8'h10 ;
			data[77603] <= 8'h10 ;
			data[77604] <= 8'h10 ;
			data[77605] <= 8'h10 ;
			data[77606] <= 8'h10 ;
			data[77607] <= 8'h10 ;
			data[77608] <= 8'h10 ;
			data[77609] <= 8'h10 ;
			data[77610] <= 8'h10 ;
			data[77611] <= 8'h10 ;
			data[77612] <= 8'h10 ;
			data[77613] <= 8'h10 ;
			data[77614] <= 8'h10 ;
			data[77615] <= 8'h10 ;
			data[77616] <= 8'h10 ;
			data[77617] <= 8'h10 ;
			data[77618] <= 8'h10 ;
			data[77619] <= 8'h10 ;
			data[77620] <= 8'h10 ;
			data[77621] <= 8'h10 ;
			data[77622] <= 8'h10 ;
			data[77623] <= 8'h10 ;
			data[77624] <= 8'h10 ;
			data[77625] <= 8'h10 ;
			data[77626] <= 8'h10 ;
			data[77627] <= 8'h10 ;
			data[77628] <= 8'h10 ;
			data[77629] <= 8'h10 ;
			data[77630] <= 8'h10 ;
			data[77631] <= 8'h10 ;
			data[77632] <= 8'h10 ;
			data[77633] <= 8'h10 ;
			data[77634] <= 8'h10 ;
			data[77635] <= 8'h10 ;
			data[77636] <= 8'h10 ;
			data[77637] <= 8'h10 ;
			data[77638] <= 8'h10 ;
			data[77639] <= 8'h10 ;
			data[77640] <= 8'h10 ;
			data[77641] <= 8'h10 ;
			data[77642] <= 8'h10 ;
			data[77643] <= 8'h10 ;
			data[77644] <= 8'h10 ;
			data[77645] <= 8'h10 ;
			data[77646] <= 8'h10 ;
			data[77647] <= 8'h10 ;
			data[77648] <= 8'h10 ;
			data[77649] <= 8'h10 ;
			data[77650] <= 8'h10 ;
			data[77651] <= 8'h10 ;
			data[77652] <= 8'h10 ;
			data[77653] <= 8'h10 ;
			data[77654] <= 8'h10 ;
			data[77655] <= 8'h10 ;
			data[77656] <= 8'h10 ;
			data[77657] <= 8'h10 ;
			data[77658] <= 8'h10 ;
			data[77659] <= 8'h10 ;
			data[77660] <= 8'h10 ;
			data[77661] <= 8'h10 ;
			data[77662] <= 8'h10 ;
			data[77663] <= 8'h10 ;
			data[77664] <= 8'h10 ;
			data[77665] <= 8'h10 ;
			data[77666] <= 8'h10 ;
			data[77667] <= 8'h10 ;
			data[77668] <= 8'h10 ;
			data[77669] <= 8'h10 ;
			data[77670] <= 8'h10 ;
			data[77671] <= 8'h10 ;
			data[77672] <= 8'h10 ;
			data[77673] <= 8'h10 ;
			data[77674] <= 8'h10 ;
			data[77675] <= 8'h10 ;
			data[77676] <= 8'h10 ;
			data[77677] <= 8'h10 ;
			data[77678] <= 8'h10 ;
			data[77679] <= 8'h10 ;
			data[77680] <= 8'h10 ;
			data[77681] <= 8'h10 ;
			data[77682] <= 8'h10 ;
			data[77683] <= 8'h10 ;
			data[77684] <= 8'h10 ;
			data[77685] <= 8'h10 ;
			data[77686] <= 8'h10 ;
			data[77687] <= 8'h10 ;
			data[77688] <= 8'h10 ;
			data[77689] <= 8'h10 ;
			data[77690] <= 8'h10 ;
			data[77691] <= 8'h10 ;
			data[77692] <= 8'h10 ;
			data[77693] <= 8'h10 ;
			data[77694] <= 8'h10 ;
			data[77695] <= 8'h10 ;
			data[77696] <= 8'h10 ;
			data[77697] <= 8'h10 ;
			data[77698] <= 8'h10 ;
			data[77699] <= 8'h10 ;
			data[77700] <= 8'h10 ;
			data[77701] <= 8'h10 ;
			data[77702] <= 8'h10 ;
			data[77703] <= 8'h10 ;
			data[77704] <= 8'h10 ;
			data[77705] <= 8'h10 ;
			data[77706] <= 8'h10 ;
			data[77707] <= 8'h10 ;
			data[77708] <= 8'h10 ;
			data[77709] <= 8'h10 ;
			data[77710] <= 8'h10 ;
			data[77711] <= 8'h10 ;
			data[77712] <= 8'h10 ;
			data[77713] <= 8'h10 ;
			data[77714] <= 8'h10 ;
			data[77715] <= 8'h10 ;
			data[77716] <= 8'h10 ;
			data[77717] <= 8'h10 ;
			data[77718] <= 8'h10 ;
			data[77719] <= 8'h10 ;
			data[77720] <= 8'h10 ;
			data[77721] <= 8'h10 ;
			data[77722] <= 8'h10 ;
			data[77723] <= 8'h10 ;
			data[77724] <= 8'h10 ;
			data[77725] <= 8'h10 ;
			data[77726] <= 8'h10 ;
			data[77727] <= 8'h10 ;
			data[77728] <= 8'h10 ;
			data[77729] <= 8'h10 ;
			data[77730] <= 8'h10 ;
			data[77731] <= 8'h10 ;
			data[77732] <= 8'h10 ;
			data[77733] <= 8'h10 ;
			data[77734] <= 8'h10 ;
			data[77735] <= 8'h10 ;
			data[77736] <= 8'h10 ;
			data[77737] <= 8'h10 ;
			data[77738] <= 8'h10 ;
			data[77739] <= 8'h10 ;
			data[77740] <= 8'h10 ;
			data[77741] <= 8'h10 ;
			data[77742] <= 8'h10 ;
			data[77743] <= 8'h10 ;
			data[77744] <= 8'h10 ;
			data[77745] <= 8'h10 ;
			data[77746] <= 8'h10 ;
			data[77747] <= 8'h10 ;
			data[77748] <= 8'h10 ;
			data[77749] <= 8'h10 ;
			data[77750] <= 8'h10 ;
			data[77751] <= 8'h10 ;
			data[77752] <= 8'h10 ;
			data[77753] <= 8'h10 ;
			data[77754] <= 8'h10 ;
			data[77755] <= 8'h10 ;
			data[77756] <= 8'h10 ;
			data[77757] <= 8'h10 ;
			data[77758] <= 8'h10 ;
			data[77759] <= 8'h10 ;
			data[77760] <= 8'h10 ;
			data[77761] <= 8'h10 ;
			data[77762] <= 8'h10 ;
			data[77763] <= 8'h10 ;
			data[77764] <= 8'h10 ;
			data[77765] <= 8'h10 ;
			data[77766] <= 8'h10 ;
			data[77767] <= 8'h10 ;
			data[77768] <= 8'h10 ;
			data[77769] <= 8'h10 ;
			data[77770] <= 8'h10 ;
			data[77771] <= 8'h10 ;
			data[77772] <= 8'h10 ;
			data[77773] <= 8'h10 ;
			data[77774] <= 8'h10 ;
			data[77775] <= 8'h10 ;
			data[77776] <= 8'h10 ;
			data[77777] <= 8'h10 ;
			data[77778] <= 8'h10 ;
			data[77779] <= 8'h10 ;
			data[77780] <= 8'h10 ;
			data[77781] <= 8'h10 ;
			data[77782] <= 8'h10 ;
			data[77783] <= 8'h10 ;
			data[77784] <= 8'h10 ;
			data[77785] <= 8'h10 ;
			data[77786] <= 8'h10 ;
			data[77787] <= 8'h10 ;
			data[77788] <= 8'h10 ;
			data[77789] <= 8'h10 ;
			data[77790] <= 8'h10 ;
			data[77791] <= 8'h10 ;
			data[77792] <= 8'h10 ;
			data[77793] <= 8'h10 ;
			data[77794] <= 8'h10 ;
			data[77795] <= 8'h10 ;
			data[77796] <= 8'h10 ;
			data[77797] <= 8'h10 ;
			data[77798] <= 8'h10 ;
			data[77799] <= 8'h10 ;
			data[77800] <= 8'h10 ;
			data[77801] <= 8'h10 ;
			data[77802] <= 8'h10 ;
			data[77803] <= 8'h10 ;
			data[77804] <= 8'h10 ;
			data[77805] <= 8'h10 ;
			data[77806] <= 8'h10 ;
			data[77807] <= 8'h10 ;
			data[77808] <= 8'h10 ;
			data[77809] <= 8'h10 ;
			data[77810] <= 8'h10 ;
			data[77811] <= 8'h10 ;
			data[77812] <= 8'h10 ;
			data[77813] <= 8'h10 ;
			data[77814] <= 8'h10 ;
			data[77815] <= 8'h10 ;
			data[77816] <= 8'h10 ;
			data[77817] <= 8'h10 ;
			data[77818] <= 8'h10 ;
			data[77819] <= 8'h10 ;
			data[77820] <= 8'h10 ;
			data[77821] <= 8'h10 ;
			data[77822] <= 8'h10 ;
			data[77823] <= 8'h10 ;
			data[77824] <= 8'h10 ;
			data[77825] <= 8'h10 ;
			data[77826] <= 8'h10 ;
			data[77827] <= 8'h10 ;
			data[77828] <= 8'h10 ;
			data[77829] <= 8'h10 ;
			data[77830] <= 8'h10 ;
			data[77831] <= 8'h10 ;
			data[77832] <= 8'h10 ;
			data[77833] <= 8'h10 ;
			data[77834] <= 8'h10 ;
			data[77835] <= 8'h10 ;
			data[77836] <= 8'h10 ;
			data[77837] <= 8'h10 ;
			data[77838] <= 8'h10 ;
			data[77839] <= 8'h10 ;
			data[77840] <= 8'h10 ;
			data[77841] <= 8'h10 ;
			data[77842] <= 8'h10 ;
			data[77843] <= 8'h10 ;
			data[77844] <= 8'h10 ;
			data[77845] <= 8'h10 ;
			data[77846] <= 8'h10 ;
			data[77847] <= 8'h10 ;
			data[77848] <= 8'h10 ;
			data[77849] <= 8'h10 ;
			data[77850] <= 8'h10 ;
			data[77851] <= 8'h10 ;
			data[77852] <= 8'h10 ;
			data[77853] <= 8'h10 ;
			data[77854] <= 8'h10 ;
			data[77855] <= 8'h10 ;
			data[77856] <= 8'h10 ;
			data[77857] <= 8'h10 ;
			data[77858] <= 8'h10 ;
			data[77859] <= 8'h10 ;
			data[77860] <= 8'h10 ;
			data[77861] <= 8'h10 ;
			data[77862] <= 8'h10 ;
			data[77863] <= 8'h10 ;
			data[77864] <= 8'h10 ;
			data[77865] <= 8'h10 ;
			data[77866] <= 8'h10 ;
			data[77867] <= 8'h10 ;
			data[77868] <= 8'h10 ;
			data[77869] <= 8'h10 ;
			data[77870] <= 8'h10 ;
			data[77871] <= 8'h10 ;
			data[77872] <= 8'h10 ;
			data[77873] <= 8'h10 ;
			data[77874] <= 8'h10 ;
			data[77875] <= 8'h10 ;
			data[77876] <= 8'h10 ;
			data[77877] <= 8'h10 ;
			data[77878] <= 8'h10 ;
			data[77879] <= 8'h10 ;
			data[77880] <= 8'h10 ;
			data[77881] <= 8'h10 ;
			data[77882] <= 8'h10 ;
			data[77883] <= 8'h10 ;
			data[77884] <= 8'h10 ;
			data[77885] <= 8'h10 ;
			data[77886] <= 8'h10 ;
			data[77887] <= 8'h10 ;
			data[77888] <= 8'h10 ;
			data[77889] <= 8'h10 ;
			data[77890] <= 8'h10 ;
			data[77891] <= 8'h10 ;
			data[77892] <= 8'h10 ;
			data[77893] <= 8'h10 ;
			data[77894] <= 8'h10 ;
			data[77895] <= 8'h10 ;
			data[77896] <= 8'h10 ;
			data[77897] <= 8'h10 ;
			data[77898] <= 8'h10 ;
			data[77899] <= 8'h10 ;
			data[77900] <= 8'h10 ;
			data[77901] <= 8'h10 ;
			data[77902] <= 8'h10 ;
			data[77903] <= 8'h10 ;
			data[77904] <= 8'h10 ;
			data[77905] <= 8'h10 ;
			data[77906] <= 8'h10 ;
			data[77907] <= 8'h10 ;
			data[77908] <= 8'h10 ;
			data[77909] <= 8'h10 ;
			data[77910] <= 8'h10 ;
			data[77911] <= 8'h10 ;
			data[77912] <= 8'h10 ;
			data[77913] <= 8'h10 ;
			data[77914] <= 8'h10 ;
			data[77915] <= 8'h10 ;
			data[77916] <= 8'h10 ;
			data[77917] <= 8'h10 ;
			data[77918] <= 8'h10 ;
			data[77919] <= 8'h10 ;
			data[77920] <= 8'h10 ;
			data[77921] <= 8'h10 ;
			data[77922] <= 8'h10 ;
			data[77923] <= 8'h10 ;
			data[77924] <= 8'h10 ;
			data[77925] <= 8'h10 ;
			data[77926] <= 8'h10 ;
			data[77927] <= 8'h10 ;
			data[77928] <= 8'h10 ;
			data[77929] <= 8'h10 ;
			data[77930] <= 8'h10 ;
			data[77931] <= 8'h10 ;
			data[77932] <= 8'h10 ;
			data[77933] <= 8'h10 ;
			data[77934] <= 8'h10 ;
			data[77935] <= 8'h10 ;
			data[77936] <= 8'h10 ;
			data[77937] <= 8'h10 ;
			data[77938] <= 8'h10 ;
			data[77939] <= 8'h10 ;
			data[77940] <= 8'h10 ;
			data[77941] <= 8'h10 ;
			data[77942] <= 8'h10 ;
			data[77943] <= 8'h10 ;
			data[77944] <= 8'h10 ;
			data[77945] <= 8'h10 ;
			data[77946] <= 8'h10 ;
			data[77947] <= 8'h10 ;
			data[77948] <= 8'h10 ;
			data[77949] <= 8'h10 ;
			data[77950] <= 8'h10 ;
			data[77951] <= 8'h10 ;
			data[77952] <= 8'h10 ;
			data[77953] <= 8'h10 ;
			data[77954] <= 8'h10 ;
			data[77955] <= 8'h10 ;
			data[77956] <= 8'h10 ;
			data[77957] <= 8'h10 ;
			data[77958] <= 8'h10 ;
			data[77959] <= 8'h10 ;
			data[77960] <= 8'h10 ;
			data[77961] <= 8'h10 ;
			data[77962] <= 8'h10 ;
			data[77963] <= 8'h10 ;
			data[77964] <= 8'h10 ;
			data[77965] <= 8'h10 ;
			data[77966] <= 8'h10 ;
			data[77967] <= 8'h10 ;
			data[77968] <= 8'h10 ;
			data[77969] <= 8'h10 ;
			data[77970] <= 8'h10 ;
			data[77971] <= 8'h10 ;
			data[77972] <= 8'h10 ;
			data[77973] <= 8'h10 ;
			data[77974] <= 8'h10 ;
			data[77975] <= 8'h10 ;
			data[77976] <= 8'h10 ;
			data[77977] <= 8'h10 ;
			data[77978] <= 8'h10 ;
			data[77979] <= 8'h10 ;
			data[77980] <= 8'h10 ;
			data[77981] <= 8'h10 ;
			data[77982] <= 8'h10 ;
			data[77983] <= 8'h10 ;
			data[77984] <= 8'h10 ;
			data[77985] <= 8'h10 ;
			data[77986] <= 8'h10 ;
			data[77987] <= 8'h10 ;
			data[77988] <= 8'h10 ;
			data[77989] <= 8'h10 ;
			data[77990] <= 8'h10 ;
			data[77991] <= 8'h10 ;
			data[77992] <= 8'h10 ;
			data[77993] <= 8'h10 ;
			data[77994] <= 8'h10 ;
			data[77995] <= 8'h10 ;
			data[77996] <= 8'h10 ;
			data[77997] <= 8'h10 ;
			data[77998] <= 8'h10 ;
			data[77999] <= 8'h10 ;
			data[78000] <= 8'h10 ;
			data[78001] <= 8'h10 ;
			data[78002] <= 8'h10 ;
			data[78003] <= 8'h10 ;
			data[78004] <= 8'h10 ;
			data[78005] <= 8'h10 ;
			data[78006] <= 8'h10 ;
			data[78007] <= 8'h10 ;
			data[78008] <= 8'h10 ;
			data[78009] <= 8'h10 ;
			data[78010] <= 8'h10 ;
			data[78011] <= 8'h10 ;
			data[78012] <= 8'h10 ;
			data[78013] <= 8'h10 ;
			data[78014] <= 8'h10 ;
			data[78015] <= 8'h10 ;
			data[78016] <= 8'h10 ;
			data[78017] <= 8'h10 ;
			data[78018] <= 8'h10 ;
			data[78019] <= 8'h10 ;
			data[78020] <= 8'h10 ;
			data[78021] <= 8'h10 ;
			data[78022] <= 8'h10 ;
			data[78023] <= 8'h10 ;
			data[78024] <= 8'h10 ;
			data[78025] <= 8'h10 ;
			data[78026] <= 8'h10 ;
			data[78027] <= 8'h10 ;
			data[78028] <= 8'h10 ;
			data[78029] <= 8'h10 ;
			data[78030] <= 8'h10 ;
			data[78031] <= 8'h10 ;
			data[78032] <= 8'h10 ;
			data[78033] <= 8'h10 ;
			data[78034] <= 8'h10 ;
			data[78035] <= 8'h10 ;
			data[78036] <= 8'h10 ;
			data[78037] <= 8'h10 ;
			data[78038] <= 8'h10 ;
			data[78039] <= 8'h10 ;
			data[78040] <= 8'h10 ;
			data[78041] <= 8'h10 ;
			data[78042] <= 8'h10 ;
			data[78043] <= 8'h10 ;
			data[78044] <= 8'h10 ;
			data[78045] <= 8'h10 ;
			data[78046] <= 8'h10 ;
			data[78047] <= 8'h10 ;
			data[78048] <= 8'h10 ;
			data[78049] <= 8'h10 ;
			data[78050] <= 8'h10 ;
			data[78051] <= 8'h10 ;
			data[78052] <= 8'h10 ;
			data[78053] <= 8'h10 ;
			data[78054] <= 8'h10 ;
			data[78055] <= 8'h10 ;
			data[78056] <= 8'h10 ;
			data[78057] <= 8'h10 ;
			data[78058] <= 8'h10 ;
			data[78059] <= 8'h10 ;
			data[78060] <= 8'h10 ;
			data[78061] <= 8'h10 ;
			data[78062] <= 8'h10 ;
			data[78063] <= 8'h10 ;
			data[78064] <= 8'h10 ;
			data[78065] <= 8'h10 ;
			data[78066] <= 8'h10 ;
			data[78067] <= 8'h10 ;
			data[78068] <= 8'h10 ;
			data[78069] <= 8'h10 ;
			data[78070] <= 8'h10 ;
			data[78071] <= 8'h10 ;
			data[78072] <= 8'h10 ;
			data[78073] <= 8'h10 ;
			data[78074] <= 8'h10 ;
			data[78075] <= 8'h10 ;
			data[78076] <= 8'h10 ;
			data[78077] <= 8'h10 ;
			data[78078] <= 8'h10 ;
			data[78079] <= 8'h10 ;
			data[78080] <= 8'h10 ;
			data[78081] <= 8'h10 ;
			data[78082] <= 8'h10 ;
			data[78083] <= 8'h10 ;
			data[78084] <= 8'h10 ;
			data[78085] <= 8'h10 ;
			data[78086] <= 8'h10 ;
			data[78087] <= 8'h10 ;
			data[78088] <= 8'h10 ;
			data[78089] <= 8'h10 ;
			data[78090] <= 8'h10 ;
			data[78091] <= 8'h10 ;
			data[78092] <= 8'h10 ;
			data[78093] <= 8'h10 ;
			data[78094] <= 8'h10 ;
			data[78095] <= 8'h10 ;
			data[78096] <= 8'h10 ;
			data[78097] <= 8'h10 ;
			data[78098] <= 8'h10 ;
			data[78099] <= 8'h10 ;
			data[78100] <= 8'h10 ;
			data[78101] <= 8'h10 ;
			data[78102] <= 8'h10 ;
			data[78103] <= 8'h10 ;
			data[78104] <= 8'h10 ;
			data[78105] <= 8'h10 ;
			data[78106] <= 8'h10 ;
			data[78107] <= 8'h10 ;
			data[78108] <= 8'h10 ;
			data[78109] <= 8'h10 ;
			data[78110] <= 8'h10 ;
			data[78111] <= 8'h10 ;
			data[78112] <= 8'h10 ;
			data[78113] <= 8'h10 ;
			data[78114] <= 8'h10 ;
			data[78115] <= 8'h10 ;
			data[78116] <= 8'h10 ;
			data[78117] <= 8'h10 ;
			data[78118] <= 8'h10 ;
			data[78119] <= 8'h10 ;
			data[78120] <= 8'h10 ;
			data[78121] <= 8'h10 ;
			data[78122] <= 8'h10 ;
			data[78123] <= 8'h10 ;
			data[78124] <= 8'h10 ;
			data[78125] <= 8'h10 ;
			data[78126] <= 8'h10 ;
			data[78127] <= 8'h10 ;
			data[78128] <= 8'h10 ;
			data[78129] <= 8'h10 ;
			data[78130] <= 8'h10 ;
			data[78131] <= 8'h10 ;
			data[78132] <= 8'h10 ;
			data[78133] <= 8'h10 ;
			data[78134] <= 8'h10 ;
			data[78135] <= 8'h10 ;
			data[78136] <= 8'h10 ;
			data[78137] <= 8'h10 ;
			data[78138] <= 8'h10 ;
			data[78139] <= 8'h10 ;
			data[78140] <= 8'h10 ;
			data[78141] <= 8'h10 ;
			data[78142] <= 8'h10 ;
			data[78143] <= 8'h10 ;
			data[78144] <= 8'h10 ;
			data[78145] <= 8'h10 ;
			data[78146] <= 8'h10 ;
			data[78147] <= 8'h10 ;
			data[78148] <= 8'h10 ;
			data[78149] <= 8'h10 ;
			data[78150] <= 8'h10 ;
			data[78151] <= 8'h10 ;
			data[78152] <= 8'h10 ;
			data[78153] <= 8'h10 ;
			data[78154] <= 8'h10 ;
			data[78155] <= 8'h10 ;
			data[78156] <= 8'h10 ;
			data[78157] <= 8'h10 ;
			data[78158] <= 8'h10 ;
			data[78159] <= 8'h10 ;
			data[78160] <= 8'h10 ;
			data[78161] <= 8'h10 ;
			data[78162] <= 8'h10 ;
			data[78163] <= 8'h10 ;
			data[78164] <= 8'h10 ;
			data[78165] <= 8'h10 ;
			data[78166] <= 8'h10 ;
			data[78167] <= 8'h10 ;
			data[78168] <= 8'h10 ;
			data[78169] <= 8'h10 ;
			data[78170] <= 8'h10 ;
			data[78171] <= 8'h10 ;
			data[78172] <= 8'h10 ;
			data[78173] <= 8'h10 ;
			data[78174] <= 8'h10 ;
			data[78175] <= 8'h10 ;
			data[78176] <= 8'h10 ;
			data[78177] <= 8'h10 ;
			data[78178] <= 8'h10 ;
			data[78179] <= 8'h10 ;
			data[78180] <= 8'h10 ;
			data[78181] <= 8'h10 ;
			data[78182] <= 8'h10 ;
			data[78183] <= 8'h10 ;
			data[78184] <= 8'h10 ;
			data[78185] <= 8'h10 ;
			data[78186] <= 8'h10 ;
			data[78187] <= 8'h10 ;
			data[78188] <= 8'h10 ;
			data[78189] <= 8'h10 ;
			data[78190] <= 8'h10 ;
			data[78191] <= 8'h10 ;
			data[78192] <= 8'h10 ;
			data[78193] <= 8'h10 ;
			data[78194] <= 8'h10 ;
			data[78195] <= 8'h10 ;
			data[78196] <= 8'h10 ;
			data[78197] <= 8'h10 ;
			data[78198] <= 8'h10 ;
			data[78199] <= 8'h10 ;
			data[78200] <= 8'h10 ;
			data[78201] <= 8'h10 ;
			data[78202] <= 8'h10 ;
			data[78203] <= 8'h10 ;
			data[78204] <= 8'h10 ;
			data[78205] <= 8'h10 ;
			data[78206] <= 8'h10 ;
			data[78207] <= 8'h10 ;
			data[78208] <= 8'h10 ;
			data[78209] <= 8'h10 ;
			data[78210] <= 8'h10 ;
			data[78211] <= 8'h10 ;
			data[78212] <= 8'h10 ;
			data[78213] <= 8'h10 ;
			data[78214] <= 8'h10 ;
			data[78215] <= 8'h10 ;
			data[78216] <= 8'h10 ;
			data[78217] <= 8'h10 ;
			data[78218] <= 8'h10 ;
			data[78219] <= 8'h10 ;
			data[78220] <= 8'h10 ;
			data[78221] <= 8'h10 ;
			data[78222] <= 8'h10 ;
			data[78223] <= 8'h10 ;
			data[78224] <= 8'h10 ;
			data[78225] <= 8'h10 ;
			data[78226] <= 8'h10 ;
			data[78227] <= 8'h10 ;
			data[78228] <= 8'h10 ;
			data[78229] <= 8'h10 ;
			data[78230] <= 8'h10 ;
			data[78231] <= 8'h10 ;
			data[78232] <= 8'h10 ;
			data[78233] <= 8'h10 ;
			data[78234] <= 8'h10 ;
			data[78235] <= 8'h10 ;
			data[78236] <= 8'h10 ;
			data[78237] <= 8'h10 ;
			data[78238] <= 8'h10 ;
			data[78239] <= 8'h10 ;
			data[78240] <= 8'h10 ;
			data[78241] <= 8'h10 ;
			data[78242] <= 8'h10 ;
			data[78243] <= 8'h10 ;
			data[78244] <= 8'h10 ;
			data[78245] <= 8'h10 ;
			data[78246] <= 8'h10 ;
			data[78247] <= 8'h10 ;
			data[78248] <= 8'h10 ;
			data[78249] <= 8'h10 ;
			data[78250] <= 8'h10 ;
			data[78251] <= 8'h10 ;
			data[78252] <= 8'h10 ;
			data[78253] <= 8'h10 ;
			data[78254] <= 8'h10 ;
			data[78255] <= 8'h10 ;
			data[78256] <= 8'h10 ;
			data[78257] <= 8'h10 ;
			data[78258] <= 8'h10 ;
			data[78259] <= 8'h10 ;
			data[78260] <= 8'h10 ;
			data[78261] <= 8'h10 ;
			data[78262] <= 8'h10 ;
			data[78263] <= 8'h10 ;
			data[78264] <= 8'h10 ;
			data[78265] <= 8'h10 ;
			data[78266] <= 8'h10 ;
			data[78267] <= 8'h10 ;
			data[78268] <= 8'h10 ;
			data[78269] <= 8'h10 ;
			data[78270] <= 8'h10 ;
			data[78271] <= 8'h10 ;
			data[78272] <= 8'h10 ;
			data[78273] <= 8'h10 ;
			data[78274] <= 8'h10 ;
			data[78275] <= 8'h10 ;
			data[78276] <= 8'h10 ;
			data[78277] <= 8'h10 ;
			data[78278] <= 8'h10 ;
			data[78279] <= 8'h10 ;
			data[78280] <= 8'h10 ;
			data[78281] <= 8'h10 ;
			data[78282] <= 8'h10 ;
			data[78283] <= 8'h10 ;
			data[78284] <= 8'h10 ;
			data[78285] <= 8'h10 ;
			data[78286] <= 8'h10 ;
			data[78287] <= 8'h10 ;
			data[78288] <= 8'h10 ;
			data[78289] <= 8'h10 ;
			data[78290] <= 8'h10 ;
			data[78291] <= 8'h10 ;
			data[78292] <= 8'h10 ;
			data[78293] <= 8'h10 ;
			data[78294] <= 8'h10 ;
			data[78295] <= 8'h10 ;
			data[78296] <= 8'h10 ;
			data[78297] <= 8'h10 ;
			data[78298] <= 8'h10 ;
			data[78299] <= 8'h10 ;
			data[78300] <= 8'h10 ;
			data[78301] <= 8'h10 ;
			data[78302] <= 8'h10 ;
			data[78303] <= 8'h10 ;
			data[78304] <= 8'h10 ;
			data[78305] <= 8'h10 ;
			data[78306] <= 8'h10 ;
			data[78307] <= 8'h10 ;
			data[78308] <= 8'h10 ;
			data[78309] <= 8'h10 ;
			data[78310] <= 8'h10 ;
			data[78311] <= 8'h10 ;
			data[78312] <= 8'h10 ;
			data[78313] <= 8'h10 ;
			data[78314] <= 8'h10 ;
			data[78315] <= 8'h10 ;
			data[78316] <= 8'h10 ;
			data[78317] <= 8'h10 ;
			data[78318] <= 8'h10 ;
			data[78319] <= 8'h10 ;
			data[78320] <= 8'h10 ;
			data[78321] <= 8'h10 ;
			data[78322] <= 8'h10 ;
			data[78323] <= 8'h10 ;
			data[78324] <= 8'h10 ;
			data[78325] <= 8'h10 ;
			data[78326] <= 8'h10 ;
			data[78327] <= 8'h10 ;
			data[78328] <= 8'h10 ;
			data[78329] <= 8'h10 ;
			data[78330] <= 8'h10 ;
			data[78331] <= 8'h10 ;
			data[78332] <= 8'h10 ;
			data[78333] <= 8'h10 ;
			data[78334] <= 8'h10 ;
			data[78335] <= 8'h10 ;
			data[78336] <= 8'h10 ;
			data[78337] <= 8'h10 ;
			data[78338] <= 8'h10 ;
			data[78339] <= 8'h10 ;
			data[78340] <= 8'h10 ;
			data[78341] <= 8'h10 ;
			data[78342] <= 8'h10 ;
			data[78343] <= 8'h10 ;
			data[78344] <= 8'h10 ;
			data[78345] <= 8'h10 ;
			data[78346] <= 8'h10 ;
			data[78347] <= 8'h10 ;
			data[78348] <= 8'h10 ;
			data[78349] <= 8'h10 ;
			data[78350] <= 8'h10 ;
			data[78351] <= 8'h10 ;
			data[78352] <= 8'h10 ;
			data[78353] <= 8'h10 ;
			data[78354] <= 8'h10 ;
			data[78355] <= 8'h10 ;
			data[78356] <= 8'h10 ;
			data[78357] <= 8'h10 ;
			data[78358] <= 8'h10 ;
			data[78359] <= 8'h10 ;
			data[78360] <= 8'h10 ;
			data[78361] <= 8'h10 ;
			data[78362] <= 8'h10 ;
			data[78363] <= 8'h10 ;
			data[78364] <= 8'h10 ;
			data[78365] <= 8'h10 ;
			data[78366] <= 8'h10 ;
			data[78367] <= 8'h10 ;
			data[78368] <= 8'h10 ;
			data[78369] <= 8'h10 ;
			data[78370] <= 8'h10 ;
			data[78371] <= 8'h10 ;
			data[78372] <= 8'h10 ;
			data[78373] <= 8'h10 ;
			data[78374] <= 8'h10 ;
			data[78375] <= 8'h10 ;
			data[78376] <= 8'h10 ;
			data[78377] <= 8'h10 ;
			data[78378] <= 8'h10 ;
			data[78379] <= 8'h10 ;
			data[78380] <= 8'h10 ;
			data[78381] <= 8'h10 ;
			data[78382] <= 8'h10 ;
			data[78383] <= 8'h10 ;
			data[78384] <= 8'h10 ;
			data[78385] <= 8'h10 ;
			data[78386] <= 8'h10 ;
			data[78387] <= 8'h10 ;
			data[78388] <= 8'h10 ;
			data[78389] <= 8'h10 ;
			data[78390] <= 8'h10 ;
			data[78391] <= 8'h10 ;
			data[78392] <= 8'h10 ;
			data[78393] <= 8'h10 ;
			data[78394] <= 8'h10 ;
			data[78395] <= 8'h10 ;
			data[78396] <= 8'h10 ;
			data[78397] <= 8'h10 ;
			data[78398] <= 8'h10 ;
			data[78399] <= 8'h10 ;
			data[78400] <= 8'h10 ;
			data[78401] <= 8'h10 ;
			data[78402] <= 8'h10 ;
			data[78403] <= 8'h10 ;
			data[78404] <= 8'h10 ;
			data[78405] <= 8'h10 ;
			data[78406] <= 8'h10 ;
			data[78407] <= 8'h10 ;
			data[78408] <= 8'h10 ;
			data[78409] <= 8'h10 ;
			data[78410] <= 8'h10 ;
			data[78411] <= 8'h10 ;
			data[78412] <= 8'h10 ;
			data[78413] <= 8'h10 ;
			data[78414] <= 8'h10 ;
			data[78415] <= 8'h10 ;
			data[78416] <= 8'h10 ;
			data[78417] <= 8'h10 ;
			data[78418] <= 8'h10 ;
			data[78419] <= 8'h10 ;
			data[78420] <= 8'h10 ;
			data[78421] <= 8'h10 ;
			data[78422] <= 8'h10 ;
			data[78423] <= 8'h10 ;
			data[78424] <= 8'h10 ;
			data[78425] <= 8'h10 ;
			data[78426] <= 8'h10 ;
			data[78427] <= 8'h10 ;
			data[78428] <= 8'h10 ;
			data[78429] <= 8'h10 ;
			data[78430] <= 8'h10 ;
			data[78431] <= 8'h10 ;
			data[78432] <= 8'h10 ;
			data[78433] <= 8'h10 ;
			data[78434] <= 8'h10 ;
			data[78435] <= 8'h10 ;
			data[78436] <= 8'h10 ;
			data[78437] <= 8'h10 ;
			data[78438] <= 8'h10 ;
			data[78439] <= 8'h10 ;
			data[78440] <= 8'h10 ;
			data[78441] <= 8'h10 ;
			data[78442] <= 8'h10 ;
			data[78443] <= 8'h10 ;
			data[78444] <= 8'h10 ;
			data[78445] <= 8'h10 ;
			data[78446] <= 8'h10 ;
			data[78447] <= 8'h10 ;
			data[78448] <= 8'h10 ;
			data[78449] <= 8'h10 ;
			data[78450] <= 8'h10 ;
			data[78451] <= 8'h10 ;
			data[78452] <= 8'h10 ;
			data[78453] <= 8'h10 ;
			data[78454] <= 8'h10 ;
			data[78455] <= 8'h10 ;
			data[78456] <= 8'h10 ;
			data[78457] <= 8'h10 ;
			data[78458] <= 8'h10 ;
			data[78459] <= 8'h10 ;
			data[78460] <= 8'h10 ;
			data[78461] <= 8'h10 ;
			data[78462] <= 8'h10 ;
			data[78463] <= 8'h10 ;
			data[78464] <= 8'h10 ;
			data[78465] <= 8'h10 ;
			data[78466] <= 8'h10 ;
			data[78467] <= 8'h10 ;
			data[78468] <= 8'h10 ;
			data[78469] <= 8'h10 ;
			data[78470] <= 8'h10 ;
			data[78471] <= 8'h10 ;
			data[78472] <= 8'h10 ;
			data[78473] <= 8'h10 ;
			data[78474] <= 8'h10 ;
			data[78475] <= 8'h10 ;
			data[78476] <= 8'h10 ;
			data[78477] <= 8'h10 ;
			data[78478] <= 8'h10 ;
			data[78479] <= 8'h10 ;
			data[78480] <= 8'h10 ;
			data[78481] <= 8'h10 ;
			data[78482] <= 8'h10 ;
			data[78483] <= 8'h10 ;
			data[78484] <= 8'h10 ;
			data[78485] <= 8'h10 ;
			data[78486] <= 8'h10 ;
			data[78487] <= 8'h10 ;
			data[78488] <= 8'h10 ;
			data[78489] <= 8'h10 ;
			data[78490] <= 8'h10 ;
			data[78491] <= 8'h10 ;
			data[78492] <= 8'h10 ;
			data[78493] <= 8'h10 ;
			data[78494] <= 8'h10 ;
			data[78495] <= 8'h10 ;
			data[78496] <= 8'h10 ;
			data[78497] <= 8'h10 ;
			data[78498] <= 8'h10 ;
			data[78499] <= 8'h10 ;
			data[78500] <= 8'h10 ;
			data[78501] <= 8'h10 ;
			data[78502] <= 8'h10 ;
			data[78503] <= 8'h10 ;
			data[78504] <= 8'h10 ;
			data[78505] <= 8'h10 ;
			data[78506] <= 8'h10 ;
			data[78507] <= 8'h10 ;
			data[78508] <= 8'h10 ;
			data[78509] <= 8'h10 ;
			data[78510] <= 8'h10 ;
			data[78511] <= 8'h10 ;
			data[78512] <= 8'h10 ;
			data[78513] <= 8'h10 ;
			data[78514] <= 8'h10 ;
			data[78515] <= 8'h10 ;
			data[78516] <= 8'h10 ;
			data[78517] <= 8'h10 ;
			data[78518] <= 8'h10 ;
			data[78519] <= 8'h10 ;
			data[78520] <= 8'h10 ;
			data[78521] <= 8'h10 ;
			data[78522] <= 8'h10 ;
			data[78523] <= 8'h10 ;
			data[78524] <= 8'h10 ;
			data[78525] <= 8'h10 ;
			data[78526] <= 8'h10 ;
			data[78527] <= 8'h10 ;
			data[78528] <= 8'h10 ;
			data[78529] <= 8'h10 ;
			data[78530] <= 8'h10 ;
			data[78531] <= 8'h10 ;
			data[78532] <= 8'h10 ;
			data[78533] <= 8'h10 ;
			data[78534] <= 8'h10 ;
			data[78535] <= 8'h10 ;
			data[78536] <= 8'h10 ;
			data[78537] <= 8'h10 ;
			data[78538] <= 8'h10 ;
			data[78539] <= 8'h10 ;
			data[78540] <= 8'h10 ;
			data[78541] <= 8'h10 ;
			data[78542] <= 8'h10 ;
			data[78543] <= 8'h10 ;
			data[78544] <= 8'h10 ;
			data[78545] <= 8'h10 ;
			data[78546] <= 8'h10 ;
			data[78547] <= 8'h10 ;
			data[78548] <= 8'h10 ;
			data[78549] <= 8'h10 ;
			data[78550] <= 8'h10 ;
			data[78551] <= 8'h10 ;
			data[78552] <= 8'h10 ;
			data[78553] <= 8'h10 ;
			data[78554] <= 8'h10 ;
			data[78555] <= 8'h10 ;
			data[78556] <= 8'h10 ;
			data[78557] <= 8'h10 ;
			data[78558] <= 8'h10 ;
			data[78559] <= 8'h10 ;
			data[78560] <= 8'h10 ;
			data[78561] <= 8'h10 ;
			data[78562] <= 8'h10 ;
			data[78563] <= 8'h10 ;
			data[78564] <= 8'h10 ;
			data[78565] <= 8'h10 ;
			data[78566] <= 8'h10 ;
			data[78567] <= 8'h10 ;
			data[78568] <= 8'h10 ;
			data[78569] <= 8'h10 ;
			data[78570] <= 8'h10 ;
			data[78571] <= 8'h10 ;
			data[78572] <= 8'h10 ;
			data[78573] <= 8'h10 ;
			data[78574] <= 8'h10 ;
			data[78575] <= 8'h10 ;
			data[78576] <= 8'h10 ;
			data[78577] <= 8'h10 ;
			data[78578] <= 8'h10 ;
			data[78579] <= 8'h10 ;
			data[78580] <= 8'h10 ;
			data[78581] <= 8'h10 ;
			data[78582] <= 8'h10 ;
			data[78583] <= 8'h10 ;
			data[78584] <= 8'h10 ;
			data[78585] <= 8'h10 ;
			data[78586] <= 8'h10 ;
			data[78587] <= 8'h10 ;
			data[78588] <= 8'h10 ;
			data[78589] <= 8'h10 ;
			data[78590] <= 8'h10 ;
			data[78591] <= 8'h10 ;
			data[78592] <= 8'h10 ;
			data[78593] <= 8'h10 ;
			data[78594] <= 8'h10 ;
			data[78595] <= 8'h10 ;
			data[78596] <= 8'h10 ;
			data[78597] <= 8'h10 ;
			data[78598] <= 8'h10 ;
			data[78599] <= 8'h10 ;
			data[78600] <= 8'h10 ;
			data[78601] <= 8'h10 ;
			data[78602] <= 8'h10 ;
			data[78603] <= 8'h10 ;
			data[78604] <= 8'h10 ;
			data[78605] <= 8'h10 ;
			data[78606] <= 8'h10 ;
			data[78607] <= 8'h10 ;
			data[78608] <= 8'h10 ;
			data[78609] <= 8'h10 ;
			data[78610] <= 8'h10 ;
			data[78611] <= 8'h10 ;
			data[78612] <= 8'h10 ;
			data[78613] <= 8'h10 ;
			data[78614] <= 8'h10 ;
			data[78615] <= 8'h10 ;
			data[78616] <= 8'h10 ;
			data[78617] <= 8'h10 ;
			data[78618] <= 8'h10 ;
			data[78619] <= 8'h10 ;
			data[78620] <= 8'h10 ;
			data[78621] <= 8'h10 ;
			data[78622] <= 8'h10 ;
			data[78623] <= 8'h10 ;
			data[78624] <= 8'h10 ;
			data[78625] <= 8'h10 ;
			data[78626] <= 8'h10 ;
			data[78627] <= 8'h10 ;
			data[78628] <= 8'h10 ;
			data[78629] <= 8'h10 ;
			data[78630] <= 8'h10 ;
			data[78631] <= 8'h10 ;
			data[78632] <= 8'h10 ;
			data[78633] <= 8'h10 ;
			data[78634] <= 8'h10 ;
			data[78635] <= 8'h10 ;
			data[78636] <= 8'h10 ;
			data[78637] <= 8'h10 ;
			data[78638] <= 8'h10 ;
			data[78639] <= 8'h10 ;
			data[78640] <= 8'h10 ;
			data[78641] <= 8'h10 ;
			data[78642] <= 8'h10 ;
			data[78643] <= 8'h10 ;
			data[78644] <= 8'h10 ;
			data[78645] <= 8'h10 ;
			data[78646] <= 8'h10 ;
			data[78647] <= 8'h10 ;
			data[78648] <= 8'h10 ;
			data[78649] <= 8'h10 ;
			data[78650] <= 8'h10 ;
			data[78651] <= 8'h10 ;
			data[78652] <= 8'h10 ;
			data[78653] <= 8'h10 ;
			data[78654] <= 8'h10 ;
			data[78655] <= 8'h10 ;
			data[78656] <= 8'h10 ;
			data[78657] <= 8'h10 ;
			data[78658] <= 8'h10 ;
			data[78659] <= 8'h10 ;
			data[78660] <= 8'h10 ;
			data[78661] <= 8'h10 ;
			data[78662] <= 8'h10 ;
			data[78663] <= 8'h10 ;
			data[78664] <= 8'h10 ;
			data[78665] <= 8'h10 ;
			data[78666] <= 8'h10 ;
			data[78667] <= 8'h10 ;
			data[78668] <= 8'h10 ;
			data[78669] <= 8'h10 ;
			data[78670] <= 8'h10 ;
			data[78671] <= 8'h10 ;
			data[78672] <= 8'h10 ;
			data[78673] <= 8'h10 ;
			data[78674] <= 8'h10 ;
			data[78675] <= 8'h10 ;
			data[78676] <= 8'h10 ;
			data[78677] <= 8'h10 ;
			data[78678] <= 8'h10 ;
			data[78679] <= 8'h10 ;
			data[78680] <= 8'h10 ;
			data[78681] <= 8'h10 ;
			data[78682] <= 8'h10 ;
			data[78683] <= 8'h10 ;
			data[78684] <= 8'h10 ;
			data[78685] <= 8'h10 ;
			data[78686] <= 8'h10 ;
			data[78687] <= 8'h10 ;
			data[78688] <= 8'h10 ;
			data[78689] <= 8'h10 ;
			data[78690] <= 8'h10 ;
			data[78691] <= 8'h10 ;
			data[78692] <= 8'h10 ;
			data[78693] <= 8'h10 ;
			data[78694] <= 8'h10 ;
			data[78695] <= 8'h10 ;
			data[78696] <= 8'h10 ;
			data[78697] <= 8'h10 ;
			data[78698] <= 8'h10 ;
			data[78699] <= 8'h10 ;
			data[78700] <= 8'h10 ;
			data[78701] <= 8'h10 ;
			data[78702] <= 8'h10 ;
			data[78703] <= 8'h10 ;
			data[78704] <= 8'h10 ;
			data[78705] <= 8'h10 ;
			data[78706] <= 8'h10 ;
			data[78707] <= 8'h10 ;
			data[78708] <= 8'h10 ;
			data[78709] <= 8'h10 ;
			data[78710] <= 8'h10 ;
			data[78711] <= 8'h10 ;
			data[78712] <= 8'h10 ;
			data[78713] <= 8'h10 ;
			data[78714] <= 8'h10 ;
			data[78715] <= 8'h10 ;
			data[78716] <= 8'h10 ;
			data[78717] <= 8'h10 ;
			data[78718] <= 8'h10 ;
			data[78719] <= 8'h10 ;
			data[78720] <= 8'h10 ;
			data[78721] <= 8'h10 ;
			data[78722] <= 8'h10 ;
			data[78723] <= 8'h10 ;
			data[78724] <= 8'h10 ;
			data[78725] <= 8'h10 ;
			data[78726] <= 8'h10 ;
			data[78727] <= 8'h10 ;
			data[78728] <= 8'h10 ;
			data[78729] <= 8'h10 ;
			data[78730] <= 8'h10 ;
			data[78731] <= 8'h10 ;
			data[78732] <= 8'h10 ;
			data[78733] <= 8'h10 ;
			data[78734] <= 8'h10 ;
			data[78735] <= 8'h10 ;
			data[78736] <= 8'h10 ;
			data[78737] <= 8'h10 ;
			data[78738] <= 8'h10 ;
			data[78739] <= 8'h10 ;
			data[78740] <= 8'h10 ;
			data[78741] <= 8'h10 ;
			data[78742] <= 8'h10 ;
			data[78743] <= 8'h10 ;
			data[78744] <= 8'h10 ;
			data[78745] <= 8'h10 ;
			data[78746] <= 8'h10 ;
			data[78747] <= 8'h10 ;
			data[78748] <= 8'h10 ;
			data[78749] <= 8'h10 ;
			data[78750] <= 8'h10 ;
			data[78751] <= 8'h10 ;
			data[78752] <= 8'h10 ;
			data[78753] <= 8'h10 ;
			data[78754] <= 8'h10 ;
			data[78755] <= 8'h10 ;
			data[78756] <= 8'h10 ;
			data[78757] <= 8'h10 ;
			data[78758] <= 8'h10 ;
			data[78759] <= 8'h10 ;
			data[78760] <= 8'h10 ;
			data[78761] <= 8'h10 ;
			data[78762] <= 8'h10 ;
			data[78763] <= 8'h10 ;
			data[78764] <= 8'h10 ;
			data[78765] <= 8'h10 ;
			data[78766] <= 8'h10 ;
			data[78767] <= 8'h10 ;
			data[78768] <= 8'h10 ;
			data[78769] <= 8'h10 ;
			data[78770] <= 8'h10 ;
			data[78771] <= 8'h10 ;
			data[78772] <= 8'h10 ;
			data[78773] <= 8'h10 ;
			data[78774] <= 8'h10 ;
			data[78775] <= 8'h10 ;
			data[78776] <= 8'h10 ;
			data[78777] <= 8'h10 ;
			data[78778] <= 8'h10 ;
			data[78779] <= 8'h10 ;
			data[78780] <= 8'h10 ;
			data[78781] <= 8'h10 ;
			data[78782] <= 8'h10 ;
			data[78783] <= 8'h10 ;
			data[78784] <= 8'h10 ;
			data[78785] <= 8'h10 ;
			data[78786] <= 8'h10 ;
			data[78787] <= 8'h10 ;
			data[78788] <= 8'h10 ;
			data[78789] <= 8'h10 ;
			data[78790] <= 8'h10 ;
			data[78791] <= 8'h10 ;
			data[78792] <= 8'h10 ;
			data[78793] <= 8'h10 ;
			data[78794] <= 8'h10 ;
			data[78795] <= 8'h10 ;
			data[78796] <= 8'h10 ;
			data[78797] <= 8'h10 ;
			data[78798] <= 8'h10 ;
			data[78799] <= 8'h10 ;
			data[78800] <= 8'h10 ;
			data[78801] <= 8'h10 ;
			data[78802] <= 8'h10 ;
			data[78803] <= 8'h10 ;
			data[78804] <= 8'h10 ;
			data[78805] <= 8'h10 ;
			data[78806] <= 8'h10 ;
			data[78807] <= 8'h10 ;
			data[78808] <= 8'h10 ;
			data[78809] <= 8'h10 ;
			data[78810] <= 8'h10 ;
			data[78811] <= 8'h10 ;
			data[78812] <= 8'h10 ;
			data[78813] <= 8'h10 ;
			data[78814] <= 8'h10 ;
			data[78815] <= 8'h10 ;
			data[78816] <= 8'h10 ;
			data[78817] <= 8'h10 ;
			data[78818] <= 8'h10 ;
			data[78819] <= 8'h10 ;
			data[78820] <= 8'h10 ;
			data[78821] <= 8'h10 ;
			data[78822] <= 8'h10 ;
			data[78823] <= 8'h10 ;
			data[78824] <= 8'h10 ;
			data[78825] <= 8'h10 ;
			data[78826] <= 8'h10 ;
			data[78827] <= 8'h10 ;
			data[78828] <= 8'h10 ;
			data[78829] <= 8'h10 ;
			data[78830] <= 8'h10 ;
			data[78831] <= 8'h10 ;
			data[78832] <= 8'h10 ;
			data[78833] <= 8'h10 ;
			data[78834] <= 8'h10 ;
			data[78835] <= 8'h10 ;
			data[78836] <= 8'h10 ;
			data[78837] <= 8'h10 ;
			data[78838] <= 8'h10 ;
			data[78839] <= 8'h10 ;
			data[78840] <= 8'h10 ;
			data[78841] <= 8'h10 ;
			data[78842] <= 8'h10 ;
			data[78843] <= 8'h10 ;
			data[78844] <= 8'h10 ;
			data[78845] <= 8'h10 ;
			data[78846] <= 8'h10 ;
			data[78847] <= 8'h10 ;
			data[78848] <= 8'h10 ;
			data[78849] <= 8'h10 ;
			data[78850] <= 8'h10 ;
			data[78851] <= 8'h10 ;
			data[78852] <= 8'h10 ;
			data[78853] <= 8'h10 ;
			data[78854] <= 8'h10 ;
			data[78855] <= 8'h10 ;
			data[78856] <= 8'h10 ;
			data[78857] <= 8'h10 ;
			data[78858] <= 8'h10 ;
			data[78859] <= 8'h10 ;
			data[78860] <= 8'h10 ;
			data[78861] <= 8'h10 ;
			data[78862] <= 8'h10 ;
			data[78863] <= 8'h10 ;
			data[78864] <= 8'h10 ;
			data[78865] <= 8'h10 ;
			data[78866] <= 8'h10 ;
			data[78867] <= 8'h10 ;
			data[78868] <= 8'h10 ;
			data[78869] <= 8'h10 ;
			data[78870] <= 8'h10 ;
			data[78871] <= 8'h10 ;
			data[78872] <= 8'h10 ;
			data[78873] <= 8'h10 ;
			data[78874] <= 8'h10 ;
			data[78875] <= 8'h10 ;
			data[78876] <= 8'h10 ;
			data[78877] <= 8'h10 ;
			data[78878] <= 8'h10 ;
			data[78879] <= 8'h10 ;
			data[78880] <= 8'h10 ;
			data[78881] <= 8'h10 ;
			data[78882] <= 8'h10 ;
			data[78883] <= 8'h10 ;
			data[78884] <= 8'h10 ;
			data[78885] <= 8'h10 ;
			data[78886] <= 8'h10 ;
			data[78887] <= 8'h10 ;
			data[78888] <= 8'h10 ;
			data[78889] <= 8'h10 ;
			data[78890] <= 8'h10 ;
			data[78891] <= 8'h10 ;
			data[78892] <= 8'h10 ;
			data[78893] <= 8'h10 ;
			data[78894] <= 8'h10 ;
			data[78895] <= 8'h10 ;
			data[78896] <= 8'h10 ;
			data[78897] <= 8'h10 ;
			data[78898] <= 8'h10 ;
			data[78899] <= 8'h10 ;
			data[78900] <= 8'h10 ;
			data[78901] <= 8'h10 ;
			data[78902] <= 8'h10 ;
			data[78903] <= 8'h10 ;
			data[78904] <= 8'h10 ;
			data[78905] <= 8'h10 ;
			data[78906] <= 8'h10 ;
			data[78907] <= 8'h10 ;
			data[78908] <= 8'h10 ;
			data[78909] <= 8'h10 ;
			data[78910] <= 8'h10 ;
			data[78911] <= 8'h10 ;
			data[78912] <= 8'h10 ;
			data[78913] <= 8'h10 ;
			data[78914] <= 8'h10 ;
			data[78915] <= 8'h10 ;
			data[78916] <= 8'h10 ;
			data[78917] <= 8'h10 ;
			data[78918] <= 8'h10 ;
			data[78919] <= 8'h10 ;
			data[78920] <= 8'h10 ;
			data[78921] <= 8'h10 ;
			data[78922] <= 8'h10 ;
			data[78923] <= 8'h10 ;
			data[78924] <= 8'h10 ;
			data[78925] <= 8'h10 ;
			data[78926] <= 8'h10 ;
			data[78927] <= 8'h10 ;
			data[78928] <= 8'h10 ;
			data[78929] <= 8'h10 ;
			data[78930] <= 8'h10 ;
			data[78931] <= 8'h10 ;
			data[78932] <= 8'h10 ;
			data[78933] <= 8'h10 ;
			data[78934] <= 8'h10 ;
			data[78935] <= 8'h10 ;
			data[78936] <= 8'h10 ;
			data[78937] <= 8'h10 ;
			data[78938] <= 8'h10 ;
			data[78939] <= 8'h10 ;
			data[78940] <= 8'h10 ;
			data[78941] <= 8'h10 ;
			data[78942] <= 8'h10 ;
			data[78943] <= 8'h10 ;
			data[78944] <= 8'h10 ;
			data[78945] <= 8'h10 ;
			data[78946] <= 8'h10 ;
			data[78947] <= 8'h10 ;
			data[78948] <= 8'h10 ;
			data[78949] <= 8'h10 ;
			data[78950] <= 8'h10 ;
			data[78951] <= 8'h10 ;
			data[78952] <= 8'h10 ;
			data[78953] <= 8'h10 ;
			data[78954] <= 8'h10 ;
			data[78955] <= 8'h10 ;
			data[78956] <= 8'h10 ;
			data[78957] <= 8'h10 ;
			data[78958] <= 8'h10 ;
			data[78959] <= 8'h10 ;
			data[78960] <= 8'h10 ;
			data[78961] <= 8'h10 ;
			data[78962] <= 8'h10 ;
			data[78963] <= 8'h10 ;
			data[78964] <= 8'h10 ;
			data[78965] <= 8'h10 ;
			data[78966] <= 8'h10 ;
			data[78967] <= 8'h10 ;
			data[78968] <= 8'h10 ;
			data[78969] <= 8'h10 ;
			data[78970] <= 8'h10 ;
			data[78971] <= 8'h10 ;
			data[78972] <= 8'h10 ;
			data[78973] <= 8'h10 ;
			data[78974] <= 8'h10 ;
			data[78975] <= 8'h10 ;
			data[78976] <= 8'h10 ;
			data[78977] <= 8'h10 ;
			data[78978] <= 8'h10 ;
			data[78979] <= 8'h10 ;
			data[78980] <= 8'h10 ;
			data[78981] <= 8'h10 ;
			data[78982] <= 8'h10 ;
			data[78983] <= 8'h10 ;
			data[78984] <= 8'h10 ;
			data[78985] <= 8'h10 ;
			data[78986] <= 8'h10 ;
			data[78987] <= 8'h10 ;
			data[78988] <= 8'h10 ;
			data[78989] <= 8'h10 ;
			data[78990] <= 8'h10 ;
			data[78991] <= 8'h10 ;
			data[78992] <= 8'h10 ;
			data[78993] <= 8'h10 ;
			data[78994] <= 8'h10 ;
			data[78995] <= 8'h10 ;
			data[78996] <= 8'h10 ;
			data[78997] <= 8'h10 ;
			data[78998] <= 8'h10 ;
			data[78999] <= 8'h10 ;
			data[79000] <= 8'h10 ;
			data[79001] <= 8'h10 ;
			data[79002] <= 8'h10 ;
			data[79003] <= 8'h10 ;
			data[79004] <= 8'h10 ;
			data[79005] <= 8'h10 ;
			data[79006] <= 8'h10 ;
			data[79007] <= 8'h10 ;
			data[79008] <= 8'h10 ;
			data[79009] <= 8'h10 ;
			data[79010] <= 8'h10 ;
			data[79011] <= 8'h10 ;
			data[79012] <= 8'h10 ;
			data[79013] <= 8'h10 ;
			data[79014] <= 8'h10 ;
			data[79015] <= 8'h10 ;
			data[79016] <= 8'h10 ;
			data[79017] <= 8'h10 ;
			data[79018] <= 8'h10 ;
			data[79019] <= 8'h10 ;
			data[79020] <= 8'h10 ;
			data[79021] <= 8'h10 ;
			data[79022] <= 8'h10 ;
			data[79023] <= 8'h10 ;
			data[79024] <= 8'h10 ;
			data[79025] <= 8'h10 ;
			data[79026] <= 8'h10 ;
			data[79027] <= 8'h10 ;
			data[79028] <= 8'h10 ;
			data[79029] <= 8'h10 ;
			data[79030] <= 8'h10 ;
			data[79031] <= 8'h10 ;
			data[79032] <= 8'h10 ;
			data[79033] <= 8'h10 ;
			data[79034] <= 8'h10 ;
			data[79035] <= 8'h10 ;
			data[79036] <= 8'h10 ;
			data[79037] <= 8'h10 ;
			data[79038] <= 8'h10 ;
			data[79039] <= 8'h10 ;
			data[79040] <= 8'h10 ;
			data[79041] <= 8'h10 ;
			data[79042] <= 8'h10 ;
			data[79043] <= 8'h10 ;
			data[79044] <= 8'h10 ;
			data[79045] <= 8'h10 ;
			data[79046] <= 8'h10 ;
			data[79047] <= 8'h10 ;
			data[79048] <= 8'h10 ;
			data[79049] <= 8'h10 ;
			data[79050] <= 8'h10 ;
			data[79051] <= 8'h10 ;
			data[79052] <= 8'h10 ;
			data[79053] <= 8'h10 ;
			data[79054] <= 8'h10 ;
			data[79055] <= 8'h10 ;
			data[79056] <= 8'h10 ;
			data[79057] <= 8'h10 ;
			data[79058] <= 8'h10 ;
			data[79059] <= 8'h10 ;
			data[79060] <= 8'h10 ;
			data[79061] <= 8'h10 ;
			data[79062] <= 8'h10 ;
			data[79063] <= 8'h10 ;
			data[79064] <= 8'h10 ;
			data[79065] <= 8'h10 ;
			data[79066] <= 8'h10 ;
			data[79067] <= 8'h10 ;
			data[79068] <= 8'h10 ;
			data[79069] <= 8'h10 ;
			data[79070] <= 8'h10 ;
			data[79071] <= 8'h10 ;
			data[79072] <= 8'h10 ;
			data[79073] <= 8'h10 ;
			data[79074] <= 8'h10 ;
			data[79075] <= 8'h10 ;
			data[79076] <= 8'h10 ;
			data[79077] <= 8'h10 ;
			data[79078] <= 8'h10 ;
			data[79079] <= 8'h10 ;
			data[79080] <= 8'h10 ;
			data[79081] <= 8'h10 ;
			data[79082] <= 8'h10 ;
			data[79083] <= 8'h10 ;
			data[79084] <= 8'h10 ;
			data[79085] <= 8'h10 ;
			data[79086] <= 8'h10 ;
			data[79087] <= 8'h10 ;
			data[79088] <= 8'h10 ;
			data[79089] <= 8'h10 ;
			data[79090] <= 8'h10 ;
			data[79091] <= 8'h10 ;
			data[79092] <= 8'h10 ;
			data[79093] <= 8'h10 ;
			data[79094] <= 8'h10 ;
			data[79095] <= 8'h10 ;
			data[79096] <= 8'h10 ;
			data[79097] <= 8'h10 ;
			data[79098] <= 8'h10 ;
			data[79099] <= 8'h10 ;
			data[79100] <= 8'h10 ;
			data[79101] <= 8'h10 ;
			data[79102] <= 8'h10 ;
			data[79103] <= 8'h10 ;
			data[79104] <= 8'h10 ;
			data[79105] <= 8'h10 ;
			data[79106] <= 8'h10 ;
			data[79107] <= 8'h10 ;
			data[79108] <= 8'h10 ;
			data[79109] <= 8'h10 ;
			data[79110] <= 8'h10 ;
			data[79111] <= 8'h10 ;
			data[79112] <= 8'h10 ;
			data[79113] <= 8'h10 ;
			data[79114] <= 8'h10 ;
			data[79115] <= 8'h10 ;
			data[79116] <= 8'h10 ;
			data[79117] <= 8'h10 ;
			data[79118] <= 8'h10 ;
			data[79119] <= 8'h10 ;
			data[79120] <= 8'h10 ;
			data[79121] <= 8'h10 ;
			data[79122] <= 8'h10 ;
			data[79123] <= 8'h10 ;
			data[79124] <= 8'h10 ;
			data[79125] <= 8'h10 ;
			data[79126] <= 8'h10 ;
			data[79127] <= 8'h10 ;
			data[79128] <= 8'h10 ;
			data[79129] <= 8'h10 ;
			data[79130] <= 8'h10 ;
			data[79131] <= 8'h10 ;
			data[79132] <= 8'h10 ;
			data[79133] <= 8'h10 ;
			data[79134] <= 8'h10 ;
			data[79135] <= 8'h10 ;
			data[79136] <= 8'h10 ;
			data[79137] <= 8'h10 ;
			data[79138] <= 8'h10 ;
			data[79139] <= 8'h10 ;
			data[79140] <= 8'h10 ;
			data[79141] <= 8'h10 ;
			data[79142] <= 8'h10 ;
			data[79143] <= 8'h10 ;
			data[79144] <= 8'h10 ;
			data[79145] <= 8'h10 ;
			data[79146] <= 8'h10 ;
			data[79147] <= 8'h10 ;
			data[79148] <= 8'h10 ;
			data[79149] <= 8'h10 ;
			data[79150] <= 8'h10 ;
			data[79151] <= 8'h10 ;
			data[79152] <= 8'h10 ;
			data[79153] <= 8'h10 ;
			data[79154] <= 8'h10 ;
			data[79155] <= 8'h10 ;
			data[79156] <= 8'h10 ;
			data[79157] <= 8'h10 ;
			data[79158] <= 8'h10 ;
			data[79159] <= 8'h10 ;
			data[79160] <= 8'h10 ;
			data[79161] <= 8'h10 ;
			data[79162] <= 8'h10 ;
			data[79163] <= 8'h10 ;
			data[79164] <= 8'h10 ;
			data[79165] <= 8'h10 ;
			data[79166] <= 8'h10 ;
			data[79167] <= 8'h10 ;
			data[79168] <= 8'h10 ;
			data[79169] <= 8'h10 ;
			data[79170] <= 8'h10 ;
			data[79171] <= 8'h10 ;
			data[79172] <= 8'h10 ;
			data[79173] <= 8'h10 ;
			data[79174] <= 8'h10 ;
			data[79175] <= 8'h10 ;
			data[79176] <= 8'h10 ;
			data[79177] <= 8'h10 ;
			data[79178] <= 8'h10 ;
			data[79179] <= 8'h10 ;
			data[79180] <= 8'h10 ;
			data[79181] <= 8'h10 ;
			data[79182] <= 8'h10 ;
			data[79183] <= 8'h10 ;
			data[79184] <= 8'h10 ;
			data[79185] <= 8'h10 ;
			data[79186] <= 8'h10 ;
			data[79187] <= 8'h10 ;
			data[79188] <= 8'h10 ;
			data[79189] <= 8'h10 ;
			data[79190] <= 8'h10 ;
			data[79191] <= 8'h10 ;
			data[79192] <= 8'h10 ;
			data[79193] <= 8'h10 ;
			data[79194] <= 8'h10 ;
			data[79195] <= 8'h10 ;
			data[79196] <= 8'h10 ;
			data[79197] <= 8'h10 ;
			data[79198] <= 8'h10 ;
			data[79199] <= 8'h10 ;
			data[79200] <= 8'h10 ;
			data[79201] <= 8'h10 ;
			data[79202] <= 8'h10 ;
			data[79203] <= 8'h10 ;
			data[79204] <= 8'h10 ;
			data[79205] <= 8'h10 ;
			data[79206] <= 8'h10 ;
			data[79207] <= 8'h10 ;
			data[79208] <= 8'h10 ;
			data[79209] <= 8'h10 ;
			data[79210] <= 8'h10 ;
			data[79211] <= 8'h10 ;
			data[79212] <= 8'h10 ;
			data[79213] <= 8'h10 ;
			data[79214] <= 8'h10 ;
			data[79215] <= 8'h10 ;
			data[79216] <= 8'h10 ;
			data[79217] <= 8'h10 ;
			data[79218] <= 8'h10 ;
			data[79219] <= 8'h10 ;
			data[79220] <= 8'h10 ;
			data[79221] <= 8'h10 ;
			data[79222] <= 8'h10 ;
			data[79223] <= 8'h10 ;
			data[79224] <= 8'h10 ;
			data[79225] <= 8'h10 ;
			data[79226] <= 8'h10 ;
			data[79227] <= 8'h10 ;
			data[79228] <= 8'h10 ;
			data[79229] <= 8'h10 ;
			data[79230] <= 8'h10 ;
			data[79231] <= 8'h10 ;
			data[79232] <= 8'h10 ;
			data[79233] <= 8'h10 ;
			data[79234] <= 8'h10 ;
			data[79235] <= 8'h10 ;
			data[79236] <= 8'h10 ;
			data[79237] <= 8'h10 ;
			data[79238] <= 8'h10 ;
			data[79239] <= 8'h10 ;
			data[79240] <= 8'h10 ;
			data[79241] <= 8'h10 ;
			data[79242] <= 8'h10 ;
			data[79243] <= 8'h10 ;
			data[79244] <= 8'h10 ;
			data[79245] <= 8'h10 ;
			data[79246] <= 8'h10 ;
			data[79247] <= 8'h10 ;
			data[79248] <= 8'h10 ;
			data[79249] <= 8'h10 ;
			data[79250] <= 8'h10 ;
			data[79251] <= 8'h10 ;
			data[79252] <= 8'h10 ;
			data[79253] <= 8'h10 ;
			data[79254] <= 8'h10 ;
			data[79255] <= 8'h10 ;
			data[79256] <= 8'h10 ;
			data[79257] <= 8'h10 ;
			data[79258] <= 8'h10 ;
			data[79259] <= 8'h10 ;
			data[79260] <= 8'h10 ;
			data[79261] <= 8'h10 ;
			data[79262] <= 8'h10 ;
			data[79263] <= 8'h10 ;
			data[79264] <= 8'h10 ;
			data[79265] <= 8'h10 ;
			data[79266] <= 8'h10 ;
			data[79267] <= 8'h10 ;
			data[79268] <= 8'h10 ;
			data[79269] <= 8'h10 ;
			data[79270] <= 8'h10 ;
			data[79271] <= 8'h10 ;
			data[79272] <= 8'h10 ;
			data[79273] <= 8'h10 ;
			data[79274] <= 8'h10 ;
			data[79275] <= 8'h10 ;
			data[79276] <= 8'h10 ;
			data[79277] <= 8'h10 ;
			data[79278] <= 8'h10 ;
			data[79279] <= 8'h10 ;
			data[79280] <= 8'h10 ;
			data[79281] <= 8'h10 ;
			data[79282] <= 8'h10 ;
			data[79283] <= 8'h10 ;
			data[79284] <= 8'h10 ;
			data[79285] <= 8'h10 ;
			data[79286] <= 8'h10 ;
			data[79287] <= 8'h10 ;
			data[79288] <= 8'h10 ;
			data[79289] <= 8'h10 ;
			data[79290] <= 8'h10 ;
			data[79291] <= 8'h10 ;
			data[79292] <= 8'h10 ;
			data[79293] <= 8'h10 ;
			data[79294] <= 8'h10 ;
			data[79295] <= 8'h10 ;
			data[79296] <= 8'h10 ;
			data[79297] <= 8'h10 ;
			data[79298] <= 8'h10 ;
			data[79299] <= 8'h10 ;
			data[79300] <= 8'h10 ;
			data[79301] <= 8'h10 ;
			data[79302] <= 8'h10 ;
			data[79303] <= 8'h10 ;
			data[79304] <= 8'h10 ;
			data[79305] <= 8'h10 ;
			data[79306] <= 8'h10 ;
			data[79307] <= 8'h10 ;
			data[79308] <= 8'h10 ;
			data[79309] <= 8'h10 ;
			data[79310] <= 8'h10 ;
			data[79311] <= 8'h10 ;
			data[79312] <= 8'h10 ;
			data[79313] <= 8'h10 ;
			data[79314] <= 8'h10 ;
			data[79315] <= 8'h10 ;
			data[79316] <= 8'h10 ;
			data[79317] <= 8'h10 ;
			data[79318] <= 8'h10 ;
			data[79319] <= 8'h10 ;
			data[79320] <= 8'h10 ;
			data[79321] <= 8'h10 ;
			data[79322] <= 8'h10 ;
			data[79323] <= 8'h10 ;
			data[79324] <= 8'h10 ;
			data[79325] <= 8'h10 ;
			data[79326] <= 8'h10 ;
			data[79327] <= 8'h10 ;
			data[79328] <= 8'h10 ;
			data[79329] <= 8'h10 ;
			data[79330] <= 8'h10 ;
			data[79331] <= 8'h10 ;
			data[79332] <= 8'h10 ;
			data[79333] <= 8'h10 ;
			data[79334] <= 8'h10 ;
			data[79335] <= 8'h10 ;
			data[79336] <= 8'h10 ;
			data[79337] <= 8'h10 ;
			data[79338] <= 8'h10 ;
			data[79339] <= 8'h10 ;
			data[79340] <= 8'h10 ;
			data[79341] <= 8'h10 ;
			data[79342] <= 8'h10 ;
			data[79343] <= 8'h10 ;
			data[79344] <= 8'h10 ;
			data[79345] <= 8'h10 ;
			data[79346] <= 8'h10 ;
			data[79347] <= 8'h10 ;
			data[79348] <= 8'h10 ;
			data[79349] <= 8'h10 ;
			data[79350] <= 8'h10 ;
			data[79351] <= 8'h10 ;
			data[79352] <= 8'h10 ;
			data[79353] <= 8'h10 ;
			data[79354] <= 8'h10 ;
			data[79355] <= 8'h10 ;
			data[79356] <= 8'h10 ;
			data[79357] <= 8'h10 ;
			data[79358] <= 8'h10 ;
			data[79359] <= 8'h10 ;
			data[79360] <= 8'h10 ;
			data[79361] <= 8'h10 ;
			data[79362] <= 8'h10 ;
			data[79363] <= 8'h10 ;
			data[79364] <= 8'h10 ;
			data[79365] <= 8'h10 ;
			data[79366] <= 8'h10 ;
			data[79367] <= 8'h10 ;
			data[79368] <= 8'h10 ;
			data[79369] <= 8'h10 ;
			data[79370] <= 8'h10 ;
			data[79371] <= 8'h10 ;
			data[79372] <= 8'h10 ;
			data[79373] <= 8'h10 ;
			data[79374] <= 8'h10 ;
			data[79375] <= 8'h10 ;
			data[79376] <= 8'h10 ;
			data[79377] <= 8'h10 ;
			data[79378] <= 8'h10 ;
			data[79379] <= 8'h10 ;
			data[79380] <= 8'h10 ;
			data[79381] <= 8'h10 ;
			data[79382] <= 8'h10 ;
			data[79383] <= 8'h10 ;
			data[79384] <= 8'h10 ;
			data[79385] <= 8'h10 ;
			data[79386] <= 8'h10 ;
			data[79387] <= 8'h10 ;
			data[79388] <= 8'h10 ;
			data[79389] <= 8'h10 ;
			data[79390] <= 8'h10 ;
			data[79391] <= 8'h10 ;
			data[79392] <= 8'h10 ;
			data[79393] <= 8'h10 ;
			data[79394] <= 8'h10 ;
			data[79395] <= 8'h10 ;
			data[79396] <= 8'h10 ;
			data[79397] <= 8'h10 ;
			data[79398] <= 8'h10 ;
			data[79399] <= 8'h10 ;
			data[79400] <= 8'h10 ;
			data[79401] <= 8'h10 ;
			data[79402] <= 8'h10 ;
			data[79403] <= 8'h10 ;
			data[79404] <= 8'h10 ;
			data[79405] <= 8'h10 ;
			data[79406] <= 8'h10 ;
			data[79407] <= 8'h10 ;
			data[79408] <= 8'h10 ;
			data[79409] <= 8'h10 ;
			data[79410] <= 8'h10 ;
			data[79411] <= 8'h10 ;
			data[79412] <= 8'h10 ;
			data[79413] <= 8'h10 ;
			data[79414] <= 8'h10 ;
			data[79415] <= 8'h10 ;
			data[79416] <= 8'h10 ;
			data[79417] <= 8'h10 ;
			data[79418] <= 8'h10 ;
			data[79419] <= 8'h10 ;
			data[79420] <= 8'h10 ;
			data[79421] <= 8'h10 ;
			data[79422] <= 8'h10 ;
			data[79423] <= 8'h10 ;
			data[79424] <= 8'h10 ;
			data[79425] <= 8'h10 ;
			data[79426] <= 8'h10 ;
			data[79427] <= 8'h10 ;
			data[79428] <= 8'h10 ;
			data[79429] <= 8'h10 ;
			data[79430] <= 8'h10 ;
			data[79431] <= 8'h10 ;
			data[79432] <= 8'h10 ;
			data[79433] <= 8'h10 ;
			data[79434] <= 8'h10 ;
			data[79435] <= 8'h10 ;
			data[79436] <= 8'h10 ;
			data[79437] <= 8'h10 ;
			data[79438] <= 8'h10 ;
			data[79439] <= 8'h10 ;
			data[79440] <= 8'h10 ;
			data[79441] <= 8'h10 ;
			data[79442] <= 8'h10 ;
			data[79443] <= 8'h10 ;
			data[79444] <= 8'h10 ;
			data[79445] <= 8'h10 ;
			data[79446] <= 8'h10 ;
			data[79447] <= 8'h10 ;
			data[79448] <= 8'h10 ;
			data[79449] <= 8'h10 ;
			data[79450] <= 8'h10 ;
			data[79451] <= 8'h10 ;
			data[79452] <= 8'h10 ;
			data[79453] <= 8'h10 ;
			data[79454] <= 8'h10 ;
			data[79455] <= 8'h10 ;
			data[79456] <= 8'h10 ;
			data[79457] <= 8'h10 ;
			data[79458] <= 8'h10 ;
			data[79459] <= 8'h10 ;
			data[79460] <= 8'h10 ;
			data[79461] <= 8'h10 ;
			data[79462] <= 8'h10 ;
			data[79463] <= 8'h10 ;
			data[79464] <= 8'h10 ;
			data[79465] <= 8'h10 ;
			data[79466] <= 8'h10 ;
			data[79467] <= 8'h10 ;
			data[79468] <= 8'h10 ;
			data[79469] <= 8'h10 ;
			data[79470] <= 8'h10 ;
			data[79471] <= 8'h10 ;
			data[79472] <= 8'h10 ;
			data[79473] <= 8'h10 ;
			data[79474] <= 8'h10 ;
			data[79475] <= 8'h10 ;
			data[79476] <= 8'h10 ;
			data[79477] <= 8'h10 ;
			data[79478] <= 8'h10 ;
			data[79479] <= 8'h10 ;
			data[79480] <= 8'h10 ;
			data[79481] <= 8'h10 ;
			data[79482] <= 8'h10 ;
			data[79483] <= 8'h10 ;
			data[79484] <= 8'h10 ;
			data[79485] <= 8'h10 ;
			data[79486] <= 8'h10 ;
			data[79487] <= 8'h10 ;
			data[79488] <= 8'h10 ;
			data[79489] <= 8'h10 ;
			data[79490] <= 8'h10 ;
			data[79491] <= 8'h10 ;
			data[79492] <= 8'h10 ;
			data[79493] <= 8'h10 ;
			data[79494] <= 8'h10 ;
			data[79495] <= 8'h10 ;
			data[79496] <= 8'h10 ;
			data[79497] <= 8'h10 ;
			data[79498] <= 8'h10 ;
			data[79499] <= 8'h10 ;
			data[79500] <= 8'h10 ;
			data[79501] <= 8'h10 ;
			data[79502] <= 8'h10 ;
			data[79503] <= 8'h10 ;
			data[79504] <= 8'h10 ;
			data[79505] <= 8'h10 ;
			data[79506] <= 8'h10 ;
			data[79507] <= 8'h10 ;
			data[79508] <= 8'h10 ;
			data[79509] <= 8'h10 ;
			data[79510] <= 8'h10 ;
			data[79511] <= 8'h10 ;
			data[79512] <= 8'h10 ;
			data[79513] <= 8'h10 ;
			data[79514] <= 8'h10 ;
			data[79515] <= 8'h10 ;
			data[79516] <= 8'h10 ;
			data[79517] <= 8'h10 ;
			data[79518] <= 8'h10 ;
			data[79519] <= 8'h10 ;
			data[79520] <= 8'h10 ;
			data[79521] <= 8'h10 ;
			data[79522] <= 8'h10 ;
			data[79523] <= 8'h10 ;
			data[79524] <= 8'h10 ;
			data[79525] <= 8'h10 ;
			data[79526] <= 8'h10 ;
			data[79527] <= 8'h10 ;
			data[79528] <= 8'h10 ;
			data[79529] <= 8'h10 ;
			data[79530] <= 8'h10 ;
			data[79531] <= 8'h10 ;
			data[79532] <= 8'h10 ;
			data[79533] <= 8'h10 ;
			data[79534] <= 8'h10 ;
			data[79535] <= 8'h10 ;
			data[79536] <= 8'h10 ;
			data[79537] <= 8'h10 ;
			data[79538] <= 8'h10 ;
			data[79539] <= 8'h10 ;
			data[79540] <= 8'h10 ;
			data[79541] <= 8'h10 ;
			data[79542] <= 8'h10 ;
			data[79543] <= 8'h10 ;
			data[79544] <= 8'h10 ;
			data[79545] <= 8'h10 ;
			data[79546] <= 8'h10 ;
			data[79547] <= 8'h10 ;
			data[79548] <= 8'h10 ;
			data[79549] <= 8'h10 ;
			data[79550] <= 8'h10 ;
			data[79551] <= 8'h10 ;
			data[79552] <= 8'h10 ;
			data[79553] <= 8'h10 ;
			data[79554] <= 8'h10 ;
			data[79555] <= 8'h10 ;
			data[79556] <= 8'h10 ;
			data[79557] <= 8'h10 ;
			data[79558] <= 8'h10 ;
			data[79559] <= 8'h10 ;
			data[79560] <= 8'h10 ;
			data[79561] <= 8'h10 ;
			data[79562] <= 8'h10 ;
			data[79563] <= 8'h10 ;
			data[79564] <= 8'h10 ;
			data[79565] <= 8'h10 ;
			data[79566] <= 8'h10 ;
			data[79567] <= 8'h10 ;
			data[79568] <= 8'h10 ;
			data[79569] <= 8'h10 ;
			data[79570] <= 8'h10 ;
			data[79571] <= 8'h10 ;
			data[79572] <= 8'h10 ;
			data[79573] <= 8'h10 ;
			data[79574] <= 8'h10 ;
			data[79575] <= 8'h10 ;
			data[79576] <= 8'h10 ;
			data[79577] <= 8'h10 ;
			data[79578] <= 8'h10 ;
			data[79579] <= 8'h10 ;
			data[79580] <= 8'h10 ;
			data[79581] <= 8'h10 ;
			data[79582] <= 8'h10 ;
			data[79583] <= 8'h10 ;
			data[79584] <= 8'h10 ;
			data[79585] <= 8'h10 ;
			data[79586] <= 8'h10 ;
			data[79587] <= 8'h10 ;
			data[79588] <= 8'h10 ;
			data[79589] <= 8'h10 ;
			data[79590] <= 8'h10 ;
			data[79591] <= 8'h10 ;
			data[79592] <= 8'h10 ;
			data[79593] <= 8'h10 ;
			data[79594] <= 8'h10 ;
			data[79595] <= 8'h10 ;
			data[79596] <= 8'h10 ;
			data[79597] <= 8'h10 ;
			data[79598] <= 8'h10 ;
			data[79599] <= 8'h10 ;
			data[79600] <= 8'h10 ;
			data[79601] <= 8'h10 ;
			data[79602] <= 8'h10 ;
			data[79603] <= 8'h10 ;
			data[79604] <= 8'h10 ;
			data[79605] <= 8'h10 ;
			data[79606] <= 8'h10 ;
			data[79607] <= 8'h10 ;
			data[79608] <= 8'h10 ;
			data[79609] <= 8'h10 ;
			data[79610] <= 8'h10 ;
			data[79611] <= 8'h10 ;
			data[79612] <= 8'h10 ;
			data[79613] <= 8'h10 ;
			data[79614] <= 8'h10 ;
			data[79615] <= 8'h10 ;
			data[79616] <= 8'h10 ;
			data[79617] <= 8'h10 ;
			data[79618] <= 8'h10 ;
			data[79619] <= 8'h10 ;
			data[79620] <= 8'h10 ;
			data[79621] <= 8'h10 ;
			data[79622] <= 8'h10 ;
			data[79623] <= 8'h10 ;
			data[79624] <= 8'h10 ;
			data[79625] <= 8'h10 ;
			data[79626] <= 8'h10 ;
			data[79627] <= 8'h10 ;
			data[79628] <= 8'h10 ;
			data[79629] <= 8'h10 ;
			data[79630] <= 8'h10 ;
			data[79631] <= 8'h10 ;
			data[79632] <= 8'h10 ;
			data[79633] <= 8'h10 ;
			data[79634] <= 8'h10 ;
			data[79635] <= 8'h10 ;
			data[79636] <= 8'h10 ;
			data[79637] <= 8'h10 ;
			data[79638] <= 8'h10 ;
			data[79639] <= 8'h10 ;
			data[79640] <= 8'h10 ;
			data[79641] <= 8'h10 ;
			data[79642] <= 8'h10 ;
			data[79643] <= 8'h10 ;
			data[79644] <= 8'h10 ;
			data[79645] <= 8'h10 ;
			data[79646] <= 8'h10 ;
			data[79647] <= 8'h10 ;
			data[79648] <= 8'h10 ;
			data[79649] <= 8'h10 ;
			data[79650] <= 8'h10 ;
			data[79651] <= 8'h10 ;
			data[79652] <= 8'h10 ;
			data[79653] <= 8'h10 ;
			data[79654] <= 8'h10 ;
			data[79655] <= 8'h10 ;
			data[79656] <= 8'h10 ;
			data[79657] <= 8'h10 ;
			data[79658] <= 8'h10 ;
			data[79659] <= 8'h10 ;
			data[79660] <= 8'h10 ;
			data[79661] <= 8'h10 ;
			data[79662] <= 8'h10 ;
			data[79663] <= 8'h10 ;
			data[79664] <= 8'h10 ;
			data[79665] <= 8'h10 ;
			data[79666] <= 8'h10 ;
			data[79667] <= 8'h10 ;
			data[79668] <= 8'h10 ;
			data[79669] <= 8'h10 ;
			data[79670] <= 8'h10 ;
			data[79671] <= 8'h10 ;
			data[79672] <= 8'h10 ;
			data[79673] <= 8'h10 ;
			data[79674] <= 8'h10 ;
			data[79675] <= 8'h10 ;
			data[79676] <= 8'h10 ;
			data[79677] <= 8'h10 ;
			data[79678] <= 8'h10 ;
			data[79679] <= 8'h10 ;
			data[79680] <= 8'h10 ;
			data[79681] <= 8'h10 ;
			data[79682] <= 8'h10 ;
			data[79683] <= 8'h10 ;
			data[79684] <= 8'h10 ;
			data[79685] <= 8'h10 ;
			data[79686] <= 8'h10 ;
			data[79687] <= 8'h10 ;
			data[79688] <= 8'h10 ;
			data[79689] <= 8'h10 ;
			data[79690] <= 8'h10 ;
			data[79691] <= 8'h10 ;
			data[79692] <= 8'h10 ;
			data[79693] <= 8'h10 ;
			data[79694] <= 8'h10 ;
			data[79695] <= 8'h10 ;
			data[79696] <= 8'h10 ;
			data[79697] <= 8'h10 ;
			data[79698] <= 8'h10 ;
			data[79699] <= 8'h10 ;
			data[79700] <= 8'h10 ;
			data[79701] <= 8'h10 ;
			data[79702] <= 8'h10 ;
			data[79703] <= 8'h10 ;
			data[79704] <= 8'h10 ;
			data[79705] <= 8'h10 ;
			data[79706] <= 8'h10 ;
			data[79707] <= 8'h10 ;
			data[79708] <= 8'h10 ;
			data[79709] <= 8'h10 ;
			data[79710] <= 8'h10 ;
			data[79711] <= 8'h10 ;
			data[79712] <= 8'h10 ;
			data[79713] <= 8'h10 ;
			data[79714] <= 8'h10 ;
			data[79715] <= 8'h10 ;
			data[79716] <= 8'h10 ;
			data[79717] <= 8'h10 ;
			data[79718] <= 8'h10 ;
			data[79719] <= 8'h10 ;
			data[79720] <= 8'h10 ;
			data[79721] <= 8'h10 ;
			data[79722] <= 8'h10 ;
			data[79723] <= 8'h10 ;
			data[79724] <= 8'h10 ;
			data[79725] <= 8'h10 ;
			data[79726] <= 8'h10 ;
			data[79727] <= 8'h10 ;
			data[79728] <= 8'h10 ;
			data[79729] <= 8'h10 ;
			data[79730] <= 8'h10 ;
			data[79731] <= 8'h10 ;
			data[79732] <= 8'h10 ;
			data[79733] <= 8'h10 ;
			data[79734] <= 8'h10 ;
			data[79735] <= 8'h10 ;
			data[79736] <= 8'h10 ;
			data[79737] <= 8'h10 ;
			data[79738] <= 8'h10 ;
			data[79739] <= 8'h10 ;
			data[79740] <= 8'h10 ;
			data[79741] <= 8'h10 ;
			data[79742] <= 8'h10 ;
			data[79743] <= 8'h10 ;
			data[79744] <= 8'h10 ;
			data[79745] <= 8'h10 ;
			data[79746] <= 8'h10 ;
			data[79747] <= 8'h10 ;
			data[79748] <= 8'h10 ;
			data[79749] <= 8'h10 ;
			data[79750] <= 8'h10 ;
			data[79751] <= 8'h10 ;
			data[79752] <= 8'h10 ;
			data[79753] <= 8'h10 ;
			data[79754] <= 8'h10 ;
			data[79755] <= 8'h10 ;
			data[79756] <= 8'h10 ;
			data[79757] <= 8'h10 ;
			data[79758] <= 8'h10 ;
			data[79759] <= 8'h10 ;
			data[79760] <= 8'h10 ;
			data[79761] <= 8'h10 ;
			data[79762] <= 8'h10 ;
			data[79763] <= 8'h10 ;
			data[79764] <= 8'h10 ;
			data[79765] <= 8'h10 ;
			data[79766] <= 8'h10 ;
			data[79767] <= 8'h10 ;
			data[79768] <= 8'h10 ;
			data[79769] <= 8'h10 ;
			data[79770] <= 8'h10 ;
			data[79771] <= 8'h10 ;
			data[79772] <= 8'h10 ;
			data[79773] <= 8'h10 ;
			data[79774] <= 8'h10 ;
			data[79775] <= 8'h10 ;
			data[79776] <= 8'h10 ;
			data[79777] <= 8'h10 ;
			data[79778] <= 8'h10 ;
			data[79779] <= 8'h10 ;
			data[79780] <= 8'h10 ;
			data[79781] <= 8'h10 ;
			data[79782] <= 8'h10 ;
			data[79783] <= 8'h10 ;
			data[79784] <= 8'h10 ;
			data[79785] <= 8'h10 ;
			data[79786] <= 8'h10 ;
			data[79787] <= 8'h10 ;
			data[79788] <= 8'h10 ;
			data[79789] <= 8'h10 ;
			data[79790] <= 8'h10 ;
			data[79791] <= 8'h10 ;
			data[79792] <= 8'h10 ;
			data[79793] <= 8'h10 ;
			data[79794] <= 8'h10 ;
			data[79795] <= 8'h10 ;
			data[79796] <= 8'h10 ;
			data[79797] <= 8'h10 ;
			data[79798] <= 8'h10 ;
			data[79799] <= 8'h10 ;
			data[79800] <= 8'h10 ;
			data[79801] <= 8'h10 ;
			data[79802] <= 8'h10 ;
			data[79803] <= 8'h10 ;
			data[79804] <= 8'h10 ;
			data[79805] <= 8'h10 ;
			data[79806] <= 8'h10 ;
			data[79807] <= 8'h10 ;
			data[79808] <= 8'h10 ;
			data[79809] <= 8'h10 ;
			data[79810] <= 8'h10 ;
			data[79811] <= 8'h10 ;
			data[79812] <= 8'h10 ;
			data[79813] <= 8'h10 ;
			data[79814] <= 8'h10 ;
			data[79815] <= 8'h10 ;
			data[79816] <= 8'h10 ;
			data[79817] <= 8'h10 ;
			data[79818] <= 8'h10 ;
			data[79819] <= 8'h10 ;
			data[79820] <= 8'h10 ;
			data[79821] <= 8'h10 ;
			data[79822] <= 8'h10 ;
			data[79823] <= 8'h10 ;
			data[79824] <= 8'h10 ;
			data[79825] <= 8'h10 ;
			data[79826] <= 8'h10 ;
			data[79827] <= 8'h10 ;
			data[79828] <= 8'h10 ;
			data[79829] <= 8'h10 ;
			data[79830] <= 8'h10 ;
			data[79831] <= 8'h10 ;
			data[79832] <= 8'h10 ;
			data[79833] <= 8'h10 ;
			data[79834] <= 8'h10 ;
			data[79835] <= 8'h10 ;
			data[79836] <= 8'h10 ;
			data[79837] <= 8'h10 ;
			data[79838] <= 8'h10 ;
			data[79839] <= 8'h10 ;
			data[79840] <= 8'h10 ;
			data[79841] <= 8'h10 ;
			data[79842] <= 8'h10 ;
			data[79843] <= 8'h10 ;
			data[79844] <= 8'h10 ;
			data[79845] <= 8'h10 ;
			data[79846] <= 8'h10 ;
			data[79847] <= 8'h10 ;
			data[79848] <= 8'h10 ;
			data[79849] <= 8'h10 ;
			data[79850] <= 8'h10 ;
			data[79851] <= 8'h10 ;
			data[79852] <= 8'h10 ;
			data[79853] <= 8'h10 ;
			data[79854] <= 8'h10 ;
			data[79855] <= 8'h10 ;
			data[79856] <= 8'h10 ;
			data[79857] <= 8'h10 ;
			data[79858] <= 8'h10 ;
			data[79859] <= 8'h10 ;
			data[79860] <= 8'h10 ;
			data[79861] <= 8'h10 ;
			data[79862] <= 8'h10 ;
			data[79863] <= 8'h10 ;
			data[79864] <= 8'h10 ;
			data[79865] <= 8'h10 ;
			data[79866] <= 8'h10 ;
			data[79867] <= 8'h10 ;
			data[79868] <= 8'h10 ;
			data[79869] <= 8'h10 ;
			data[79870] <= 8'h10 ;
			data[79871] <= 8'h10 ;
			data[79872] <= 8'h10 ;
			data[79873] <= 8'h10 ;
			data[79874] <= 8'h10 ;
			data[79875] <= 8'h10 ;
			data[79876] <= 8'h10 ;
			data[79877] <= 8'h10 ;
			data[79878] <= 8'h10 ;
			data[79879] <= 8'h10 ;
			data[79880] <= 8'h10 ;
			data[79881] <= 8'h10 ;
			data[79882] <= 8'h10 ;
			data[79883] <= 8'h10 ;
			data[79884] <= 8'h10 ;
			data[79885] <= 8'h10 ;
			data[79886] <= 8'h10 ;
			data[79887] <= 8'h10 ;
			data[79888] <= 8'h10 ;
			data[79889] <= 8'h10 ;
			data[79890] <= 8'h10 ;
			data[79891] <= 8'h10 ;
			data[79892] <= 8'h10 ;
			data[79893] <= 8'h10 ;
			data[79894] <= 8'h10 ;
			data[79895] <= 8'h10 ;
			data[79896] <= 8'h10 ;
			data[79897] <= 8'h10 ;
			data[79898] <= 8'h10 ;
			data[79899] <= 8'h10 ;
			data[79900] <= 8'h10 ;
			data[79901] <= 8'h10 ;
			data[79902] <= 8'h10 ;
			data[79903] <= 8'h10 ;
			data[79904] <= 8'h10 ;
			data[79905] <= 8'h10 ;
			data[79906] <= 8'h10 ;
			data[79907] <= 8'h10 ;
			data[79908] <= 8'h10 ;
			data[79909] <= 8'h10 ;
			data[79910] <= 8'h10 ;
			data[79911] <= 8'h10 ;
			data[79912] <= 8'h10 ;
			data[79913] <= 8'h10 ;
			data[79914] <= 8'h10 ;
			data[79915] <= 8'h10 ;
			data[79916] <= 8'h10 ;
			data[79917] <= 8'h10 ;
			data[79918] <= 8'h10 ;
			data[79919] <= 8'h10 ;
			data[79920] <= 8'h10 ;
			data[79921] <= 8'h10 ;
			data[79922] <= 8'h10 ;
			data[79923] <= 8'h10 ;
			data[79924] <= 8'h10 ;
			data[79925] <= 8'h10 ;
			data[79926] <= 8'h10 ;
			data[79927] <= 8'h10 ;
			data[79928] <= 8'h10 ;
			data[79929] <= 8'h10 ;
			data[79930] <= 8'h10 ;
			data[79931] <= 8'h10 ;
			data[79932] <= 8'h10 ;
			data[79933] <= 8'h10 ;
			data[79934] <= 8'h10 ;
			data[79935] <= 8'h10 ;
			data[79936] <= 8'h10 ;
			data[79937] <= 8'h10 ;
			data[79938] <= 8'h10 ;
			data[79939] <= 8'h10 ;
			data[79940] <= 8'h10 ;
			data[79941] <= 8'h10 ;
			data[79942] <= 8'h10 ;
			data[79943] <= 8'h10 ;
			data[79944] <= 8'h10 ;
			data[79945] <= 8'h10 ;
			data[79946] <= 8'h10 ;
			data[79947] <= 8'h10 ;
			data[79948] <= 8'h10 ;
			data[79949] <= 8'h10 ;
			data[79950] <= 8'h10 ;
			data[79951] <= 8'h10 ;
			data[79952] <= 8'h10 ;
			data[79953] <= 8'h10 ;
			data[79954] <= 8'h10 ;
			data[79955] <= 8'h10 ;
			data[79956] <= 8'h10 ;
			data[79957] <= 8'h10 ;
			data[79958] <= 8'h10 ;
			data[79959] <= 8'h10 ;
			data[79960] <= 8'h10 ;
			data[79961] <= 8'h10 ;
			data[79962] <= 8'h10 ;
			data[79963] <= 8'h10 ;
			data[79964] <= 8'h10 ;
			data[79965] <= 8'h10 ;
			data[79966] <= 8'h10 ;
			data[79967] <= 8'h10 ;
			data[79968] <= 8'h10 ;
			data[79969] <= 8'h10 ;
			data[79970] <= 8'h10 ;
			data[79971] <= 8'h10 ;
			data[79972] <= 8'h10 ;
			data[79973] <= 8'h10 ;
			data[79974] <= 8'h10 ;
			data[79975] <= 8'h10 ;
			data[79976] <= 8'h10 ;
			data[79977] <= 8'h10 ;
			data[79978] <= 8'h10 ;
			data[79979] <= 8'h10 ;
			data[79980] <= 8'h10 ;
			data[79981] <= 8'h10 ;
			data[79982] <= 8'h10 ;
			data[79983] <= 8'h10 ;
			data[79984] <= 8'h10 ;
			data[79985] <= 8'h10 ;
			data[79986] <= 8'h10 ;
			data[79987] <= 8'h10 ;
			data[79988] <= 8'h10 ;
			data[79989] <= 8'h10 ;
			data[79990] <= 8'h10 ;
			data[79991] <= 8'h10 ;
			data[79992] <= 8'h10 ;
			data[79993] <= 8'h10 ;
			data[79994] <= 8'h10 ;
			data[79995] <= 8'h10 ;
			data[79996] <= 8'h10 ;
			data[79997] <= 8'h10 ;
			data[79998] <= 8'h10 ;
			data[79999] <= 8'h10 ;
			data[80000] <= 8'h10 ;
			data[80001] <= 8'h10 ;
			data[80002] <= 8'h10 ;
			data[80003] <= 8'h10 ;
			data[80004] <= 8'h10 ;
			data[80005] <= 8'h10 ;
			data[80006] <= 8'h10 ;
			data[80007] <= 8'h10 ;
			data[80008] <= 8'h10 ;
			data[80009] <= 8'h10 ;
			data[80010] <= 8'h10 ;
			data[80011] <= 8'h10 ;
			data[80012] <= 8'h10 ;
			data[80013] <= 8'h10 ;
			data[80014] <= 8'h10 ;
			data[80015] <= 8'h10 ;
			data[80016] <= 8'h10 ;
			data[80017] <= 8'h10 ;
			data[80018] <= 8'h10 ;
			data[80019] <= 8'h10 ;
			data[80020] <= 8'h10 ;
			data[80021] <= 8'h10 ;
			data[80022] <= 8'h10 ;
			data[80023] <= 8'h10 ;
			data[80024] <= 8'h10 ;
			data[80025] <= 8'h10 ;
			data[80026] <= 8'h10 ;
			data[80027] <= 8'h10 ;
			data[80028] <= 8'h10 ;
			data[80029] <= 8'h10 ;
			data[80030] <= 8'h10 ;
			data[80031] <= 8'h10 ;
			data[80032] <= 8'h10 ;
			data[80033] <= 8'h10 ;
			data[80034] <= 8'h10 ;
			data[80035] <= 8'h10 ;
			data[80036] <= 8'h10 ;
			data[80037] <= 8'h10 ;
			data[80038] <= 8'h10 ;
			data[80039] <= 8'h10 ;
			data[80040] <= 8'h10 ;
			data[80041] <= 8'h10 ;
			data[80042] <= 8'h10 ;
			data[80043] <= 8'h10 ;
			data[80044] <= 8'h10 ;
			data[80045] <= 8'h10 ;
			data[80046] <= 8'h10 ;
			data[80047] <= 8'h10 ;
			data[80048] <= 8'h10 ;
			data[80049] <= 8'h10 ;
			data[80050] <= 8'h10 ;
			data[80051] <= 8'h10 ;
			data[80052] <= 8'h10 ;
			data[80053] <= 8'h10 ;
			data[80054] <= 8'h10 ;
			data[80055] <= 8'h10 ;
			data[80056] <= 8'h10 ;
			data[80057] <= 8'h10 ;
			data[80058] <= 8'h10 ;
			data[80059] <= 8'h10 ;
			data[80060] <= 8'h10 ;
			data[80061] <= 8'h10 ;
			data[80062] <= 8'h10 ;
			data[80063] <= 8'h10 ;
			data[80064] <= 8'h10 ;
			data[80065] <= 8'h10 ;
			data[80066] <= 8'h10 ;
			data[80067] <= 8'h10 ;
			data[80068] <= 8'h10 ;
			data[80069] <= 8'h10 ;
			data[80070] <= 8'h10 ;
			data[80071] <= 8'h10 ;
			data[80072] <= 8'h10 ;
			data[80073] <= 8'h10 ;
			data[80074] <= 8'h10 ;
			data[80075] <= 8'h10 ;
			data[80076] <= 8'h10 ;
			data[80077] <= 8'h10 ;
			data[80078] <= 8'h10 ;
			data[80079] <= 8'h10 ;
			data[80080] <= 8'h10 ;
			data[80081] <= 8'h10 ;
			data[80082] <= 8'h10 ;
			data[80083] <= 8'h10 ;
			data[80084] <= 8'h10 ;
			data[80085] <= 8'h10 ;
			data[80086] <= 8'h10 ;
			data[80087] <= 8'h10 ;
			data[80088] <= 8'h10 ;
			data[80089] <= 8'h10 ;
			data[80090] <= 8'h10 ;
			data[80091] <= 8'h10 ;
			data[80092] <= 8'h10 ;
			data[80093] <= 8'h10 ;
			data[80094] <= 8'h10 ;
			data[80095] <= 8'h10 ;
			data[80096] <= 8'h10 ;
			data[80097] <= 8'h10 ;
			data[80098] <= 8'h10 ;
			data[80099] <= 8'h10 ;
			data[80100] <= 8'h10 ;
			data[80101] <= 8'h10 ;
			data[80102] <= 8'h10 ;
			data[80103] <= 8'h10 ;
			data[80104] <= 8'h10 ;
			data[80105] <= 8'h10 ;
			data[80106] <= 8'h10 ;
			data[80107] <= 8'h10 ;
			data[80108] <= 8'h10 ;
			data[80109] <= 8'h10 ;
			data[80110] <= 8'h10 ;
			data[80111] <= 8'h10 ;
			data[80112] <= 8'h10 ;
			data[80113] <= 8'h10 ;
			data[80114] <= 8'h10 ;
			data[80115] <= 8'h10 ;
			data[80116] <= 8'h10 ;
			data[80117] <= 8'h10 ;
			data[80118] <= 8'h10 ;
			data[80119] <= 8'h10 ;
			data[80120] <= 8'h10 ;
			data[80121] <= 8'h10 ;
			data[80122] <= 8'h10 ;
			data[80123] <= 8'h10 ;
			data[80124] <= 8'h10 ;
			data[80125] <= 8'h10 ;
			data[80126] <= 8'h10 ;
			data[80127] <= 8'h10 ;
			data[80128] <= 8'h10 ;
			data[80129] <= 8'h10 ;
			data[80130] <= 8'h10 ;
			data[80131] <= 8'h10 ;
			data[80132] <= 8'h10 ;
			data[80133] <= 8'h10 ;
			data[80134] <= 8'h10 ;
			data[80135] <= 8'h10 ;
			data[80136] <= 8'h10 ;
			data[80137] <= 8'h10 ;
			data[80138] <= 8'h10 ;
			data[80139] <= 8'h10 ;
			data[80140] <= 8'h10 ;
			data[80141] <= 8'h10 ;
			data[80142] <= 8'h10 ;
			data[80143] <= 8'h10 ;
			data[80144] <= 8'h10 ;
			data[80145] <= 8'h10 ;
			data[80146] <= 8'h10 ;
			data[80147] <= 8'h10 ;
			data[80148] <= 8'h10 ;
			data[80149] <= 8'h10 ;
			data[80150] <= 8'h10 ;
			data[80151] <= 8'h10 ;
			data[80152] <= 8'h10 ;
			data[80153] <= 8'h10 ;
			data[80154] <= 8'h10 ;
			data[80155] <= 8'h10 ;
			data[80156] <= 8'h10 ;
			data[80157] <= 8'h10 ;
			data[80158] <= 8'h10 ;
			data[80159] <= 8'h10 ;
			data[80160] <= 8'h10 ;
			data[80161] <= 8'h10 ;
			data[80162] <= 8'h10 ;
			data[80163] <= 8'h10 ;
			data[80164] <= 8'h10 ;
			data[80165] <= 8'h10 ;
			data[80166] <= 8'h10 ;
			data[80167] <= 8'h10 ;
			data[80168] <= 8'h10 ;
			data[80169] <= 8'h10 ;
			data[80170] <= 8'h10 ;
			data[80171] <= 8'h10 ;
			data[80172] <= 8'h10 ;
			data[80173] <= 8'h10 ;
			data[80174] <= 8'h10 ;
			data[80175] <= 8'h10 ;
			data[80176] <= 8'h10 ;
			data[80177] <= 8'h10 ;
			data[80178] <= 8'h10 ;
			data[80179] <= 8'h10 ;
			data[80180] <= 8'h10 ;
			data[80181] <= 8'h10 ;
			data[80182] <= 8'h10 ;
			data[80183] <= 8'h10 ;
			data[80184] <= 8'h10 ;
			data[80185] <= 8'h10 ;
			data[80186] <= 8'h10 ;
			data[80187] <= 8'h10 ;
			data[80188] <= 8'h10 ;
			data[80189] <= 8'h10 ;
			data[80190] <= 8'h10 ;
			data[80191] <= 8'h10 ;
			data[80192] <= 8'h10 ;
			data[80193] <= 8'h10 ;
			data[80194] <= 8'h10 ;
			data[80195] <= 8'h10 ;
			data[80196] <= 8'h10 ;
			data[80197] <= 8'h10 ;
			data[80198] <= 8'h10 ;
			data[80199] <= 8'h10 ;
			data[80200] <= 8'h10 ;
			data[80201] <= 8'h10 ;
			data[80202] <= 8'h10 ;
			data[80203] <= 8'h10 ;
			data[80204] <= 8'h10 ;
			data[80205] <= 8'h10 ;
			data[80206] <= 8'h10 ;
			data[80207] <= 8'h10 ;
			data[80208] <= 8'h10 ;
			data[80209] <= 8'h10 ;
			data[80210] <= 8'h10 ;
			data[80211] <= 8'h10 ;
			data[80212] <= 8'h10 ;
			data[80213] <= 8'h10 ;
			data[80214] <= 8'h10 ;
			data[80215] <= 8'h10 ;
			data[80216] <= 8'h10 ;
			data[80217] <= 8'h10 ;
			data[80218] <= 8'h10 ;
			data[80219] <= 8'h10 ;
			data[80220] <= 8'h10 ;
			data[80221] <= 8'h10 ;
			data[80222] <= 8'h10 ;
			data[80223] <= 8'h10 ;
			data[80224] <= 8'h10 ;
			data[80225] <= 8'h10 ;
			data[80226] <= 8'h10 ;
			data[80227] <= 8'h10 ;
			data[80228] <= 8'h10 ;
			data[80229] <= 8'h10 ;
			data[80230] <= 8'h10 ;
			data[80231] <= 8'h10 ;
			data[80232] <= 8'h10 ;
			data[80233] <= 8'h10 ;
			data[80234] <= 8'h10 ;
			data[80235] <= 8'h10 ;
			data[80236] <= 8'h10 ;
			data[80237] <= 8'h10 ;
			data[80238] <= 8'h10 ;
			data[80239] <= 8'h10 ;
			data[80240] <= 8'h10 ;
			data[80241] <= 8'h10 ;
			data[80242] <= 8'h10 ;
			data[80243] <= 8'h10 ;
			data[80244] <= 8'h10 ;
			data[80245] <= 8'h10 ;
			data[80246] <= 8'h10 ;
			data[80247] <= 8'h10 ;
			data[80248] <= 8'h10 ;
			data[80249] <= 8'h10 ;
			data[80250] <= 8'h10 ;
			data[80251] <= 8'h10 ;
			data[80252] <= 8'h10 ;
			data[80253] <= 8'h10 ;
			data[80254] <= 8'h10 ;
			data[80255] <= 8'h10 ;
			data[80256] <= 8'h10 ;
			data[80257] <= 8'h10 ;
			data[80258] <= 8'h10 ;
			data[80259] <= 8'h10 ;
			data[80260] <= 8'h10 ;
			data[80261] <= 8'h10 ;
			data[80262] <= 8'h10 ;
			data[80263] <= 8'h10 ;
			data[80264] <= 8'h10 ;
			data[80265] <= 8'h10 ;
			data[80266] <= 8'h10 ;
			data[80267] <= 8'h10 ;
			data[80268] <= 8'h10 ;
			data[80269] <= 8'h10 ;
			data[80270] <= 8'h10 ;
			data[80271] <= 8'h10 ;
			data[80272] <= 8'h10 ;
			data[80273] <= 8'h10 ;
			data[80274] <= 8'h10 ;
			data[80275] <= 8'h10 ;
			data[80276] <= 8'h10 ;
			data[80277] <= 8'h10 ;
			data[80278] <= 8'h10 ;
			data[80279] <= 8'h10 ;
			data[80280] <= 8'h10 ;
			data[80281] <= 8'h10 ;
			data[80282] <= 8'h10 ;
			data[80283] <= 8'h10 ;
			data[80284] <= 8'h10 ;
			data[80285] <= 8'h10 ;
			data[80286] <= 8'h10 ;
			data[80287] <= 8'h10 ;
			data[80288] <= 8'h10 ;
			data[80289] <= 8'h10 ;
			data[80290] <= 8'h10 ;
			data[80291] <= 8'h10 ;
			data[80292] <= 8'h10 ;
			data[80293] <= 8'h10 ;
			data[80294] <= 8'h10 ;
			data[80295] <= 8'h10 ;
			data[80296] <= 8'h10 ;
			data[80297] <= 8'h10 ;
			data[80298] <= 8'h10 ;
			data[80299] <= 8'h10 ;
			data[80300] <= 8'h10 ;
			data[80301] <= 8'h10 ;
			data[80302] <= 8'h10 ;
			data[80303] <= 8'h10 ;
			data[80304] <= 8'h10 ;
			data[80305] <= 8'h10 ;
			data[80306] <= 8'h10 ;
			data[80307] <= 8'h10 ;
			data[80308] <= 8'h10 ;
			data[80309] <= 8'h10 ;
			data[80310] <= 8'h10 ;
			data[80311] <= 8'h10 ;
			data[80312] <= 8'h10 ;
			data[80313] <= 8'h10 ;
			data[80314] <= 8'h10 ;
			data[80315] <= 8'h10 ;
			data[80316] <= 8'h10 ;
			data[80317] <= 8'h10 ;
			data[80318] <= 8'h10 ;
			data[80319] <= 8'h10 ;
			data[80320] <= 8'h10 ;
			data[80321] <= 8'h10 ;
			data[80322] <= 8'h10 ;
			data[80323] <= 8'h10 ;
			data[80324] <= 8'h10 ;
			data[80325] <= 8'h10 ;
			data[80326] <= 8'h10 ;
			data[80327] <= 8'h10 ;
			data[80328] <= 8'h10 ;
			data[80329] <= 8'h10 ;
			data[80330] <= 8'h10 ;
			data[80331] <= 8'h10 ;
			data[80332] <= 8'h10 ;
			data[80333] <= 8'h10 ;
			data[80334] <= 8'h10 ;
			data[80335] <= 8'h10 ;
			data[80336] <= 8'h10 ;
			data[80337] <= 8'h10 ;
			data[80338] <= 8'h10 ;
			data[80339] <= 8'h10 ;
			data[80340] <= 8'h10 ;
			data[80341] <= 8'h10 ;
			data[80342] <= 8'h10 ;
			data[80343] <= 8'h10 ;
			data[80344] <= 8'h10 ;
			data[80345] <= 8'h10 ;
			data[80346] <= 8'h10 ;
			data[80347] <= 8'h10 ;
			data[80348] <= 8'h10 ;
			data[80349] <= 8'h10 ;
			data[80350] <= 8'h10 ;
			data[80351] <= 8'h10 ;
			data[80352] <= 8'h10 ;
			data[80353] <= 8'h10 ;
			data[80354] <= 8'h10 ;
			data[80355] <= 8'h10 ;
			data[80356] <= 8'h10 ;
			data[80357] <= 8'h10 ;
			data[80358] <= 8'h10 ;
			data[80359] <= 8'h10 ;
			data[80360] <= 8'h10 ;
			data[80361] <= 8'h10 ;
			data[80362] <= 8'h10 ;
			data[80363] <= 8'h10 ;
			data[80364] <= 8'h10 ;
			data[80365] <= 8'h10 ;
			data[80366] <= 8'h10 ;
			data[80367] <= 8'h10 ;
			data[80368] <= 8'h10 ;
			data[80369] <= 8'h10 ;
			data[80370] <= 8'h10 ;
			data[80371] <= 8'h10 ;
			data[80372] <= 8'h10 ;
			data[80373] <= 8'h10 ;
			data[80374] <= 8'h10 ;
			data[80375] <= 8'h10 ;
			data[80376] <= 8'h10 ;
			data[80377] <= 8'h10 ;
			data[80378] <= 8'h10 ;
			data[80379] <= 8'h10 ;
			data[80380] <= 8'h10 ;
			data[80381] <= 8'h10 ;
			data[80382] <= 8'h10 ;
			data[80383] <= 8'h10 ;
			data[80384] <= 8'h10 ;
			data[80385] <= 8'h10 ;
			data[80386] <= 8'h10 ;
			data[80387] <= 8'h10 ;
			data[80388] <= 8'h10 ;
			data[80389] <= 8'h10 ;
			data[80390] <= 8'h10 ;
			data[80391] <= 8'h10 ;
			data[80392] <= 8'h10 ;
			data[80393] <= 8'h10 ;
			data[80394] <= 8'h10 ;
			data[80395] <= 8'h10 ;
			data[80396] <= 8'h10 ;
			data[80397] <= 8'h10 ;
			data[80398] <= 8'h10 ;
			data[80399] <= 8'h10 ;
			data[80400] <= 8'h10 ;
			data[80401] <= 8'h10 ;
			data[80402] <= 8'h10 ;
			data[80403] <= 8'h10 ;
			data[80404] <= 8'h10 ;
			data[80405] <= 8'h10 ;
			data[80406] <= 8'h10 ;
			data[80407] <= 8'h10 ;
			data[80408] <= 8'h10 ;
			data[80409] <= 8'h10 ;
			data[80410] <= 8'h10 ;
			data[80411] <= 8'h10 ;
			data[80412] <= 8'h10 ;
			data[80413] <= 8'h10 ;
			data[80414] <= 8'h10 ;
			data[80415] <= 8'h10 ;
			data[80416] <= 8'h10 ;
			data[80417] <= 8'h10 ;
			data[80418] <= 8'h10 ;
			data[80419] <= 8'h10 ;
			data[80420] <= 8'h10 ;
			data[80421] <= 8'h10 ;
			data[80422] <= 8'h10 ;
			data[80423] <= 8'h10 ;
			data[80424] <= 8'h10 ;
			data[80425] <= 8'h10 ;
			data[80426] <= 8'h10 ;
			data[80427] <= 8'h10 ;
			data[80428] <= 8'h10 ;
			data[80429] <= 8'h10 ;
			data[80430] <= 8'h10 ;
			data[80431] <= 8'h10 ;
			data[80432] <= 8'h10 ;
			data[80433] <= 8'h10 ;
			data[80434] <= 8'h10 ;
			data[80435] <= 8'h10 ;
			data[80436] <= 8'h10 ;
			data[80437] <= 8'h10 ;
			data[80438] <= 8'h10 ;
			data[80439] <= 8'h10 ;
			data[80440] <= 8'h10 ;
			data[80441] <= 8'h10 ;
			data[80442] <= 8'h10 ;
			data[80443] <= 8'h10 ;
			data[80444] <= 8'h10 ;
			data[80445] <= 8'h10 ;
			data[80446] <= 8'h10 ;
			data[80447] <= 8'h10 ;
			data[80448] <= 8'h10 ;
			data[80449] <= 8'h10 ;
			data[80450] <= 8'h10 ;
			data[80451] <= 8'h10 ;
			data[80452] <= 8'h10 ;
			data[80453] <= 8'h10 ;
			data[80454] <= 8'h10 ;
			data[80455] <= 8'h10 ;
			data[80456] <= 8'h10 ;
			data[80457] <= 8'h10 ;
			data[80458] <= 8'h10 ;
			data[80459] <= 8'h10 ;
			data[80460] <= 8'h10 ;
			data[80461] <= 8'h10 ;
			data[80462] <= 8'h10 ;
			data[80463] <= 8'h10 ;
			data[80464] <= 8'h10 ;
			data[80465] <= 8'h10 ;
			data[80466] <= 8'h10 ;
			data[80467] <= 8'h10 ;
			data[80468] <= 8'h10 ;
			data[80469] <= 8'h10 ;
			data[80470] <= 8'h10 ;
			data[80471] <= 8'h10 ;
			data[80472] <= 8'h10 ;
			data[80473] <= 8'h10 ;
			data[80474] <= 8'h10 ;
			data[80475] <= 8'h10 ;
			data[80476] <= 8'h10 ;
			data[80477] <= 8'h10 ;
			data[80478] <= 8'h10 ;
			data[80479] <= 8'h10 ;
			data[80480] <= 8'h10 ;
			data[80481] <= 8'h10 ;
			data[80482] <= 8'h10 ;
			data[80483] <= 8'h10 ;
			data[80484] <= 8'h10 ;
			data[80485] <= 8'h10 ;
			data[80486] <= 8'h10 ;
			data[80487] <= 8'h10 ;
			data[80488] <= 8'h10 ;
			data[80489] <= 8'h10 ;
			data[80490] <= 8'h10 ;
			data[80491] <= 8'h10 ;
			data[80492] <= 8'h10 ;
			data[80493] <= 8'h10 ;
			data[80494] <= 8'h10 ;
			data[80495] <= 8'h10 ;
			data[80496] <= 8'h10 ;
			data[80497] <= 8'h10 ;
			data[80498] <= 8'h10 ;
			data[80499] <= 8'h10 ;
			data[80500] <= 8'h10 ;
			data[80501] <= 8'h10 ;
			data[80502] <= 8'h10 ;
			data[80503] <= 8'h10 ;
			data[80504] <= 8'h10 ;
			data[80505] <= 8'h10 ;
			data[80506] <= 8'h10 ;
			data[80507] <= 8'h10 ;
			data[80508] <= 8'h10 ;
			data[80509] <= 8'h10 ;
			data[80510] <= 8'h10 ;
			data[80511] <= 8'h10 ;
			data[80512] <= 8'h10 ;
			data[80513] <= 8'h10 ;
			data[80514] <= 8'h10 ;
			data[80515] <= 8'h10 ;
			data[80516] <= 8'h10 ;
			data[80517] <= 8'h10 ;
			data[80518] <= 8'h10 ;
			data[80519] <= 8'h10 ;
			data[80520] <= 8'h10 ;
			data[80521] <= 8'h10 ;
			data[80522] <= 8'h10 ;
			data[80523] <= 8'h10 ;
			data[80524] <= 8'h10 ;
			data[80525] <= 8'h10 ;
			data[80526] <= 8'h10 ;
			data[80527] <= 8'h10 ;
			data[80528] <= 8'h10 ;
			data[80529] <= 8'h10 ;
			data[80530] <= 8'h10 ;
			data[80531] <= 8'h10 ;
			data[80532] <= 8'h10 ;
			data[80533] <= 8'h10 ;
			data[80534] <= 8'h10 ;
			data[80535] <= 8'h10 ;
			data[80536] <= 8'h10 ;
			data[80537] <= 8'h10 ;
			data[80538] <= 8'h10 ;
			data[80539] <= 8'h10 ;
			data[80540] <= 8'h10 ;
			data[80541] <= 8'h10 ;
			data[80542] <= 8'h10 ;
			data[80543] <= 8'h10 ;
			data[80544] <= 8'h10 ;
			data[80545] <= 8'h10 ;
			data[80546] <= 8'h10 ;
			data[80547] <= 8'h10 ;
			data[80548] <= 8'h10 ;
			data[80549] <= 8'h10 ;
			data[80550] <= 8'h10 ;
			data[80551] <= 8'h10 ;
			data[80552] <= 8'h10 ;
			data[80553] <= 8'h10 ;
			data[80554] <= 8'h10 ;
			data[80555] <= 8'h10 ;
			data[80556] <= 8'h10 ;
			data[80557] <= 8'h10 ;
			data[80558] <= 8'h10 ;
			data[80559] <= 8'h10 ;
			data[80560] <= 8'h10 ;
			data[80561] <= 8'h10 ;
			data[80562] <= 8'h10 ;
			data[80563] <= 8'h10 ;
			data[80564] <= 8'h10 ;
			data[80565] <= 8'h10 ;
			data[80566] <= 8'h10 ;
			data[80567] <= 8'h10 ;
			data[80568] <= 8'h10 ;
			data[80569] <= 8'h10 ;
			data[80570] <= 8'h10 ;
			data[80571] <= 8'h10 ;
			data[80572] <= 8'h10 ;
			data[80573] <= 8'h10 ;
			data[80574] <= 8'h10 ;
			data[80575] <= 8'h10 ;
			data[80576] <= 8'h10 ;
			data[80577] <= 8'h10 ;
			data[80578] <= 8'h10 ;
			data[80579] <= 8'h10 ;
			data[80580] <= 8'h10 ;
			data[80581] <= 8'h10 ;
			data[80582] <= 8'h10 ;
			data[80583] <= 8'h10 ;
			data[80584] <= 8'h10 ;
			data[80585] <= 8'h10 ;
			data[80586] <= 8'h10 ;
			data[80587] <= 8'h10 ;
			data[80588] <= 8'h10 ;
			data[80589] <= 8'h10 ;
			data[80590] <= 8'h10 ;
			data[80591] <= 8'h10 ;
			data[80592] <= 8'h10 ;
			data[80593] <= 8'h10 ;
			data[80594] <= 8'h10 ;
			data[80595] <= 8'h10 ;
			data[80596] <= 8'h10 ;
			data[80597] <= 8'h10 ;
			data[80598] <= 8'h10 ;
			data[80599] <= 8'h10 ;
			data[80600] <= 8'h10 ;
			data[80601] <= 8'h10 ;
			data[80602] <= 8'h10 ;
			data[80603] <= 8'h10 ;
			data[80604] <= 8'h10 ;
			data[80605] <= 8'h10 ;
			data[80606] <= 8'h10 ;
			data[80607] <= 8'h10 ;
			data[80608] <= 8'h10 ;
			data[80609] <= 8'h10 ;
			data[80610] <= 8'h10 ;
			data[80611] <= 8'h10 ;
			data[80612] <= 8'h10 ;
			data[80613] <= 8'h10 ;
			data[80614] <= 8'h10 ;
			data[80615] <= 8'h10 ;
			data[80616] <= 8'h10 ;
			data[80617] <= 8'h10 ;
			data[80618] <= 8'h10 ;
			data[80619] <= 8'h10 ;
			data[80620] <= 8'h10 ;
			data[80621] <= 8'h10 ;
			data[80622] <= 8'h10 ;
			data[80623] <= 8'h10 ;
			data[80624] <= 8'h10 ;
			data[80625] <= 8'h10 ;
			data[80626] <= 8'h10 ;
			data[80627] <= 8'h10 ;
			data[80628] <= 8'h10 ;
			data[80629] <= 8'h10 ;
			data[80630] <= 8'h10 ;
			data[80631] <= 8'h10 ;
			data[80632] <= 8'h10 ;
			data[80633] <= 8'h10 ;
			data[80634] <= 8'h10 ;
			data[80635] <= 8'h10 ;
			data[80636] <= 8'h10 ;
			data[80637] <= 8'h10 ;
			data[80638] <= 8'h10 ;
			data[80639] <= 8'h10 ;
			data[80640] <= 8'h10 ;
			data[80641] <= 8'h10 ;
			data[80642] <= 8'h10 ;
			data[80643] <= 8'h10 ;
			data[80644] <= 8'h10 ;
			data[80645] <= 8'h10 ;
			data[80646] <= 8'h10 ;
			data[80647] <= 8'h10 ;
			data[80648] <= 8'h10 ;
			data[80649] <= 8'h10 ;
			data[80650] <= 8'h10 ;
			data[80651] <= 8'h10 ;
			data[80652] <= 8'h10 ;
			data[80653] <= 8'h10 ;
			data[80654] <= 8'h10 ;
			data[80655] <= 8'h10 ;
			data[80656] <= 8'h10 ;
			data[80657] <= 8'h10 ;
			data[80658] <= 8'h10 ;
			data[80659] <= 8'h10 ;
			data[80660] <= 8'h10 ;
			data[80661] <= 8'h10 ;
			data[80662] <= 8'h10 ;
			data[80663] <= 8'h10 ;
			data[80664] <= 8'h10 ;
			data[80665] <= 8'h10 ;
			data[80666] <= 8'h10 ;
			data[80667] <= 8'h10 ;
			data[80668] <= 8'h10 ;
			data[80669] <= 8'h10 ;
			data[80670] <= 8'h10 ;
			data[80671] <= 8'h10 ;
			data[80672] <= 8'h10 ;
			data[80673] <= 8'h10 ;
			data[80674] <= 8'h10 ;
			data[80675] <= 8'h10 ;
			data[80676] <= 8'h10 ;
			data[80677] <= 8'h10 ;
			data[80678] <= 8'h10 ;
			data[80679] <= 8'h10 ;
			data[80680] <= 8'h10 ;
			data[80681] <= 8'h10 ;
			data[80682] <= 8'h10 ;
			data[80683] <= 8'h10 ;
			data[80684] <= 8'h10 ;
			data[80685] <= 8'h10 ;
			data[80686] <= 8'h10 ;
			data[80687] <= 8'h10 ;
			data[80688] <= 8'h10 ;
			data[80689] <= 8'h10 ;
			data[80690] <= 8'h10 ;
			data[80691] <= 8'h10 ;
			data[80692] <= 8'h10 ;
			data[80693] <= 8'h10 ;
			data[80694] <= 8'h10 ;
			data[80695] <= 8'h10 ;
			data[80696] <= 8'h10 ;
			data[80697] <= 8'h10 ;
			data[80698] <= 8'h10 ;
			data[80699] <= 8'h10 ;
			data[80700] <= 8'h10 ;
			data[80701] <= 8'h10 ;
			data[80702] <= 8'h10 ;
			data[80703] <= 8'h10 ;
			data[80704] <= 8'h10 ;
			data[80705] <= 8'h10 ;
			data[80706] <= 8'h10 ;
			data[80707] <= 8'h10 ;
			data[80708] <= 8'h10 ;
			data[80709] <= 8'h10 ;
			data[80710] <= 8'h10 ;
			data[80711] <= 8'h10 ;
			data[80712] <= 8'h10 ;
			data[80713] <= 8'h10 ;
			data[80714] <= 8'h10 ;
			data[80715] <= 8'h10 ;
			data[80716] <= 8'h10 ;
			data[80717] <= 8'h10 ;
			data[80718] <= 8'h10 ;
			data[80719] <= 8'h10 ;
			data[80720] <= 8'h10 ;
			data[80721] <= 8'h10 ;
			data[80722] <= 8'h10 ;
			data[80723] <= 8'h10 ;
			data[80724] <= 8'h10 ;
			data[80725] <= 8'h10 ;
			data[80726] <= 8'h10 ;
			data[80727] <= 8'h10 ;
			data[80728] <= 8'h10 ;
			data[80729] <= 8'h10 ;
			data[80730] <= 8'h10 ;
			data[80731] <= 8'h10 ;
			data[80732] <= 8'h10 ;
			data[80733] <= 8'h10 ;
			data[80734] <= 8'h10 ;
			data[80735] <= 8'h10 ;
			data[80736] <= 8'h10 ;
			data[80737] <= 8'h10 ;
			data[80738] <= 8'h10 ;
			data[80739] <= 8'h10 ;
			data[80740] <= 8'h10 ;
			data[80741] <= 8'h10 ;
			data[80742] <= 8'h10 ;
			data[80743] <= 8'h10 ;
			data[80744] <= 8'h10 ;
			data[80745] <= 8'h10 ;
			data[80746] <= 8'h10 ;
			data[80747] <= 8'h10 ;
			data[80748] <= 8'h10 ;
			data[80749] <= 8'h10 ;
			data[80750] <= 8'h10 ;
			data[80751] <= 8'h10 ;
			data[80752] <= 8'h10 ;
			data[80753] <= 8'h10 ;
			data[80754] <= 8'h10 ;
			data[80755] <= 8'h10 ;
			data[80756] <= 8'h10 ;
			data[80757] <= 8'h10 ;
			data[80758] <= 8'h10 ;
			data[80759] <= 8'h10 ;
			data[80760] <= 8'h10 ;
			data[80761] <= 8'h10 ;
			data[80762] <= 8'h10 ;
			data[80763] <= 8'h10 ;
			data[80764] <= 8'h10 ;
			data[80765] <= 8'h10 ;
			data[80766] <= 8'h10 ;
			data[80767] <= 8'h10 ;
			data[80768] <= 8'h10 ;
			data[80769] <= 8'h10 ;
			data[80770] <= 8'h10 ;
			data[80771] <= 8'h10 ;
			data[80772] <= 8'h10 ;
			data[80773] <= 8'h10 ;
			data[80774] <= 8'h10 ;
			data[80775] <= 8'h10 ;
			data[80776] <= 8'h10 ;
			data[80777] <= 8'h10 ;
			data[80778] <= 8'h10 ;
			data[80779] <= 8'h10 ;
			data[80780] <= 8'h10 ;
			data[80781] <= 8'h10 ;
			data[80782] <= 8'h10 ;
			data[80783] <= 8'h10 ;
			data[80784] <= 8'h10 ;
			data[80785] <= 8'h10 ;
			data[80786] <= 8'h10 ;
			data[80787] <= 8'h10 ;
			data[80788] <= 8'h10 ;
			data[80789] <= 8'h10 ;
			data[80790] <= 8'h10 ;
			data[80791] <= 8'h10 ;
			data[80792] <= 8'h10 ;
			data[80793] <= 8'h10 ;
			data[80794] <= 8'h10 ;
			data[80795] <= 8'h10 ;
			data[80796] <= 8'h10 ;
			data[80797] <= 8'h10 ;
			data[80798] <= 8'h10 ;
			data[80799] <= 8'h10 ;
			data[80800] <= 8'h10 ;
			data[80801] <= 8'h10 ;
			data[80802] <= 8'h10 ;
			data[80803] <= 8'h10 ;
			data[80804] <= 8'h10 ;
			data[80805] <= 8'h10 ;
			data[80806] <= 8'h10 ;
			data[80807] <= 8'h10 ;
			data[80808] <= 8'h10 ;
			data[80809] <= 8'h10 ;
			data[80810] <= 8'h10 ;
			data[80811] <= 8'h10 ;
			data[80812] <= 8'h10 ;
			data[80813] <= 8'h10 ;
			data[80814] <= 8'h10 ;
			data[80815] <= 8'h10 ;
			data[80816] <= 8'h10 ;
			data[80817] <= 8'h10 ;
			data[80818] <= 8'h10 ;
			data[80819] <= 8'h10 ;
			data[80820] <= 8'h10 ;
			data[80821] <= 8'h10 ;
			data[80822] <= 8'h10 ;
			data[80823] <= 8'h10 ;
			data[80824] <= 8'h10 ;
			data[80825] <= 8'h10 ;
			data[80826] <= 8'h10 ;
			data[80827] <= 8'h10 ;
			data[80828] <= 8'h10 ;
			data[80829] <= 8'h10 ;
			data[80830] <= 8'h10 ;
			data[80831] <= 8'h10 ;
			data[80832] <= 8'h10 ;
			data[80833] <= 8'h10 ;
			data[80834] <= 8'h10 ;
			data[80835] <= 8'h10 ;
			data[80836] <= 8'h10 ;
			data[80837] <= 8'h10 ;
			data[80838] <= 8'h10 ;
			data[80839] <= 8'h10 ;
			data[80840] <= 8'h10 ;
			data[80841] <= 8'h10 ;
			data[80842] <= 8'h10 ;
			data[80843] <= 8'h10 ;
			data[80844] <= 8'h10 ;
			data[80845] <= 8'h10 ;
			data[80846] <= 8'h10 ;
			data[80847] <= 8'h10 ;
			data[80848] <= 8'h10 ;
			data[80849] <= 8'h10 ;
			data[80850] <= 8'h10 ;
			data[80851] <= 8'h10 ;
			data[80852] <= 8'h10 ;
			data[80853] <= 8'h10 ;
			data[80854] <= 8'h10 ;
			data[80855] <= 8'h10 ;
			data[80856] <= 8'h10 ;
			data[80857] <= 8'h10 ;
			data[80858] <= 8'h10 ;
			data[80859] <= 8'h10 ;
			data[80860] <= 8'h10 ;
			data[80861] <= 8'h10 ;
			data[80862] <= 8'h10 ;
			data[80863] <= 8'h10 ;
			data[80864] <= 8'h10 ;
			data[80865] <= 8'h10 ;
			data[80866] <= 8'h10 ;
			data[80867] <= 8'h10 ;
			data[80868] <= 8'h10 ;
			data[80869] <= 8'h10 ;
			data[80870] <= 8'h10 ;
			data[80871] <= 8'h10 ;
			data[80872] <= 8'h10 ;
			data[80873] <= 8'h10 ;
			data[80874] <= 8'h10 ;
			data[80875] <= 8'h10 ;
			data[80876] <= 8'h10 ;
			data[80877] <= 8'h10 ;
			data[80878] <= 8'h10 ;
			data[80879] <= 8'h10 ;
			data[80880] <= 8'h10 ;
			data[80881] <= 8'h10 ;
			data[80882] <= 8'h10 ;
			data[80883] <= 8'h10 ;
			data[80884] <= 8'h10 ;
			data[80885] <= 8'h10 ;
			data[80886] <= 8'h10 ;
			data[80887] <= 8'h10 ;
			data[80888] <= 8'h10 ;
			data[80889] <= 8'h10 ;
			data[80890] <= 8'h10 ;
			data[80891] <= 8'h10 ;
			data[80892] <= 8'h10 ;
			data[80893] <= 8'h10 ;
			data[80894] <= 8'h10 ;
			data[80895] <= 8'h10 ;
			data[80896] <= 8'h10 ;
			data[80897] <= 8'h10 ;
			data[80898] <= 8'h10 ;
			data[80899] <= 8'h10 ;
			data[80900] <= 8'h10 ;
			data[80901] <= 8'h10 ;
			data[80902] <= 8'h10 ;
			data[80903] <= 8'h10 ;
			data[80904] <= 8'h10 ;
			data[80905] <= 8'h10 ;
			data[80906] <= 8'h10 ;
			data[80907] <= 8'h10 ;
			data[80908] <= 8'h10 ;
			data[80909] <= 8'h10 ;
			data[80910] <= 8'h10 ;
			data[80911] <= 8'h10 ;
			data[80912] <= 8'h10 ;
			data[80913] <= 8'h10 ;
			data[80914] <= 8'h10 ;
			data[80915] <= 8'h10 ;
			data[80916] <= 8'h10 ;
			data[80917] <= 8'h10 ;
			data[80918] <= 8'h10 ;
			data[80919] <= 8'h10 ;
			data[80920] <= 8'h10 ;
			data[80921] <= 8'h10 ;
			data[80922] <= 8'h10 ;
			data[80923] <= 8'h10 ;
			data[80924] <= 8'h10 ;
			data[80925] <= 8'h10 ;
			data[80926] <= 8'h10 ;
			data[80927] <= 8'h10 ;
			data[80928] <= 8'h10 ;
			data[80929] <= 8'h10 ;
			data[80930] <= 8'h10 ;
			data[80931] <= 8'h10 ;
			data[80932] <= 8'h10 ;
			data[80933] <= 8'h10 ;
			data[80934] <= 8'h10 ;
			data[80935] <= 8'h10 ;
			data[80936] <= 8'h10 ;
			data[80937] <= 8'h10 ;
			data[80938] <= 8'h10 ;
			data[80939] <= 8'h10 ;
			data[80940] <= 8'h10 ;
			data[80941] <= 8'h10 ;
			data[80942] <= 8'h10 ;
			data[80943] <= 8'h10 ;
			data[80944] <= 8'h10 ;
			data[80945] <= 8'h10 ;
			data[80946] <= 8'h10 ;
			data[80947] <= 8'h10 ;
			data[80948] <= 8'h10 ;
			data[80949] <= 8'h10 ;
			data[80950] <= 8'h10 ;
			data[80951] <= 8'h10 ;
			data[80952] <= 8'h10 ;
			data[80953] <= 8'h10 ;
			data[80954] <= 8'h10 ;
			data[80955] <= 8'h10 ;
			data[80956] <= 8'h10 ;
			data[80957] <= 8'h10 ;
			data[80958] <= 8'h10 ;
			data[80959] <= 8'h10 ;
			data[80960] <= 8'h10 ;
			data[80961] <= 8'h10 ;
			data[80962] <= 8'h10 ;
			data[80963] <= 8'h10 ;
			data[80964] <= 8'h10 ;
			data[80965] <= 8'h10 ;
			data[80966] <= 8'h10 ;
			data[80967] <= 8'h10 ;
			data[80968] <= 8'h10 ;
			data[80969] <= 8'h10 ;
			data[80970] <= 8'h10 ;
			data[80971] <= 8'h10 ;
			data[80972] <= 8'h10 ;
			data[80973] <= 8'h10 ;
			data[80974] <= 8'h10 ;
			data[80975] <= 8'h10 ;
			data[80976] <= 8'h10 ;
			data[80977] <= 8'h10 ;
			data[80978] <= 8'h10 ;
			data[80979] <= 8'h10 ;
			data[80980] <= 8'h10 ;
			data[80981] <= 8'h10 ;
			data[80982] <= 8'h10 ;
			data[80983] <= 8'h10 ;
			data[80984] <= 8'h10 ;
			data[80985] <= 8'h10 ;
			data[80986] <= 8'h10 ;
			data[80987] <= 8'h10 ;
			data[80988] <= 8'h10 ;
			data[80989] <= 8'h10 ;
			data[80990] <= 8'h10 ;
			data[80991] <= 8'h10 ;
			data[80992] <= 8'h10 ;
			data[80993] <= 8'h10 ;
			data[80994] <= 8'h10 ;
			data[80995] <= 8'h10 ;
			data[80996] <= 8'h10 ;
			data[80997] <= 8'h10 ;
			data[80998] <= 8'h10 ;
			data[80999] <= 8'h10 ;
			data[81000] <= 8'h10 ;
			data[81001] <= 8'h10 ;
			data[81002] <= 8'h10 ;
			data[81003] <= 8'h10 ;
			data[81004] <= 8'h10 ;
			data[81005] <= 8'h10 ;
			data[81006] <= 8'h10 ;
			data[81007] <= 8'h10 ;
			data[81008] <= 8'h10 ;
			data[81009] <= 8'h10 ;
			data[81010] <= 8'h10 ;
			data[81011] <= 8'h10 ;
			data[81012] <= 8'h10 ;
			data[81013] <= 8'h10 ;
			data[81014] <= 8'h10 ;
			data[81015] <= 8'h10 ;
			data[81016] <= 8'h10 ;
			data[81017] <= 8'h10 ;
			data[81018] <= 8'h10 ;
			data[81019] <= 8'h10 ;
			data[81020] <= 8'h10 ;
			data[81021] <= 8'h10 ;
			data[81022] <= 8'h10 ;
			data[81023] <= 8'h10 ;
			data[81024] <= 8'h10 ;
			data[81025] <= 8'h10 ;
			data[81026] <= 8'h10 ;
			data[81027] <= 8'h10 ;
			data[81028] <= 8'h10 ;
			data[81029] <= 8'h10 ;
			data[81030] <= 8'h10 ;
			data[81031] <= 8'h10 ;
			data[81032] <= 8'h10 ;
			data[81033] <= 8'h10 ;
			data[81034] <= 8'h10 ;
			data[81035] <= 8'h10 ;
			data[81036] <= 8'h10 ;
			data[81037] <= 8'h10 ;
			data[81038] <= 8'h10 ;
			data[81039] <= 8'h10 ;
			data[81040] <= 8'h10 ;
			data[81041] <= 8'h10 ;
			data[81042] <= 8'h10 ;
			data[81043] <= 8'h10 ;
			data[81044] <= 8'h10 ;
			data[81045] <= 8'h10 ;
			data[81046] <= 8'h10 ;
			data[81047] <= 8'h10 ;
			data[81048] <= 8'h10 ;
			data[81049] <= 8'h10 ;
			data[81050] <= 8'h10 ;
			data[81051] <= 8'h10 ;
			data[81052] <= 8'h10 ;
			data[81053] <= 8'h10 ;
			data[81054] <= 8'h10 ;
			data[81055] <= 8'h10 ;
			data[81056] <= 8'h10 ;
			data[81057] <= 8'h10 ;
			data[81058] <= 8'h10 ;
			data[81059] <= 8'h10 ;
			data[81060] <= 8'h10 ;
			data[81061] <= 8'h10 ;
			data[81062] <= 8'h10 ;
			data[81063] <= 8'h10 ;
			data[81064] <= 8'h10 ;
			data[81065] <= 8'h10 ;
			data[81066] <= 8'h10 ;
			data[81067] <= 8'h10 ;
			data[81068] <= 8'h10 ;
			data[81069] <= 8'h10 ;
			data[81070] <= 8'h10 ;
			data[81071] <= 8'h10 ;
			data[81072] <= 8'h10 ;
			data[81073] <= 8'h10 ;
			data[81074] <= 8'h10 ;
			data[81075] <= 8'h10 ;
			data[81076] <= 8'h10 ;
			data[81077] <= 8'h10 ;
			data[81078] <= 8'h10 ;
			data[81079] <= 8'h10 ;
			data[81080] <= 8'h10 ;
			data[81081] <= 8'h10 ;
			data[81082] <= 8'h10 ;
			data[81083] <= 8'h10 ;
			data[81084] <= 8'h10 ;
			data[81085] <= 8'h10 ;
			data[81086] <= 8'h10 ;
			data[81087] <= 8'h10 ;
			data[81088] <= 8'h10 ;
			data[81089] <= 8'h10 ;
			data[81090] <= 8'h10 ;
			data[81091] <= 8'h10 ;
			data[81092] <= 8'h10 ;
			data[81093] <= 8'h10 ;
			data[81094] <= 8'h10 ;
			data[81095] <= 8'h10 ;
			data[81096] <= 8'h10 ;
			data[81097] <= 8'h10 ;
			data[81098] <= 8'h10 ;
			data[81099] <= 8'h10 ;
			data[81100] <= 8'h10 ;
			data[81101] <= 8'h10 ;
			data[81102] <= 8'h10 ;
			data[81103] <= 8'h10 ;
			data[81104] <= 8'h10 ;
			data[81105] <= 8'h10 ;
			data[81106] <= 8'h10 ;
			data[81107] <= 8'h10 ;
			data[81108] <= 8'h10 ;
			data[81109] <= 8'h10 ;
			data[81110] <= 8'h10 ;
			data[81111] <= 8'h10 ;
			data[81112] <= 8'h10 ;
			data[81113] <= 8'h10 ;
			data[81114] <= 8'h10 ;
			data[81115] <= 8'h10 ;
			data[81116] <= 8'h10 ;
			data[81117] <= 8'h10 ;
			data[81118] <= 8'h10 ;
			data[81119] <= 8'h10 ;
			data[81120] <= 8'h10 ;
			data[81121] <= 8'h10 ;
			data[81122] <= 8'h10 ;
			data[81123] <= 8'h10 ;
			data[81124] <= 8'h10 ;
			data[81125] <= 8'h10 ;
			data[81126] <= 8'h10 ;
			data[81127] <= 8'h10 ;
			data[81128] <= 8'h10 ;
			data[81129] <= 8'h10 ;
			data[81130] <= 8'h10 ;
			data[81131] <= 8'h10 ;
			data[81132] <= 8'h10 ;
			data[81133] <= 8'h10 ;
			data[81134] <= 8'h10 ;
			data[81135] <= 8'h10 ;
			data[81136] <= 8'h10 ;
			data[81137] <= 8'h10 ;
			data[81138] <= 8'h10 ;
			data[81139] <= 8'h10 ;
			data[81140] <= 8'h10 ;
			data[81141] <= 8'h10 ;
			data[81142] <= 8'h10 ;
			data[81143] <= 8'h10 ;
			data[81144] <= 8'h10 ;
			data[81145] <= 8'h10 ;
			data[81146] <= 8'h10 ;
			data[81147] <= 8'h10 ;
			data[81148] <= 8'h10 ;
			data[81149] <= 8'h10 ;
			data[81150] <= 8'h10 ;
			data[81151] <= 8'h10 ;
			data[81152] <= 8'h10 ;
			data[81153] <= 8'h10 ;
			data[81154] <= 8'h10 ;
			data[81155] <= 8'h10 ;
			data[81156] <= 8'h10 ;
			data[81157] <= 8'h10 ;
			data[81158] <= 8'h10 ;
			data[81159] <= 8'h10 ;
			data[81160] <= 8'h10 ;
			data[81161] <= 8'h10 ;
			data[81162] <= 8'h10 ;
			data[81163] <= 8'h10 ;
			data[81164] <= 8'h10 ;
			data[81165] <= 8'h10 ;
			data[81166] <= 8'h10 ;
			data[81167] <= 8'h10 ;
			data[81168] <= 8'h10 ;
			data[81169] <= 8'h10 ;
			data[81170] <= 8'h10 ;
			data[81171] <= 8'h10 ;
			data[81172] <= 8'h10 ;
			data[81173] <= 8'h10 ;
			data[81174] <= 8'h10 ;
			data[81175] <= 8'h10 ;
			data[81176] <= 8'h10 ;
			data[81177] <= 8'h10 ;
			data[81178] <= 8'h10 ;
			data[81179] <= 8'h10 ;
			data[81180] <= 8'h10 ;
			data[81181] <= 8'h10 ;
			data[81182] <= 8'h10 ;
			data[81183] <= 8'h10 ;
			data[81184] <= 8'h10 ;
			data[81185] <= 8'h10 ;
			data[81186] <= 8'h10 ;
			data[81187] <= 8'h10 ;
			data[81188] <= 8'h10 ;
			data[81189] <= 8'h10 ;
			data[81190] <= 8'h10 ;
			data[81191] <= 8'h10 ;
			data[81192] <= 8'h10 ;
			data[81193] <= 8'h10 ;
			data[81194] <= 8'h10 ;
			data[81195] <= 8'h10 ;
			data[81196] <= 8'h10 ;
			data[81197] <= 8'h10 ;
			data[81198] <= 8'h10 ;
			data[81199] <= 8'h10 ;
			data[81200] <= 8'h10 ;
			data[81201] <= 8'h10 ;
			data[81202] <= 8'h10 ;
			data[81203] <= 8'h10 ;
			data[81204] <= 8'h10 ;
			data[81205] <= 8'h10 ;
			data[81206] <= 8'h10 ;
			data[81207] <= 8'h10 ;
			data[81208] <= 8'h10 ;
			data[81209] <= 8'h10 ;
			data[81210] <= 8'h10 ;
			data[81211] <= 8'h10 ;
			data[81212] <= 8'h10 ;
			data[81213] <= 8'h10 ;
			data[81214] <= 8'h10 ;
			data[81215] <= 8'h10 ;
			data[81216] <= 8'h10 ;
			data[81217] <= 8'h10 ;
			data[81218] <= 8'h10 ;
			data[81219] <= 8'h10 ;
			data[81220] <= 8'h10 ;
			data[81221] <= 8'h10 ;
			data[81222] <= 8'h10 ;
			data[81223] <= 8'h10 ;
			data[81224] <= 8'h10 ;
			data[81225] <= 8'h10 ;
			data[81226] <= 8'h10 ;
			data[81227] <= 8'h10 ;
			data[81228] <= 8'h10 ;
			data[81229] <= 8'h10 ;
			data[81230] <= 8'h10 ;
			data[81231] <= 8'h10 ;
			data[81232] <= 8'h10 ;
			data[81233] <= 8'h10 ;
			data[81234] <= 8'h10 ;
			data[81235] <= 8'h10 ;
			data[81236] <= 8'h10 ;
			data[81237] <= 8'h10 ;
			data[81238] <= 8'h10 ;
			data[81239] <= 8'h10 ;
			data[81240] <= 8'h10 ;
			data[81241] <= 8'h10 ;
			data[81242] <= 8'h10 ;
			data[81243] <= 8'h10 ;
			data[81244] <= 8'h10 ;
			data[81245] <= 8'h10 ;
			data[81246] <= 8'h10 ;
			data[81247] <= 8'h10 ;
			data[81248] <= 8'h10 ;
			data[81249] <= 8'h10 ;
			data[81250] <= 8'h10 ;
			data[81251] <= 8'h10 ;
			data[81252] <= 8'h10 ;
			data[81253] <= 8'h10 ;
			data[81254] <= 8'h10 ;
			data[81255] <= 8'h10 ;
			data[81256] <= 8'h10 ;
			data[81257] <= 8'h10 ;
			data[81258] <= 8'h10 ;
			data[81259] <= 8'h10 ;
			data[81260] <= 8'h10 ;
			data[81261] <= 8'h10 ;
			data[81262] <= 8'h10 ;
			data[81263] <= 8'h10 ;
			data[81264] <= 8'h10 ;
			data[81265] <= 8'h10 ;
			data[81266] <= 8'h10 ;
			data[81267] <= 8'h10 ;
			data[81268] <= 8'h10 ;
			data[81269] <= 8'h10 ;
			data[81270] <= 8'h10 ;
			data[81271] <= 8'h10 ;
			data[81272] <= 8'h10 ;
			data[81273] <= 8'h10 ;
			data[81274] <= 8'h10 ;
			data[81275] <= 8'h10 ;
			data[81276] <= 8'h10 ;
			data[81277] <= 8'h10 ;
			data[81278] <= 8'h10 ;
			data[81279] <= 8'h10 ;
			data[81280] <= 8'h10 ;
			data[81281] <= 8'h10 ;
			data[81282] <= 8'h10 ;
			data[81283] <= 8'h10 ;
			data[81284] <= 8'h10 ;
			data[81285] <= 8'h10 ;
			data[81286] <= 8'h10 ;
			data[81287] <= 8'h10 ;
			data[81288] <= 8'h10 ;
			data[81289] <= 8'h10 ;
			data[81290] <= 8'h10 ;
			data[81291] <= 8'h10 ;
			data[81292] <= 8'h10 ;
			data[81293] <= 8'h10 ;
			data[81294] <= 8'h10 ;
			data[81295] <= 8'h10 ;
			data[81296] <= 8'h10 ;
			data[81297] <= 8'h10 ;
			data[81298] <= 8'h10 ;
			data[81299] <= 8'h10 ;
			data[81300] <= 8'h10 ;
			data[81301] <= 8'h10 ;
			data[81302] <= 8'h10 ;
			data[81303] <= 8'h10 ;
			data[81304] <= 8'h10 ;
			data[81305] <= 8'h10 ;
			data[81306] <= 8'h10 ;
			data[81307] <= 8'h10 ;
			data[81308] <= 8'h10 ;
			data[81309] <= 8'h10 ;
			data[81310] <= 8'h10 ;
			data[81311] <= 8'h10 ;
			data[81312] <= 8'h10 ;
			data[81313] <= 8'h10 ;
			data[81314] <= 8'h10 ;
			data[81315] <= 8'h10 ;
			data[81316] <= 8'h10 ;
			data[81317] <= 8'h10 ;
			data[81318] <= 8'h10 ;
			data[81319] <= 8'h10 ;
			data[81320] <= 8'h10 ;
			data[81321] <= 8'h10 ;
			data[81322] <= 8'h10 ;
			data[81323] <= 8'h10 ;
			data[81324] <= 8'h10 ;
			data[81325] <= 8'h10 ;
			data[81326] <= 8'h10 ;
			data[81327] <= 8'h10 ;
			data[81328] <= 8'h10 ;
			data[81329] <= 8'h10 ;
			data[81330] <= 8'h10 ;
			data[81331] <= 8'h10 ;
			data[81332] <= 8'h10 ;
			data[81333] <= 8'h10 ;
			data[81334] <= 8'h10 ;
			data[81335] <= 8'h10 ;
			data[81336] <= 8'h10 ;
			data[81337] <= 8'h10 ;
			data[81338] <= 8'h10 ;
			data[81339] <= 8'h10 ;
			data[81340] <= 8'h10 ;
			data[81341] <= 8'h10 ;
			data[81342] <= 8'h10 ;
			data[81343] <= 8'h10 ;
			data[81344] <= 8'h10 ;
			data[81345] <= 8'h10 ;
			data[81346] <= 8'h10 ;
			data[81347] <= 8'h10 ;
			data[81348] <= 8'h10 ;
			data[81349] <= 8'h10 ;
			data[81350] <= 8'h10 ;
			data[81351] <= 8'h10 ;
			data[81352] <= 8'h10 ;
			data[81353] <= 8'h10 ;
			data[81354] <= 8'h10 ;
			data[81355] <= 8'h10 ;
			data[81356] <= 8'h10 ;
			data[81357] <= 8'h10 ;
			data[81358] <= 8'h10 ;
			data[81359] <= 8'h10 ;
			data[81360] <= 8'h10 ;
			data[81361] <= 8'h10 ;
			data[81362] <= 8'h10 ;
			data[81363] <= 8'h10 ;
			data[81364] <= 8'h10 ;
			data[81365] <= 8'h10 ;
			data[81366] <= 8'h10 ;
			data[81367] <= 8'h10 ;
			data[81368] <= 8'h10 ;
			data[81369] <= 8'h10 ;
			data[81370] <= 8'h10 ;
			data[81371] <= 8'h10 ;
			data[81372] <= 8'h10 ;
			data[81373] <= 8'h10 ;
			data[81374] <= 8'h10 ;
			data[81375] <= 8'h10 ;
			data[81376] <= 8'h10 ;
			data[81377] <= 8'h10 ;
			data[81378] <= 8'h10 ;
			data[81379] <= 8'h10 ;
			data[81380] <= 8'h10 ;
			data[81381] <= 8'h10 ;
			data[81382] <= 8'h10 ;
			data[81383] <= 8'h10 ;
			data[81384] <= 8'h10 ;
			data[81385] <= 8'h10 ;
			data[81386] <= 8'h10 ;
			data[81387] <= 8'h10 ;
			data[81388] <= 8'h10 ;
			data[81389] <= 8'h10 ;
			data[81390] <= 8'h10 ;
			data[81391] <= 8'h10 ;
			data[81392] <= 8'h10 ;
			data[81393] <= 8'h10 ;
			data[81394] <= 8'h10 ;
			data[81395] <= 8'h10 ;
			data[81396] <= 8'h10 ;
			data[81397] <= 8'h10 ;
			data[81398] <= 8'h10 ;
			data[81399] <= 8'h10 ;
			data[81400] <= 8'h10 ;
			data[81401] <= 8'h10 ;
			data[81402] <= 8'h10 ;
			data[81403] <= 8'h10 ;
			data[81404] <= 8'h10 ;
			data[81405] <= 8'h10 ;
			data[81406] <= 8'h10 ;
			data[81407] <= 8'h10 ;
			data[81408] <= 8'h10 ;
			data[81409] <= 8'h10 ;
			data[81410] <= 8'h10 ;
			data[81411] <= 8'h10 ;
			data[81412] <= 8'h10 ;
			data[81413] <= 8'h10 ;
			data[81414] <= 8'h10 ;
			data[81415] <= 8'h10 ;
			data[81416] <= 8'h10 ;
			data[81417] <= 8'h10 ;
			data[81418] <= 8'h10 ;
			data[81419] <= 8'h10 ;
			data[81420] <= 8'h10 ;
			data[81421] <= 8'h10 ;
			data[81422] <= 8'h10 ;
			data[81423] <= 8'h10 ;
			data[81424] <= 8'h10 ;
			data[81425] <= 8'h10 ;
			data[81426] <= 8'h10 ;
			data[81427] <= 8'h10 ;
			data[81428] <= 8'h10 ;
			data[81429] <= 8'h10 ;
			data[81430] <= 8'h10 ;
			data[81431] <= 8'h10 ;
			data[81432] <= 8'h10 ;
			data[81433] <= 8'h10 ;
			data[81434] <= 8'h10 ;
			data[81435] <= 8'h10 ;
			data[81436] <= 8'h10 ;
			data[81437] <= 8'h10 ;
			data[81438] <= 8'h10 ;
			data[81439] <= 8'h10 ;
			data[81440] <= 8'h10 ;
			data[81441] <= 8'h10 ;
			data[81442] <= 8'h10 ;
			data[81443] <= 8'h10 ;
			data[81444] <= 8'h10 ;
			data[81445] <= 8'h10 ;
			data[81446] <= 8'h10 ;
			data[81447] <= 8'h10 ;
			data[81448] <= 8'h10 ;
			data[81449] <= 8'h10 ;
			data[81450] <= 8'h10 ;
			data[81451] <= 8'h10 ;
			data[81452] <= 8'h10 ;
			data[81453] <= 8'h10 ;
			data[81454] <= 8'h10 ;
			data[81455] <= 8'h10 ;
			data[81456] <= 8'h10 ;
			data[81457] <= 8'h10 ;
			data[81458] <= 8'h10 ;
			data[81459] <= 8'h10 ;
			data[81460] <= 8'h10 ;
			data[81461] <= 8'h10 ;
			data[81462] <= 8'h10 ;
			data[81463] <= 8'h10 ;
			data[81464] <= 8'h10 ;
			data[81465] <= 8'h10 ;
			data[81466] <= 8'h10 ;
			data[81467] <= 8'h10 ;
			data[81468] <= 8'h10 ;
			data[81469] <= 8'h10 ;
			data[81470] <= 8'h10 ;
			data[81471] <= 8'h10 ;
			data[81472] <= 8'h10 ;
			data[81473] <= 8'h10 ;
			data[81474] <= 8'h10 ;
			data[81475] <= 8'h10 ;
			data[81476] <= 8'h10 ;
			data[81477] <= 8'h10 ;
			data[81478] <= 8'h10 ;
			data[81479] <= 8'h10 ;
			data[81480] <= 8'h10 ;
			data[81481] <= 8'h10 ;
			data[81482] <= 8'h10 ;
			data[81483] <= 8'h10 ;
			data[81484] <= 8'h10 ;
			data[81485] <= 8'h10 ;
			data[81486] <= 8'h10 ;
			data[81487] <= 8'h10 ;
			data[81488] <= 8'h10 ;
			data[81489] <= 8'h10 ;
			data[81490] <= 8'h10 ;
			data[81491] <= 8'h10 ;
			data[81492] <= 8'h10 ;
			data[81493] <= 8'h10 ;
			data[81494] <= 8'h10 ;
			data[81495] <= 8'h10 ;
			data[81496] <= 8'h10 ;
			data[81497] <= 8'h10 ;
			data[81498] <= 8'h10 ;
			data[81499] <= 8'h10 ;
			data[81500] <= 8'h10 ;
			data[81501] <= 8'h10 ;
			data[81502] <= 8'h10 ;
			data[81503] <= 8'h10 ;
			data[81504] <= 8'h10 ;
			data[81505] <= 8'h10 ;
			data[81506] <= 8'h10 ;
			data[81507] <= 8'h10 ;
			data[81508] <= 8'h10 ;
			data[81509] <= 8'h10 ;
			data[81510] <= 8'h10 ;
			data[81511] <= 8'h10 ;
			data[81512] <= 8'h10 ;
			data[81513] <= 8'h10 ;
			data[81514] <= 8'h10 ;
			data[81515] <= 8'h10 ;
			data[81516] <= 8'h10 ;
			data[81517] <= 8'h10 ;
			data[81518] <= 8'h10 ;
			data[81519] <= 8'h10 ;
			data[81520] <= 8'h10 ;
			data[81521] <= 8'h10 ;
			data[81522] <= 8'h10 ;
			data[81523] <= 8'h10 ;
			data[81524] <= 8'h10 ;
			data[81525] <= 8'h10 ;
			data[81526] <= 8'h10 ;
			data[81527] <= 8'h10 ;
			data[81528] <= 8'h10 ;
			data[81529] <= 8'h10 ;
			data[81530] <= 8'h10 ;
			data[81531] <= 8'h10 ;
			data[81532] <= 8'h10 ;
			data[81533] <= 8'h10 ;
			data[81534] <= 8'h10 ;
			data[81535] <= 8'h10 ;
			data[81536] <= 8'h10 ;
			data[81537] <= 8'h10 ;
			data[81538] <= 8'h10 ;
			data[81539] <= 8'h10 ;
			data[81540] <= 8'h10 ;
			data[81541] <= 8'h10 ;
			data[81542] <= 8'h10 ;
			data[81543] <= 8'h10 ;
			data[81544] <= 8'h10 ;
			data[81545] <= 8'h10 ;
			data[81546] <= 8'h10 ;
			data[81547] <= 8'h10 ;
			data[81548] <= 8'h10 ;
			data[81549] <= 8'h10 ;
			data[81550] <= 8'h10 ;
			data[81551] <= 8'h10 ;
			data[81552] <= 8'h10 ;
			data[81553] <= 8'h10 ;
			data[81554] <= 8'h10 ;
			data[81555] <= 8'h10 ;
			data[81556] <= 8'h10 ;
			data[81557] <= 8'h10 ;
			data[81558] <= 8'h10 ;
			data[81559] <= 8'h10 ;
			data[81560] <= 8'h10 ;
			data[81561] <= 8'h10 ;
			data[81562] <= 8'h10 ;
			data[81563] <= 8'h10 ;
			data[81564] <= 8'h10 ;
			data[81565] <= 8'h10 ;
			data[81566] <= 8'h10 ;
			data[81567] <= 8'h10 ;
			data[81568] <= 8'h10 ;
			data[81569] <= 8'h10 ;
			data[81570] <= 8'h10 ;
			data[81571] <= 8'h10 ;
			data[81572] <= 8'h10 ;
			data[81573] <= 8'h10 ;
			data[81574] <= 8'h10 ;
			data[81575] <= 8'h10 ;
			data[81576] <= 8'h10 ;
			data[81577] <= 8'h10 ;
			data[81578] <= 8'h10 ;
			data[81579] <= 8'h10 ;
			data[81580] <= 8'h10 ;
			data[81581] <= 8'h10 ;
			data[81582] <= 8'h10 ;
			data[81583] <= 8'h10 ;
			data[81584] <= 8'h10 ;
			data[81585] <= 8'h10 ;
			data[81586] <= 8'h10 ;
			data[81587] <= 8'h10 ;
			data[81588] <= 8'h10 ;
			data[81589] <= 8'h10 ;
			data[81590] <= 8'h10 ;
			data[81591] <= 8'h10 ;
			data[81592] <= 8'h10 ;
			data[81593] <= 8'h10 ;
			data[81594] <= 8'h10 ;
			data[81595] <= 8'h10 ;
			data[81596] <= 8'h10 ;
			data[81597] <= 8'h10 ;
			data[81598] <= 8'h10 ;
			data[81599] <= 8'h10 ;
			data[81600] <= 8'h10 ;
			data[81601] <= 8'h10 ;
			data[81602] <= 8'h10 ;
			data[81603] <= 8'h10 ;
			data[81604] <= 8'h10 ;
			data[81605] <= 8'h10 ;
			data[81606] <= 8'h10 ;
			data[81607] <= 8'h10 ;
			data[81608] <= 8'h10 ;
			data[81609] <= 8'h10 ;
			data[81610] <= 8'h10 ;
			data[81611] <= 8'h10 ;
			data[81612] <= 8'h10 ;
			data[81613] <= 8'h10 ;
			data[81614] <= 8'h10 ;
			data[81615] <= 8'h10 ;
			data[81616] <= 8'h10 ;
			data[81617] <= 8'h10 ;
			data[81618] <= 8'h10 ;
			data[81619] <= 8'h10 ;
			data[81620] <= 8'h10 ;
			data[81621] <= 8'h10 ;
			data[81622] <= 8'h10 ;
			data[81623] <= 8'h10 ;
			data[81624] <= 8'h10 ;
			data[81625] <= 8'h10 ;
			data[81626] <= 8'h10 ;
			data[81627] <= 8'h10 ;
			data[81628] <= 8'h10 ;
			data[81629] <= 8'h10 ;
			data[81630] <= 8'h10 ;
			data[81631] <= 8'h10 ;
			data[81632] <= 8'h10 ;
			data[81633] <= 8'h10 ;
			data[81634] <= 8'h10 ;
			data[81635] <= 8'h10 ;
			data[81636] <= 8'h10 ;
			data[81637] <= 8'h10 ;
			data[81638] <= 8'h10 ;
			data[81639] <= 8'h10 ;
			data[81640] <= 8'h10 ;
			data[81641] <= 8'h10 ;
			data[81642] <= 8'h10 ;
			data[81643] <= 8'h10 ;
			data[81644] <= 8'h10 ;
			data[81645] <= 8'h10 ;
			data[81646] <= 8'h10 ;
			data[81647] <= 8'h10 ;
			data[81648] <= 8'h10 ;
			data[81649] <= 8'h10 ;
			data[81650] <= 8'h10 ;
			data[81651] <= 8'h10 ;
			data[81652] <= 8'h10 ;
			data[81653] <= 8'h10 ;
			data[81654] <= 8'h10 ;
			data[81655] <= 8'h10 ;
			data[81656] <= 8'h10 ;
			data[81657] <= 8'h10 ;
			data[81658] <= 8'h10 ;
			data[81659] <= 8'h10 ;
			data[81660] <= 8'h10 ;
			data[81661] <= 8'h10 ;
			data[81662] <= 8'h10 ;
			data[81663] <= 8'h10 ;
			data[81664] <= 8'h10 ;
			data[81665] <= 8'h10 ;
			data[81666] <= 8'h10 ;
			data[81667] <= 8'h10 ;
			data[81668] <= 8'h10 ;
			data[81669] <= 8'h10 ;
			data[81670] <= 8'h10 ;
			data[81671] <= 8'h10 ;
			data[81672] <= 8'h10 ;
			data[81673] <= 8'h10 ;
			data[81674] <= 8'h10 ;
			data[81675] <= 8'h10 ;
			data[81676] <= 8'h10 ;
			data[81677] <= 8'h10 ;
			data[81678] <= 8'h10 ;
			data[81679] <= 8'h10 ;
			data[81680] <= 8'h10 ;
			data[81681] <= 8'h10 ;
			data[81682] <= 8'h10 ;
			data[81683] <= 8'h10 ;
			data[81684] <= 8'h10 ;
			data[81685] <= 8'h10 ;
			data[81686] <= 8'h10 ;
			data[81687] <= 8'h10 ;
			data[81688] <= 8'h10 ;
			data[81689] <= 8'h10 ;
			data[81690] <= 8'h10 ;
			data[81691] <= 8'h10 ;
			data[81692] <= 8'h10 ;
			data[81693] <= 8'h10 ;
			data[81694] <= 8'h10 ;
			data[81695] <= 8'h10 ;
			data[81696] <= 8'h10 ;
			data[81697] <= 8'h10 ;
			data[81698] <= 8'h10 ;
			data[81699] <= 8'h10 ;
			data[81700] <= 8'h10 ;
			data[81701] <= 8'h10 ;
			data[81702] <= 8'h10 ;
			data[81703] <= 8'h10 ;
			data[81704] <= 8'h10 ;
			data[81705] <= 8'h10 ;
			data[81706] <= 8'h10 ;
			data[81707] <= 8'h10 ;
			data[81708] <= 8'h10 ;
			data[81709] <= 8'h10 ;
			data[81710] <= 8'h10 ;
			data[81711] <= 8'h10 ;
			data[81712] <= 8'h10 ;
			data[81713] <= 8'h10 ;
			data[81714] <= 8'h10 ;
			data[81715] <= 8'h10 ;
			data[81716] <= 8'h10 ;
			data[81717] <= 8'h10 ;
			data[81718] <= 8'h10 ;
			data[81719] <= 8'h10 ;
			data[81720] <= 8'h10 ;
			data[81721] <= 8'h10 ;
			data[81722] <= 8'h10 ;
			data[81723] <= 8'h10 ;
			data[81724] <= 8'h10 ;
			data[81725] <= 8'h10 ;
			data[81726] <= 8'h10 ;
			data[81727] <= 8'h10 ;
			data[81728] <= 8'h10 ;
			data[81729] <= 8'h10 ;
			data[81730] <= 8'h10 ;
			data[81731] <= 8'h10 ;
			data[81732] <= 8'h10 ;
			data[81733] <= 8'h10 ;
			data[81734] <= 8'h10 ;
			data[81735] <= 8'h10 ;
			data[81736] <= 8'h10 ;
			data[81737] <= 8'h10 ;
			data[81738] <= 8'h10 ;
			data[81739] <= 8'h10 ;
			data[81740] <= 8'h10 ;
			data[81741] <= 8'h10 ;
			data[81742] <= 8'h10 ;
			data[81743] <= 8'h10 ;
			data[81744] <= 8'h10 ;
			data[81745] <= 8'h10 ;
			data[81746] <= 8'h10 ;
			data[81747] <= 8'h10 ;
			data[81748] <= 8'h10 ;
			data[81749] <= 8'h10 ;
			data[81750] <= 8'h10 ;
			data[81751] <= 8'h10 ;
			data[81752] <= 8'h10 ;
			data[81753] <= 8'h10 ;
			data[81754] <= 8'h10 ;
			data[81755] <= 8'h10 ;
			data[81756] <= 8'h10 ;
			data[81757] <= 8'h10 ;
			data[81758] <= 8'h10 ;
			data[81759] <= 8'h10 ;
			data[81760] <= 8'h10 ;
			data[81761] <= 8'h10 ;
			data[81762] <= 8'h10 ;
			data[81763] <= 8'h10 ;
			data[81764] <= 8'h10 ;
			data[81765] <= 8'h10 ;
			data[81766] <= 8'h10 ;
			data[81767] <= 8'h10 ;
			data[81768] <= 8'h10 ;
			data[81769] <= 8'h10 ;
			data[81770] <= 8'h10 ;
			data[81771] <= 8'h10 ;
			data[81772] <= 8'h10 ;
			data[81773] <= 8'h10 ;
			data[81774] <= 8'h10 ;
			data[81775] <= 8'h10 ;
			data[81776] <= 8'h10 ;
			data[81777] <= 8'h10 ;
			data[81778] <= 8'h10 ;
			data[81779] <= 8'h10 ;
			data[81780] <= 8'h10 ;
			data[81781] <= 8'h10 ;
			data[81782] <= 8'h10 ;
			data[81783] <= 8'h10 ;
			data[81784] <= 8'h10 ;
			data[81785] <= 8'h10 ;
			data[81786] <= 8'h10 ;
			data[81787] <= 8'h10 ;
			data[81788] <= 8'h10 ;
			data[81789] <= 8'h10 ;
			data[81790] <= 8'h10 ;
			data[81791] <= 8'h10 ;
			data[81792] <= 8'h10 ;
			data[81793] <= 8'h10 ;
			data[81794] <= 8'h10 ;
			data[81795] <= 8'h10 ;
			data[81796] <= 8'h10 ;
			data[81797] <= 8'h10 ;
			data[81798] <= 8'h10 ;
			data[81799] <= 8'h10 ;
			data[81800] <= 8'h10 ;
			data[81801] <= 8'h10 ;
			data[81802] <= 8'h10 ;
			data[81803] <= 8'h10 ;
			data[81804] <= 8'h10 ;
			data[81805] <= 8'h10 ;
			data[81806] <= 8'h10 ;
			data[81807] <= 8'h10 ;
			data[81808] <= 8'h10 ;
			data[81809] <= 8'h10 ;
			data[81810] <= 8'h10 ;
			data[81811] <= 8'h10 ;
			data[81812] <= 8'h10 ;
			data[81813] <= 8'h10 ;
			data[81814] <= 8'h10 ;
			data[81815] <= 8'h10 ;
			data[81816] <= 8'h10 ;
			data[81817] <= 8'h10 ;
			data[81818] <= 8'h10 ;
			data[81819] <= 8'h10 ;
			data[81820] <= 8'h10 ;
			data[81821] <= 8'h10 ;
			data[81822] <= 8'h10 ;
			data[81823] <= 8'h10 ;
			data[81824] <= 8'h10 ;
			data[81825] <= 8'h10 ;
			data[81826] <= 8'h10 ;
			data[81827] <= 8'h10 ;
			data[81828] <= 8'h10 ;
			data[81829] <= 8'h10 ;
			data[81830] <= 8'h10 ;
			data[81831] <= 8'h10 ;
			data[81832] <= 8'h10 ;
			data[81833] <= 8'h10 ;
			data[81834] <= 8'h10 ;
			data[81835] <= 8'h10 ;
			data[81836] <= 8'h10 ;
			data[81837] <= 8'h10 ;
			data[81838] <= 8'h10 ;
			data[81839] <= 8'h10 ;
			data[81840] <= 8'h10 ;
			data[81841] <= 8'h10 ;
			data[81842] <= 8'h10 ;
			data[81843] <= 8'h10 ;
			data[81844] <= 8'h10 ;
			data[81845] <= 8'h10 ;
			data[81846] <= 8'h10 ;
			data[81847] <= 8'h10 ;
			data[81848] <= 8'h10 ;
			data[81849] <= 8'h10 ;
			data[81850] <= 8'h10 ;
			data[81851] <= 8'h10 ;
			data[81852] <= 8'h10 ;
			data[81853] <= 8'h10 ;
			data[81854] <= 8'h10 ;
			data[81855] <= 8'h10 ;
			data[81856] <= 8'h10 ;
			data[81857] <= 8'h10 ;
			data[81858] <= 8'h10 ;
			data[81859] <= 8'h10 ;
			data[81860] <= 8'h10 ;
			data[81861] <= 8'h10 ;
			data[81862] <= 8'h10 ;
			data[81863] <= 8'h10 ;
			data[81864] <= 8'h10 ;
			data[81865] <= 8'h10 ;
			data[81866] <= 8'h10 ;
			data[81867] <= 8'h10 ;
			data[81868] <= 8'h10 ;
			data[81869] <= 8'h10 ;
			data[81870] <= 8'h10 ;
			data[81871] <= 8'h10 ;
			data[81872] <= 8'h10 ;
			data[81873] <= 8'h10 ;
			data[81874] <= 8'h10 ;
			data[81875] <= 8'h10 ;
			data[81876] <= 8'h10 ;
			data[81877] <= 8'h10 ;
			data[81878] <= 8'h10 ;
			data[81879] <= 8'h10 ;
			data[81880] <= 8'h10 ;
			data[81881] <= 8'h10 ;
			data[81882] <= 8'h10 ;
			data[81883] <= 8'h10 ;
			data[81884] <= 8'h10 ;
			data[81885] <= 8'h10 ;
			data[81886] <= 8'h10 ;
			data[81887] <= 8'h10 ;
			data[81888] <= 8'h10 ;
			data[81889] <= 8'h10 ;
			data[81890] <= 8'h10 ;
			data[81891] <= 8'h10 ;
			data[81892] <= 8'h10 ;
			data[81893] <= 8'h10 ;
			data[81894] <= 8'h10 ;
			data[81895] <= 8'h10 ;
			data[81896] <= 8'h10 ;
			data[81897] <= 8'h10 ;
			data[81898] <= 8'h10 ;
			data[81899] <= 8'h10 ;
			data[81900] <= 8'h10 ;
			data[81901] <= 8'h10 ;
			data[81902] <= 8'h10 ;
			data[81903] <= 8'h10 ;
			data[81904] <= 8'h10 ;
			data[81905] <= 8'h10 ;
			data[81906] <= 8'h10 ;
			data[81907] <= 8'h10 ;
			data[81908] <= 8'h10 ;
			data[81909] <= 8'h10 ;
			data[81910] <= 8'h10 ;
			data[81911] <= 8'h10 ;
			data[81912] <= 8'h10 ;
			data[81913] <= 8'h10 ;
			data[81914] <= 8'h10 ;
			data[81915] <= 8'h10 ;
			data[81916] <= 8'h10 ;
			data[81917] <= 8'h10 ;
			data[81918] <= 8'h10 ;
			data[81919] <= 8'h10 ;
			data[81920] <= 8'h10 ;
			data[81921] <= 8'h10 ;
			data[81922] <= 8'h10 ;
			data[81923] <= 8'h10 ;
			data[81924] <= 8'h10 ;
			data[81925] <= 8'h10 ;
			data[81926] <= 8'h10 ;
			data[81927] <= 8'h10 ;
			data[81928] <= 8'h10 ;
			data[81929] <= 8'h10 ;
			data[81930] <= 8'h10 ;
			data[81931] <= 8'h10 ;
			data[81932] <= 8'h10 ;
			data[81933] <= 8'h10 ;
			data[81934] <= 8'h10 ;
			data[81935] <= 8'h10 ;
			data[81936] <= 8'h10 ;
			data[81937] <= 8'h10 ;
			data[81938] <= 8'h10 ;
			data[81939] <= 8'h10 ;
			data[81940] <= 8'h10 ;
			data[81941] <= 8'h10 ;
			data[81942] <= 8'h10 ;
			data[81943] <= 8'h10 ;
			data[81944] <= 8'h10 ;
			data[81945] <= 8'h10 ;
			data[81946] <= 8'h10 ;
			data[81947] <= 8'h10 ;
			data[81948] <= 8'h10 ;
			data[81949] <= 8'h10 ;
			data[81950] <= 8'h10 ;
			data[81951] <= 8'h10 ;
			data[81952] <= 8'h10 ;
			data[81953] <= 8'h10 ;
			data[81954] <= 8'h10 ;
			data[81955] <= 8'h10 ;
			data[81956] <= 8'h10 ;
			data[81957] <= 8'h10 ;
			data[81958] <= 8'h10 ;
			data[81959] <= 8'h10 ;
			data[81960] <= 8'h10 ;
			data[81961] <= 8'h10 ;
			data[81962] <= 8'h10 ;
			data[81963] <= 8'h10 ;
			data[81964] <= 8'h10 ;
			data[81965] <= 8'h10 ;
			data[81966] <= 8'h10 ;
			data[81967] <= 8'h10 ;
			data[81968] <= 8'h10 ;
			data[81969] <= 8'h10 ;
			data[81970] <= 8'h10 ;
			data[81971] <= 8'h10 ;
			data[81972] <= 8'h10 ;
			data[81973] <= 8'h10 ;
			data[81974] <= 8'h10 ;
			data[81975] <= 8'h10 ;
			data[81976] <= 8'h10 ;
			data[81977] <= 8'h10 ;
			data[81978] <= 8'h10 ;
			data[81979] <= 8'h10 ;
			data[81980] <= 8'h10 ;
			data[81981] <= 8'h10 ;
			data[81982] <= 8'h10 ;
			data[81983] <= 8'h10 ;
			data[81984] <= 8'h10 ;
			data[81985] <= 8'h10 ;
			data[81986] <= 8'h10 ;
			data[81987] <= 8'h10 ;
			data[81988] <= 8'h10 ;
			data[81989] <= 8'h10 ;
			data[81990] <= 8'h10 ;
			data[81991] <= 8'h10 ;
			data[81992] <= 8'h10 ;
			data[81993] <= 8'h10 ;
			data[81994] <= 8'h10 ;
			data[81995] <= 8'h10 ;
			data[81996] <= 8'h10 ;
			data[81997] <= 8'h10 ;
			data[81998] <= 8'h10 ;
			data[81999] <= 8'h10 ;
			data[82000] <= 8'h10 ;
			data[82001] <= 8'h10 ;
			data[82002] <= 8'h10 ;
			data[82003] <= 8'h10 ;
			data[82004] <= 8'h10 ;
			data[82005] <= 8'h10 ;
			data[82006] <= 8'h10 ;
			data[82007] <= 8'h10 ;
			data[82008] <= 8'h10 ;
			data[82009] <= 8'h10 ;
			data[82010] <= 8'h10 ;
			data[82011] <= 8'h10 ;
			data[82012] <= 8'h10 ;
			data[82013] <= 8'h10 ;
			data[82014] <= 8'h10 ;
			data[82015] <= 8'h10 ;
			data[82016] <= 8'h10 ;
			data[82017] <= 8'h10 ;
			data[82018] <= 8'h10 ;
			data[82019] <= 8'h10 ;
			data[82020] <= 8'h10 ;
			data[82021] <= 8'h10 ;
			data[82022] <= 8'h10 ;
			data[82023] <= 8'h10 ;
			data[82024] <= 8'h10 ;
			data[82025] <= 8'h10 ;
			data[82026] <= 8'h10 ;
			data[82027] <= 8'h10 ;
			data[82028] <= 8'h10 ;
			data[82029] <= 8'h10 ;
			data[82030] <= 8'h10 ;
			data[82031] <= 8'h10 ;
			data[82032] <= 8'h10 ;
			data[82033] <= 8'h10 ;
			data[82034] <= 8'h10 ;
			data[82035] <= 8'h10 ;
			data[82036] <= 8'h10 ;
			data[82037] <= 8'h10 ;
			data[82038] <= 8'h10 ;
			data[82039] <= 8'h10 ;
			data[82040] <= 8'h10 ;
			data[82041] <= 8'h10 ;
			data[82042] <= 8'h10 ;
			data[82043] <= 8'h10 ;
			data[82044] <= 8'h10 ;
			data[82045] <= 8'h10 ;
			data[82046] <= 8'h10 ;
			data[82047] <= 8'h10 ;
			data[82048] <= 8'h10 ;
			data[82049] <= 8'h10 ;
			data[82050] <= 8'h10 ;
			data[82051] <= 8'h10 ;
			data[82052] <= 8'h10 ;
			data[82053] <= 8'h10 ;
			data[82054] <= 8'h10 ;
			data[82055] <= 8'h10 ;
			data[82056] <= 8'h10 ;
			data[82057] <= 8'h10 ;
			data[82058] <= 8'h10 ;
			data[82059] <= 8'h10 ;
			data[82060] <= 8'h10 ;
			data[82061] <= 8'h10 ;
			data[82062] <= 8'h10 ;
			data[82063] <= 8'h10 ;
			data[82064] <= 8'h10 ;
			data[82065] <= 8'h10 ;
			data[82066] <= 8'h10 ;
			data[82067] <= 8'h10 ;
			data[82068] <= 8'h10 ;
			data[82069] <= 8'h10 ;
			data[82070] <= 8'h10 ;
			data[82071] <= 8'h10 ;
			data[82072] <= 8'h10 ;
			data[82073] <= 8'h10 ;
			data[82074] <= 8'h10 ;
			data[82075] <= 8'h10 ;
			data[82076] <= 8'h10 ;
			data[82077] <= 8'h10 ;
			data[82078] <= 8'h10 ;
			data[82079] <= 8'h10 ;
			data[82080] <= 8'h10 ;
			data[82081] <= 8'h10 ;
			data[82082] <= 8'h10 ;
			data[82083] <= 8'h10 ;
			data[82084] <= 8'h10 ;
			data[82085] <= 8'h10 ;
			data[82086] <= 8'h10 ;
			data[82087] <= 8'h10 ;
			data[82088] <= 8'h10 ;
			data[82089] <= 8'h10 ;
			data[82090] <= 8'h10 ;
			data[82091] <= 8'h10 ;
			data[82092] <= 8'h10 ;
			data[82093] <= 8'h10 ;
			data[82094] <= 8'h10 ;
			data[82095] <= 8'h10 ;
			data[82096] <= 8'h10 ;
			data[82097] <= 8'h10 ;
			data[82098] <= 8'h10 ;
			data[82099] <= 8'h10 ;
			data[82100] <= 8'h10 ;
			data[82101] <= 8'h10 ;
			data[82102] <= 8'h10 ;
			data[82103] <= 8'h10 ;
			data[82104] <= 8'h10 ;
			data[82105] <= 8'h10 ;
			data[82106] <= 8'h10 ;
			data[82107] <= 8'h10 ;
			data[82108] <= 8'h10 ;
			data[82109] <= 8'h10 ;
			data[82110] <= 8'h10 ;
			data[82111] <= 8'h10 ;
			data[82112] <= 8'h10 ;
			data[82113] <= 8'h10 ;
			data[82114] <= 8'h10 ;
			data[82115] <= 8'h10 ;
			data[82116] <= 8'h10 ;
			data[82117] <= 8'h10 ;
			data[82118] <= 8'h10 ;
			data[82119] <= 8'h10 ;
			data[82120] <= 8'h10 ;
			data[82121] <= 8'h10 ;
			data[82122] <= 8'h10 ;
			data[82123] <= 8'h10 ;
			data[82124] <= 8'h10 ;
			data[82125] <= 8'h10 ;
			data[82126] <= 8'h10 ;
			data[82127] <= 8'h10 ;
			data[82128] <= 8'h10 ;
			data[82129] <= 8'h10 ;
			data[82130] <= 8'h10 ;
			data[82131] <= 8'h10 ;
			data[82132] <= 8'h10 ;
			data[82133] <= 8'h10 ;
			data[82134] <= 8'h10 ;
			data[82135] <= 8'h10 ;
			data[82136] <= 8'h10 ;
			data[82137] <= 8'h10 ;
			data[82138] <= 8'h10 ;
			data[82139] <= 8'h10 ;
			data[82140] <= 8'h10 ;
			data[82141] <= 8'h10 ;
			data[82142] <= 8'h10 ;
			data[82143] <= 8'h10 ;
			data[82144] <= 8'h10 ;
			data[82145] <= 8'h10 ;
			data[82146] <= 8'h10 ;
			data[82147] <= 8'h10 ;
			data[82148] <= 8'h10 ;
			data[82149] <= 8'h10 ;
			data[82150] <= 8'h10 ;
			data[82151] <= 8'h10 ;
			data[82152] <= 8'h10 ;
			data[82153] <= 8'h10 ;
			data[82154] <= 8'h10 ;
			data[82155] <= 8'h10 ;
			data[82156] <= 8'h10 ;
			data[82157] <= 8'h10 ;
			data[82158] <= 8'h10 ;
			data[82159] <= 8'h10 ;
			data[82160] <= 8'h10 ;
			data[82161] <= 8'h10 ;
			data[82162] <= 8'h10 ;
			data[82163] <= 8'h10 ;
			data[82164] <= 8'h10 ;
			data[82165] <= 8'h10 ;
			data[82166] <= 8'h10 ;
			data[82167] <= 8'h10 ;
			data[82168] <= 8'h10 ;
			data[82169] <= 8'h10 ;
			data[82170] <= 8'h10 ;
			data[82171] <= 8'h10 ;
			data[82172] <= 8'h10 ;
			data[82173] <= 8'h10 ;
			data[82174] <= 8'h10 ;
			data[82175] <= 8'h10 ;
			data[82176] <= 8'h10 ;
			data[82177] <= 8'h10 ;
			data[82178] <= 8'h10 ;
			data[82179] <= 8'h10 ;
			data[82180] <= 8'h10 ;
			data[82181] <= 8'h10 ;
			data[82182] <= 8'h10 ;
			data[82183] <= 8'h10 ;
			data[82184] <= 8'h10 ;
			data[82185] <= 8'h10 ;
			data[82186] <= 8'h10 ;
			data[82187] <= 8'h10 ;
			data[82188] <= 8'h10 ;
			data[82189] <= 8'h10 ;
			data[82190] <= 8'h10 ;
			data[82191] <= 8'h10 ;
			data[82192] <= 8'h10 ;
			data[82193] <= 8'h10 ;
			data[82194] <= 8'h10 ;
			data[82195] <= 8'h10 ;
			data[82196] <= 8'h10 ;
			data[82197] <= 8'h10 ;
			data[82198] <= 8'h10 ;
			data[82199] <= 8'h10 ;
			data[82200] <= 8'h10 ;
			data[82201] <= 8'h10 ;
			data[82202] <= 8'h10 ;
			data[82203] <= 8'h10 ;
			data[82204] <= 8'h10 ;
			data[82205] <= 8'h10 ;
			data[82206] <= 8'h10 ;
			data[82207] <= 8'h10 ;
			data[82208] <= 8'h10 ;
			data[82209] <= 8'h10 ;
			data[82210] <= 8'h10 ;
			data[82211] <= 8'h10 ;
			data[82212] <= 8'h10 ;
			data[82213] <= 8'h10 ;
			data[82214] <= 8'h10 ;
			data[82215] <= 8'h10 ;
			data[82216] <= 8'h10 ;
			data[82217] <= 8'h10 ;
			data[82218] <= 8'h10 ;
			data[82219] <= 8'h10 ;
			data[82220] <= 8'h10 ;
			data[82221] <= 8'h10 ;
			data[82222] <= 8'h10 ;
			data[82223] <= 8'h10 ;
			data[82224] <= 8'h10 ;
			data[82225] <= 8'h10 ;
			data[82226] <= 8'h10 ;
			data[82227] <= 8'h10 ;
			data[82228] <= 8'h10 ;
			data[82229] <= 8'h10 ;
			data[82230] <= 8'h10 ;
			data[82231] <= 8'h10 ;
			data[82232] <= 8'h10 ;
			data[82233] <= 8'h10 ;
			data[82234] <= 8'h10 ;
			data[82235] <= 8'h10 ;
			data[82236] <= 8'h10 ;
			data[82237] <= 8'h10 ;
			data[82238] <= 8'h10 ;
			data[82239] <= 8'h10 ;
			data[82240] <= 8'h10 ;
			data[82241] <= 8'h10 ;
			data[82242] <= 8'h10 ;
			data[82243] <= 8'h10 ;
			data[82244] <= 8'h10 ;
			data[82245] <= 8'h10 ;
			data[82246] <= 8'h10 ;
			data[82247] <= 8'h10 ;
			data[82248] <= 8'h10 ;
			data[82249] <= 8'h10 ;
			data[82250] <= 8'h10 ;
			data[82251] <= 8'h10 ;
			data[82252] <= 8'h10 ;
			data[82253] <= 8'h10 ;
			data[82254] <= 8'h10 ;
			data[82255] <= 8'h10 ;
			data[82256] <= 8'h10 ;
			data[82257] <= 8'h10 ;
			data[82258] <= 8'h10 ;
			data[82259] <= 8'h10 ;
			data[82260] <= 8'h10 ;
			data[82261] <= 8'h10 ;
			data[82262] <= 8'h10 ;
			data[82263] <= 8'h10 ;
			data[82264] <= 8'h10 ;
			data[82265] <= 8'h10 ;
			data[82266] <= 8'h10 ;
			data[82267] <= 8'h10 ;
			data[82268] <= 8'h10 ;
			data[82269] <= 8'h10 ;
			data[82270] <= 8'h10 ;
			data[82271] <= 8'h10 ;
			data[82272] <= 8'h10 ;
			data[82273] <= 8'h10 ;
			data[82274] <= 8'h10 ;
			data[82275] <= 8'h10 ;
			data[82276] <= 8'h10 ;
			data[82277] <= 8'h10 ;
			data[82278] <= 8'h10 ;
			data[82279] <= 8'h10 ;
			data[82280] <= 8'h10 ;
			data[82281] <= 8'h10 ;
			data[82282] <= 8'h10 ;
			data[82283] <= 8'h10 ;
			data[82284] <= 8'h10 ;
			data[82285] <= 8'h10 ;
			data[82286] <= 8'h10 ;
			data[82287] <= 8'h10 ;
			data[82288] <= 8'h10 ;
			data[82289] <= 8'h10 ;
			data[82290] <= 8'h10 ;
			data[82291] <= 8'h10 ;
			data[82292] <= 8'h10 ;
			data[82293] <= 8'h10 ;
			data[82294] <= 8'h10 ;
			data[82295] <= 8'h10 ;
			data[82296] <= 8'h10 ;
			data[82297] <= 8'h10 ;
			data[82298] <= 8'h10 ;
			data[82299] <= 8'h10 ;
			data[82300] <= 8'h10 ;
			data[82301] <= 8'h10 ;
			data[82302] <= 8'h10 ;
			data[82303] <= 8'h10 ;
			data[82304] <= 8'h10 ;
			data[82305] <= 8'h10 ;
			data[82306] <= 8'h10 ;
			data[82307] <= 8'h10 ;
			data[82308] <= 8'h10 ;
			data[82309] <= 8'h10 ;
			data[82310] <= 8'h10 ;
			data[82311] <= 8'h10 ;
			data[82312] <= 8'h10 ;
			data[82313] <= 8'h10 ;
			data[82314] <= 8'h10 ;
			data[82315] <= 8'h10 ;
			data[82316] <= 8'h10 ;
			data[82317] <= 8'h10 ;
			data[82318] <= 8'h10 ;
			data[82319] <= 8'h10 ;
			data[82320] <= 8'h10 ;
			data[82321] <= 8'h10 ;
			data[82322] <= 8'h10 ;
			data[82323] <= 8'h10 ;
			data[82324] <= 8'h10 ;
			data[82325] <= 8'h10 ;
			data[82326] <= 8'h10 ;
			data[82327] <= 8'h10 ;
			data[82328] <= 8'h10 ;
			data[82329] <= 8'h10 ;
			data[82330] <= 8'h10 ;
			data[82331] <= 8'h10 ;
			data[82332] <= 8'h10 ;
			data[82333] <= 8'h10 ;
			data[82334] <= 8'h10 ;
			data[82335] <= 8'h10 ;
			data[82336] <= 8'h10 ;
			data[82337] <= 8'h10 ;
			data[82338] <= 8'h10 ;
			data[82339] <= 8'h10 ;
			data[82340] <= 8'h10 ;
			data[82341] <= 8'h10 ;
			data[82342] <= 8'h10 ;
			data[82343] <= 8'h10 ;
			data[82344] <= 8'h10 ;
			data[82345] <= 8'h10 ;
			data[82346] <= 8'h10 ;
			data[82347] <= 8'h10 ;
			data[82348] <= 8'h10 ;
			data[82349] <= 8'h10 ;
			data[82350] <= 8'h10 ;
			data[82351] <= 8'h10 ;
			data[82352] <= 8'h10 ;
			data[82353] <= 8'h10 ;
			data[82354] <= 8'h10 ;
			data[82355] <= 8'h10 ;
			data[82356] <= 8'h10 ;
			data[82357] <= 8'h10 ;
			data[82358] <= 8'h10 ;
			data[82359] <= 8'h10 ;
			data[82360] <= 8'h10 ;
			data[82361] <= 8'h10 ;
			data[82362] <= 8'h10 ;
			data[82363] <= 8'h10 ;
			data[82364] <= 8'h10 ;
			data[82365] <= 8'h10 ;
			data[82366] <= 8'h10 ;
			data[82367] <= 8'h10 ;
			data[82368] <= 8'h10 ;
			data[82369] <= 8'h10 ;
			data[82370] <= 8'h10 ;
			data[82371] <= 8'h10 ;
			data[82372] <= 8'h10 ;
			data[82373] <= 8'h10 ;
			data[82374] <= 8'h10 ;
			data[82375] <= 8'h10 ;
			data[82376] <= 8'h10 ;
			data[82377] <= 8'h10 ;
			data[82378] <= 8'h10 ;
			data[82379] <= 8'h10 ;
			data[82380] <= 8'h10 ;
			data[82381] <= 8'h10 ;
			data[82382] <= 8'h10 ;
			data[82383] <= 8'h10 ;
			data[82384] <= 8'h10 ;
			data[82385] <= 8'h10 ;
			data[82386] <= 8'h10 ;
			data[82387] <= 8'h10 ;
			data[82388] <= 8'h10 ;
			data[82389] <= 8'h10 ;
			data[82390] <= 8'h10 ;
			data[82391] <= 8'h10 ;
			data[82392] <= 8'h10 ;
			data[82393] <= 8'h10 ;
			data[82394] <= 8'h10 ;
			data[82395] <= 8'h10 ;
			data[82396] <= 8'h10 ;
			data[82397] <= 8'h10 ;
			data[82398] <= 8'h10 ;
			data[82399] <= 8'h10 ;
			data[82400] <= 8'h10 ;
			data[82401] <= 8'h10 ;
			data[82402] <= 8'h10 ;
			data[82403] <= 8'h10 ;
			data[82404] <= 8'h10 ;
			data[82405] <= 8'h10 ;
			data[82406] <= 8'h10 ;
			data[82407] <= 8'h10 ;
			data[82408] <= 8'h10 ;
			data[82409] <= 8'h10 ;
			data[82410] <= 8'h10 ;
			data[82411] <= 8'h10 ;
			data[82412] <= 8'h10 ;
			data[82413] <= 8'h10 ;
			data[82414] <= 8'h10 ;
			data[82415] <= 8'h10 ;
			data[82416] <= 8'h10 ;
			data[82417] <= 8'h10 ;
			data[82418] <= 8'h10 ;
			data[82419] <= 8'h10 ;
			data[82420] <= 8'h10 ;
			data[82421] <= 8'h10 ;
			data[82422] <= 8'h10 ;
			data[82423] <= 8'h10 ;
			data[82424] <= 8'h10 ;
			data[82425] <= 8'h10 ;
			data[82426] <= 8'h10 ;
			data[82427] <= 8'h10 ;
			data[82428] <= 8'h10 ;
			data[82429] <= 8'h10 ;
			data[82430] <= 8'h10 ;
			data[82431] <= 8'h10 ;
			data[82432] <= 8'h10 ;
			data[82433] <= 8'h10 ;
			data[82434] <= 8'h10 ;
			data[82435] <= 8'h10 ;
			data[82436] <= 8'h10 ;
			data[82437] <= 8'h10 ;
			data[82438] <= 8'h10 ;
			data[82439] <= 8'h10 ;
			data[82440] <= 8'h10 ;
			data[82441] <= 8'h10 ;
			data[82442] <= 8'h10 ;
			data[82443] <= 8'h10 ;
			data[82444] <= 8'h10 ;
			data[82445] <= 8'h10 ;
			data[82446] <= 8'h10 ;
			data[82447] <= 8'h10 ;
			data[82448] <= 8'h10 ;
			data[82449] <= 8'h10 ;
			data[82450] <= 8'h10 ;
			data[82451] <= 8'h10 ;
			data[82452] <= 8'h10 ;
			data[82453] <= 8'h10 ;
			data[82454] <= 8'h10 ;
			data[82455] <= 8'h10 ;
			data[82456] <= 8'h10 ;
			data[82457] <= 8'h10 ;
			data[82458] <= 8'h10 ;
			data[82459] <= 8'h10 ;
			data[82460] <= 8'h10 ;
			data[82461] <= 8'h10 ;
			data[82462] <= 8'h10 ;
			data[82463] <= 8'h10 ;
			data[82464] <= 8'h10 ;
			data[82465] <= 8'h10 ;
			data[82466] <= 8'h10 ;
			data[82467] <= 8'h10 ;
			data[82468] <= 8'h10 ;
			data[82469] <= 8'h10 ;
			data[82470] <= 8'h10 ;
			data[82471] <= 8'h10 ;
			data[82472] <= 8'h10 ;
			data[82473] <= 8'h10 ;
			data[82474] <= 8'h10 ;
			data[82475] <= 8'h10 ;
			data[82476] <= 8'h10 ;
			data[82477] <= 8'h10 ;
			data[82478] <= 8'h10 ;
			data[82479] <= 8'h10 ;
			data[82480] <= 8'h10 ;
			data[82481] <= 8'h10 ;
			data[82482] <= 8'h10 ;
			data[82483] <= 8'h10 ;
			data[82484] <= 8'h10 ;
			data[82485] <= 8'h10 ;
			data[82486] <= 8'h10 ;
			data[82487] <= 8'h10 ;
			data[82488] <= 8'h10 ;
			data[82489] <= 8'h10 ;
			data[82490] <= 8'h10 ;
			data[82491] <= 8'h10 ;
			data[82492] <= 8'h10 ;
			data[82493] <= 8'h10 ;
			data[82494] <= 8'h10 ;
			data[82495] <= 8'h10 ;
			data[82496] <= 8'h10 ;
			data[82497] <= 8'h10 ;
			data[82498] <= 8'h10 ;
			data[82499] <= 8'h10 ;
			data[82500] <= 8'h10 ;
			data[82501] <= 8'h10 ;
			data[82502] <= 8'h10 ;
			data[82503] <= 8'h10 ;
			data[82504] <= 8'h10 ;
			data[82505] <= 8'h10 ;
			data[82506] <= 8'h10 ;
			data[82507] <= 8'h10 ;
			data[82508] <= 8'h10 ;
			data[82509] <= 8'h10 ;
			data[82510] <= 8'h10 ;
			data[82511] <= 8'h10 ;
			data[82512] <= 8'h10 ;
			data[82513] <= 8'h10 ;
			data[82514] <= 8'h10 ;
			data[82515] <= 8'h10 ;
			data[82516] <= 8'h10 ;
			data[82517] <= 8'h10 ;
			data[82518] <= 8'h10 ;
			data[82519] <= 8'h10 ;
			data[82520] <= 8'h10 ;
			data[82521] <= 8'h10 ;
			data[82522] <= 8'h10 ;
			data[82523] <= 8'h10 ;
			data[82524] <= 8'h10 ;
			data[82525] <= 8'h10 ;
			data[82526] <= 8'h10 ;
			data[82527] <= 8'h10 ;
			data[82528] <= 8'h10 ;
			data[82529] <= 8'h10 ;
			data[82530] <= 8'h10 ;
			data[82531] <= 8'h10 ;
			data[82532] <= 8'h10 ;
			data[82533] <= 8'h10 ;
			data[82534] <= 8'h10 ;
			data[82535] <= 8'h10 ;
			data[82536] <= 8'h10 ;
			data[82537] <= 8'h10 ;
			data[82538] <= 8'h10 ;
			data[82539] <= 8'h10 ;
			data[82540] <= 8'h10 ;
			data[82541] <= 8'h10 ;
			data[82542] <= 8'h10 ;
			data[82543] <= 8'h10 ;
			data[82544] <= 8'h10 ;
			data[82545] <= 8'h10 ;
			data[82546] <= 8'h10 ;
			data[82547] <= 8'h10 ;
			data[82548] <= 8'h10 ;
			data[82549] <= 8'h10 ;
			data[82550] <= 8'h10 ;
			data[82551] <= 8'h10 ;
			data[82552] <= 8'h10 ;
			data[82553] <= 8'h10 ;
			data[82554] <= 8'h10 ;
			data[82555] <= 8'h10 ;
			data[82556] <= 8'h10 ;
			data[82557] <= 8'h10 ;
			data[82558] <= 8'h10 ;
			data[82559] <= 8'h10 ;
			data[82560] <= 8'h10 ;
			data[82561] <= 8'h10 ;
			data[82562] <= 8'h10 ;
			data[82563] <= 8'h10 ;
			data[82564] <= 8'h10 ;
			data[82565] <= 8'h10 ;
			data[82566] <= 8'h10 ;
			data[82567] <= 8'h10 ;
			data[82568] <= 8'h10 ;
			data[82569] <= 8'h10 ;
			data[82570] <= 8'h10 ;
			data[82571] <= 8'h10 ;
			data[82572] <= 8'h10 ;
			data[82573] <= 8'h10 ;
			data[82574] <= 8'h10 ;
			data[82575] <= 8'h10 ;
			data[82576] <= 8'h10 ;
			data[82577] <= 8'h10 ;
			data[82578] <= 8'h10 ;
			data[82579] <= 8'h10 ;
			data[82580] <= 8'h10 ;
			data[82581] <= 8'h10 ;
			data[82582] <= 8'h10 ;
			data[82583] <= 8'h10 ;
			data[82584] <= 8'h10 ;
			data[82585] <= 8'h10 ;
			data[82586] <= 8'h10 ;
			data[82587] <= 8'h10 ;
			data[82588] <= 8'h10 ;
			data[82589] <= 8'h10 ;
			data[82590] <= 8'h10 ;
			data[82591] <= 8'h10 ;
			data[82592] <= 8'h10 ;
			data[82593] <= 8'h10 ;
			data[82594] <= 8'h10 ;
			data[82595] <= 8'h10 ;
			data[82596] <= 8'h10 ;
			data[82597] <= 8'h10 ;
			data[82598] <= 8'h10 ;
			data[82599] <= 8'h10 ;
			data[82600] <= 8'h10 ;
			data[82601] <= 8'h10 ;
			data[82602] <= 8'h10 ;
			data[82603] <= 8'h10 ;
			data[82604] <= 8'h10 ;
			data[82605] <= 8'h10 ;
			data[82606] <= 8'h10 ;
			data[82607] <= 8'h10 ;
			data[82608] <= 8'h10 ;
			data[82609] <= 8'h10 ;
			data[82610] <= 8'h10 ;
			data[82611] <= 8'h10 ;
			data[82612] <= 8'h10 ;
			data[82613] <= 8'h10 ;
			data[82614] <= 8'h10 ;
			data[82615] <= 8'h10 ;
			data[82616] <= 8'h10 ;
			data[82617] <= 8'h10 ;
			data[82618] <= 8'h10 ;
			data[82619] <= 8'h10 ;
			data[82620] <= 8'h10 ;
			data[82621] <= 8'h10 ;
			data[82622] <= 8'h10 ;
			data[82623] <= 8'h10 ;
			data[82624] <= 8'h10 ;
			data[82625] <= 8'h10 ;
			data[82626] <= 8'h10 ;
			data[82627] <= 8'h10 ;
			data[82628] <= 8'h10 ;
			data[82629] <= 8'h10 ;
			data[82630] <= 8'h10 ;
			data[82631] <= 8'h10 ;
			data[82632] <= 8'h10 ;
			data[82633] <= 8'h10 ;
			data[82634] <= 8'h10 ;
			data[82635] <= 8'h10 ;
			data[82636] <= 8'h10 ;
			data[82637] <= 8'h10 ;
			data[82638] <= 8'h10 ;
			data[82639] <= 8'h10 ;
			data[82640] <= 8'h10 ;
			data[82641] <= 8'h10 ;
			data[82642] <= 8'h10 ;
			data[82643] <= 8'h10 ;
			data[82644] <= 8'h10 ;
			data[82645] <= 8'h10 ;
			data[82646] <= 8'h10 ;
			data[82647] <= 8'h10 ;
			data[82648] <= 8'h10 ;
			data[82649] <= 8'h10 ;
			data[82650] <= 8'h10 ;
			data[82651] <= 8'h10 ;
			data[82652] <= 8'h10 ;
			data[82653] <= 8'h10 ;
			data[82654] <= 8'h10 ;
			data[82655] <= 8'h10 ;
			data[82656] <= 8'h10 ;
			data[82657] <= 8'h10 ;
			data[82658] <= 8'h10 ;
			data[82659] <= 8'h10 ;
			data[82660] <= 8'h10 ;
			data[82661] <= 8'h10 ;
			data[82662] <= 8'h10 ;
			data[82663] <= 8'h10 ;
			data[82664] <= 8'h10 ;
			data[82665] <= 8'h10 ;
			data[82666] <= 8'h10 ;
			data[82667] <= 8'h10 ;
			data[82668] <= 8'h10 ;
			data[82669] <= 8'h10 ;
			data[82670] <= 8'h10 ;
			data[82671] <= 8'h10 ;
			data[82672] <= 8'h10 ;
			data[82673] <= 8'h10 ;
			data[82674] <= 8'h10 ;
			data[82675] <= 8'h10 ;
			data[82676] <= 8'h10 ;
			data[82677] <= 8'h10 ;
			data[82678] <= 8'h10 ;
			data[82679] <= 8'h10 ;
			data[82680] <= 8'h10 ;
			data[82681] <= 8'h10 ;
			data[82682] <= 8'h10 ;
			data[82683] <= 8'h10 ;
			data[82684] <= 8'h10 ;
			data[82685] <= 8'h10 ;
			data[82686] <= 8'h10 ;
			data[82687] <= 8'h10 ;
			data[82688] <= 8'h10 ;
			data[82689] <= 8'h10 ;
			data[82690] <= 8'h10 ;
			data[82691] <= 8'h10 ;
			data[82692] <= 8'h10 ;
			data[82693] <= 8'h10 ;
			data[82694] <= 8'h10 ;
			data[82695] <= 8'h10 ;
			data[82696] <= 8'h10 ;
			data[82697] <= 8'h10 ;
			data[82698] <= 8'h10 ;
			data[82699] <= 8'h10 ;
			data[82700] <= 8'h10 ;
			data[82701] <= 8'h10 ;
			data[82702] <= 8'h10 ;
			data[82703] <= 8'h10 ;
			data[82704] <= 8'h10 ;
			data[82705] <= 8'h10 ;
			data[82706] <= 8'h10 ;
			data[82707] <= 8'h10 ;
			data[82708] <= 8'h10 ;
			data[82709] <= 8'h10 ;
			data[82710] <= 8'h10 ;
			data[82711] <= 8'h10 ;
			data[82712] <= 8'h10 ;
			data[82713] <= 8'h10 ;
			data[82714] <= 8'h10 ;
			data[82715] <= 8'h10 ;
			data[82716] <= 8'h10 ;
			data[82717] <= 8'h10 ;
			data[82718] <= 8'h10 ;
			data[82719] <= 8'h10 ;
			data[82720] <= 8'h10 ;
			data[82721] <= 8'h10 ;
			data[82722] <= 8'h10 ;
			data[82723] <= 8'h10 ;
			data[82724] <= 8'h10 ;
			data[82725] <= 8'h10 ;
			data[82726] <= 8'h10 ;
			data[82727] <= 8'h10 ;
			data[82728] <= 8'h10 ;
			data[82729] <= 8'h10 ;
			data[82730] <= 8'h10 ;
			data[82731] <= 8'h10 ;
			data[82732] <= 8'h10 ;
			data[82733] <= 8'h10 ;
			data[82734] <= 8'h10 ;
			data[82735] <= 8'h10 ;
			data[82736] <= 8'h10 ;
			data[82737] <= 8'h10 ;
			data[82738] <= 8'h10 ;
			data[82739] <= 8'h10 ;
			data[82740] <= 8'h10 ;
			data[82741] <= 8'h10 ;
			data[82742] <= 8'h10 ;
			data[82743] <= 8'h10 ;
			data[82744] <= 8'h10 ;
			data[82745] <= 8'h10 ;
			data[82746] <= 8'h10 ;
			data[82747] <= 8'h10 ;
			data[82748] <= 8'h10 ;
			data[82749] <= 8'h10 ;
			data[82750] <= 8'h10 ;
			data[82751] <= 8'h10 ;
			data[82752] <= 8'h10 ;
			data[82753] <= 8'h10 ;
			data[82754] <= 8'h10 ;
			data[82755] <= 8'h10 ;
			data[82756] <= 8'h10 ;
			data[82757] <= 8'h10 ;
			data[82758] <= 8'h10 ;
			data[82759] <= 8'h10 ;
			data[82760] <= 8'h10 ;
			data[82761] <= 8'h10 ;
			data[82762] <= 8'h10 ;
			data[82763] <= 8'h10 ;
			data[82764] <= 8'h10 ;
			data[82765] <= 8'h10 ;
			data[82766] <= 8'h10 ;
			data[82767] <= 8'h10 ;
			data[82768] <= 8'h10 ;
			data[82769] <= 8'h10 ;
			data[82770] <= 8'h10 ;
			data[82771] <= 8'h10 ;
			data[82772] <= 8'h10 ;
			data[82773] <= 8'h10 ;
			data[82774] <= 8'h10 ;
			data[82775] <= 8'h10 ;
			data[82776] <= 8'h10 ;
			data[82777] <= 8'h10 ;
			data[82778] <= 8'h10 ;
			data[82779] <= 8'h10 ;
			data[82780] <= 8'h10 ;
			data[82781] <= 8'h10 ;
			data[82782] <= 8'h10 ;
			data[82783] <= 8'h10 ;
			data[82784] <= 8'h10 ;
			data[82785] <= 8'h10 ;
			data[82786] <= 8'h10 ;
			data[82787] <= 8'h10 ;
			data[82788] <= 8'h10 ;
			data[82789] <= 8'h10 ;
			data[82790] <= 8'h10 ;
			data[82791] <= 8'h10 ;
			data[82792] <= 8'h10 ;
			data[82793] <= 8'h10 ;
			data[82794] <= 8'h10 ;
			data[82795] <= 8'h10 ;
			data[82796] <= 8'h10 ;
			data[82797] <= 8'h10 ;
			data[82798] <= 8'h10 ;
			data[82799] <= 8'h10 ;
			data[82800] <= 8'h10 ;
			data[82801] <= 8'h10 ;
			data[82802] <= 8'h10 ;
			data[82803] <= 8'h10 ;
			data[82804] <= 8'h10 ;
			data[82805] <= 8'h10 ;
			data[82806] <= 8'h10 ;
			data[82807] <= 8'h10 ;
			data[82808] <= 8'h10 ;
			data[82809] <= 8'h10 ;
			data[82810] <= 8'h10 ;
			data[82811] <= 8'h10 ;
			data[82812] <= 8'h10 ;
			data[82813] <= 8'h10 ;
			data[82814] <= 8'h10 ;
			data[82815] <= 8'h10 ;
			data[82816] <= 8'h10 ;
			data[82817] <= 8'h10 ;
			data[82818] <= 8'h10 ;
			data[82819] <= 8'h10 ;
			data[82820] <= 8'h10 ;
			data[82821] <= 8'h10 ;
			data[82822] <= 8'h10 ;
			data[82823] <= 8'h10 ;
			data[82824] <= 8'h10 ;
			data[82825] <= 8'h10 ;
			data[82826] <= 8'h10 ;
			data[82827] <= 8'h10 ;
			data[82828] <= 8'h10 ;
			data[82829] <= 8'h10 ;
			data[82830] <= 8'h10 ;
			data[82831] <= 8'h10 ;
			data[82832] <= 8'h10 ;
			data[82833] <= 8'h10 ;
			data[82834] <= 8'h10 ;
			data[82835] <= 8'h10 ;
			data[82836] <= 8'h10 ;
			data[82837] <= 8'h10 ;
			data[82838] <= 8'h10 ;
			data[82839] <= 8'h10 ;
			data[82840] <= 8'h10 ;
			data[82841] <= 8'h10 ;
			data[82842] <= 8'h10 ;
			data[82843] <= 8'h10 ;
			data[82844] <= 8'h10 ;
			data[82845] <= 8'h10 ;
			data[82846] <= 8'h10 ;
			data[82847] <= 8'h10 ;
			data[82848] <= 8'h10 ;
			data[82849] <= 8'h10 ;
			data[82850] <= 8'h10 ;
			data[82851] <= 8'h10 ;
			data[82852] <= 8'h10 ;
			data[82853] <= 8'h10 ;
			data[82854] <= 8'h10 ;
			data[82855] <= 8'h10 ;
			data[82856] <= 8'h10 ;
			data[82857] <= 8'h10 ;
			data[82858] <= 8'h10 ;
			data[82859] <= 8'h10 ;
			data[82860] <= 8'h10 ;
			data[82861] <= 8'h10 ;
			data[82862] <= 8'h10 ;
			data[82863] <= 8'h10 ;
			data[82864] <= 8'h10 ;
			data[82865] <= 8'h10 ;
			data[82866] <= 8'h10 ;
			data[82867] <= 8'h10 ;
			data[82868] <= 8'h10 ;
			data[82869] <= 8'h10 ;
			data[82870] <= 8'h10 ;
			data[82871] <= 8'h10 ;
			data[82872] <= 8'h10 ;
			data[82873] <= 8'h10 ;
			data[82874] <= 8'h10 ;
			data[82875] <= 8'h10 ;
			data[82876] <= 8'h10 ;
			data[82877] <= 8'h10 ;
			data[82878] <= 8'h10 ;
			data[82879] <= 8'h10 ;
			data[82880] <= 8'h10 ;
			data[82881] <= 8'h10 ;
			data[82882] <= 8'h10 ;
			data[82883] <= 8'h10 ;
			data[82884] <= 8'h10 ;
			data[82885] <= 8'h10 ;
			data[82886] <= 8'h10 ;
			data[82887] <= 8'h10 ;
			data[82888] <= 8'h10 ;
			data[82889] <= 8'h10 ;
			data[82890] <= 8'h10 ;
			data[82891] <= 8'h10 ;
			data[82892] <= 8'h10 ;
			data[82893] <= 8'h10 ;
			data[82894] <= 8'h10 ;
			data[82895] <= 8'h10 ;
			data[82896] <= 8'h10 ;
			data[82897] <= 8'h10 ;
			data[82898] <= 8'h10 ;
			data[82899] <= 8'h10 ;
			data[82900] <= 8'h10 ;
			data[82901] <= 8'h10 ;
			data[82902] <= 8'h10 ;
			data[82903] <= 8'h10 ;
			data[82904] <= 8'h10 ;
			data[82905] <= 8'h10 ;
			data[82906] <= 8'h10 ;
			data[82907] <= 8'h10 ;
			data[82908] <= 8'h10 ;
			data[82909] <= 8'h10 ;
			data[82910] <= 8'h10 ;
			data[82911] <= 8'h10 ;
			data[82912] <= 8'h10 ;
			data[82913] <= 8'h10 ;
			data[82914] <= 8'h10 ;
			data[82915] <= 8'h10 ;
			data[82916] <= 8'h10 ;
			data[82917] <= 8'h10 ;
			data[82918] <= 8'h10 ;
			data[82919] <= 8'h10 ;
			data[82920] <= 8'h10 ;
			data[82921] <= 8'h10 ;
			data[82922] <= 8'h10 ;
			data[82923] <= 8'h10 ;
			data[82924] <= 8'h10 ;
			data[82925] <= 8'h10 ;
			data[82926] <= 8'h10 ;
			data[82927] <= 8'h10 ;
			data[82928] <= 8'h10 ;
			data[82929] <= 8'h10 ;
			data[82930] <= 8'h10 ;
			data[82931] <= 8'h10 ;
			data[82932] <= 8'h10 ;
			data[82933] <= 8'h10 ;
			data[82934] <= 8'h10 ;
			data[82935] <= 8'h10 ;
			data[82936] <= 8'h10 ;
			data[82937] <= 8'h10 ;
			data[82938] <= 8'h10 ;
			data[82939] <= 8'h10 ;
			data[82940] <= 8'h10 ;
			data[82941] <= 8'h10 ;
			data[82942] <= 8'h10 ;
			data[82943] <= 8'h10 ;
			data[82944] <= 8'h10 ;
			data[82945] <= 8'h10 ;
			data[82946] <= 8'h10 ;
			data[82947] <= 8'h10 ;
			data[82948] <= 8'h10 ;
			data[82949] <= 8'h10 ;
			data[82950] <= 8'h10 ;
			data[82951] <= 8'h10 ;
			data[82952] <= 8'h10 ;
			data[82953] <= 8'h10 ;
			data[82954] <= 8'h10 ;
			data[82955] <= 8'h10 ;
			data[82956] <= 8'h10 ;
			data[82957] <= 8'h10 ;
			data[82958] <= 8'h10 ;
			data[82959] <= 8'h10 ;
			data[82960] <= 8'h10 ;
			data[82961] <= 8'h10 ;
			data[82962] <= 8'h10 ;
			data[82963] <= 8'h10 ;
			data[82964] <= 8'h10 ;
			data[82965] <= 8'h10 ;
			data[82966] <= 8'h10 ;
			data[82967] <= 8'h10 ;
			data[82968] <= 8'h10 ;
			data[82969] <= 8'h10 ;
			data[82970] <= 8'h10 ;
			data[82971] <= 8'h10 ;
			data[82972] <= 8'h10 ;
			data[82973] <= 8'h10 ;
			data[82974] <= 8'h10 ;
			data[82975] <= 8'h10 ;
			data[82976] <= 8'h10 ;
			data[82977] <= 8'h10 ;
			data[82978] <= 8'h10 ;
			data[82979] <= 8'h10 ;
			data[82980] <= 8'h10 ;
			data[82981] <= 8'h10 ;
			data[82982] <= 8'h10 ;
			data[82983] <= 8'h10 ;
			data[82984] <= 8'h10 ;
			data[82985] <= 8'h10 ;
			data[82986] <= 8'h10 ;
			data[82987] <= 8'h10 ;
			data[82988] <= 8'h10 ;
			data[82989] <= 8'h10 ;
			data[82990] <= 8'h10 ;
			data[82991] <= 8'h10 ;
			data[82992] <= 8'h10 ;
			data[82993] <= 8'h10 ;
			data[82994] <= 8'h10 ;
			data[82995] <= 8'h10 ;
			data[82996] <= 8'h10 ;
			data[82997] <= 8'h10 ;
			data[82998] <= 8'h10 ;
			data[82999] <= 8'h10 ;
			data[83000] <= 8'h10 ;
			data[83001] <= 8'h10 ;
			data[83002] <= 8'h10 ;
			data[83003] <= 8'h10 ;
			data[83004] <= 8'h10 ;
			data[83005] <= 8'h10 ;
			data[83006] <= 8'h10 ;
			data[83007] <= 8'h10 ;
			data[83008] <= 8'h10 ;
			data[83009] <= 8'h10 ;
			data[83010] <= 8'h10 ;
			data[83011] <= 8'h10 ;
			data[83012] <= 8'h10 ;
			data[83013] <= 8'h10 ;
			data[83014] <= 8'h10 ;
			data[83015] <= 8'h10 ;
			data[83016] <= 8'h10 ;
			data[83017] <= 8'h10 ;
			data[83018] <= 8'h10 ;
			data[83019] <= 8'h10 ;
			data[83020] <= 8'h10 ;
			data[83021] <= 8'h10 ;
			data[83022] <= 8'h10 ;
			data[83023] <= 8'h10 ;
			data[83024] <= 8'h10 ;
			data[83025] <= 8'h10 ;
			data[83026] <= 8'h10 ;
			data[83027] <= 8'h10 ;
			data[83028] <= 8'h10 ;
			data[83029] <= 8'h10 ;
			data[83030] <= 8'h10 ;
			data[83031] <= 8'h10 ;
			data[83032] <= 8'h10 ;
			data[83033] <= 8'h10 ;
			data[83034] <= 8'h10 ;
			data[83035] <= 8'h10 ;
			data[83036] <= 8'h10 ;
			data[83037] <= 8'h10 ;
			data[83038] <= 8'h10 ;
			data[83039] <= 8'h10 ;
			data[83040] <= 8'h10 ;
			data[83041] <= 8'h10 ;
			data[83042] <= 8'h10 ;
			data[83043] <= 8'h10 ;
			data[83044] <= 8'h10 ;
			data[83045] <= 8'h10 ;
			data[83046] <= 8'h10 ;
			data[83047] <= 8'h10 ;
			data[83048] <= 8'h10 ;
			data[83049] <= 8'h10 ;
			data[83050] <= 8'h10 ;
			data[83051] <= 8'h10 ;
			data[83052] <= 8'h10 ;
			data[83053] <= 8'h10 ;
			data[83054] <= 8'h10 ;
			data[83055] <= 8'h10 ;
			data[83056] <= 8'h10 ;
			data[83057] <= 8'h10 ;
			data[83058] <= 8'h10 ;
			data[83059] <= 8'h10 ;
			data[83060] <= 8'h10 ;
			data[83061] <= 8'h10 ;
			data[83062] <= 8'h10 ;
			data[83063] <= 8'h10 ;
			data[83064] <= 8'h10 ;
			data[83065] <= 8'h10 ;
			data[83066] <= 8'h10 ;
			data[83067] <= 8'h10 ;
			data[83068] <= 8'h10 ;
			data[83069] <= 8'h10 ;
			data[83070] <= 8'h10 ;
			data[83071] <= 8'h10 ;
			data[83072] <= 8'h10 ;
			data[83073] <= 8'h10 ;
			data[83074] <= 8'h10 ;
			data[83075] <= 8'h10 ;
			data[83076] <= 8'h10 ;
			data[83077] <= 8'h10 ;
			data[83078] <= 8'h10 ;
			data[83079] <= 8'h10 ;
			data[83080] <= 8'h10 ;
			data[83081] <= 8'h10 ;
			data[83082] <= 8'h10 ;
			data[83083] <= 8'h10 ;
			data[83084] <= 8'h10 ;
			data[83085] <= 8'h10 ;
			data[83086] <= 8'h10 ;
			data[83087] <= 8'h10 ;
			data[83088] <= 8'h10 ;
			data[83089] <= 8'h10 ;
			data[83090] <= 8'h10 ;
			data[83091] <= 8'h10 ;
			data[83092] <= 8'h10 ;
			data[83093] <= 8'h10 ;
			data[83094] <= 8'h10 ;
			data[83095] <= 8'h10 ;
			data[83096] <= 8'h10 ;
			data[83097] <= 8'h10 ;
			data[83098] <= 8'h10 ;
			data[83099] <= 8'h10 ;
			data[83100] <= 8'h10 ;
			data[83101] <= 8'h10 ;
			data[83102] <= 8'h10 ;
			data[83103] <= 8'h10 ;
			data[83104] <= 8'h10 ;
			data[83105] <= 8'h10 ;
			data[83106] <= 8'h10 ;
			data[83107] <= 8'h10 ;
			data[83108] <= 8'h10 ;
			data[83109] <= 8'h10 ;
			data[83110] <= 8'h10 ;
			data[83111] <= 8'h10 ;
			data[83112] <= 8'h10 ;
			data[83113] <= 8'h10 ;
			data[83114] <= 8'h10 ;
			data[83115] <= 8'h10 ;
			data[83116] <= 8'h10 ;
			data[83117] <= 8'h10 ;
			data[83118] <= 8'h10 ;
			data[83119] <= 8'h10 ;
			data[83120] <= 8'h10 ;
			data[83121] <= 8'h10 ;
			data[83122] <= 8'h10 ;
			data[83123] <= 8'h10 ;
			data[83124] <= 8'h10 ;
			data[83125] <= 8'h10 ;
			data[83126] <= 8'h10 ;
			data[83127] <= 8'h10 ;
			data[83128] <= 8'h10 ;
			data[83129] <= 8'h10 ;
			data[83130] <= 8'h10 ;
			data[83131] <= 8'h10 ;
			data[83132] <= 8'h10 ;
			data[83133] <= 8'h10 ;
			data[83134] <= 8'h10 ;
			data[83135] <= 8'h10 ;
			data[83136] <= 8'h10 ;
			data[83137] <= 8'h10 ;
			data[83138] <= 8'h10 ;
			data[83139] <= 8'h10 ;
			data[83140] <= 8'h10 ;
			data[83141] <= 8'h10 ;
			data[83142] <= 8'h10 ;
			data[83143] <= 8'h10 ;
			data[83144] <= 8'h10 ;
			data[83145] <= 8'h10 ;
			data[83146] <= 8'h10 ;
			data[83147] <= 8'h10 ;
			data[83148] <= 8'h10 ;
			data[83149] <= 8'h10 ;
			data[83150] <= 8'h10 ;
			data[83151] <= 8'h10 ;
			data[83152] <= 8'h10 ;
			data[83153] <= 8'h10 ;
			data[83154] <= 8'h10 ;
			data[83155] <= 8'h10 ;
			data[83156] <= 8'h10 ;
			data[83157] <= 8'h10 ;
			data[83158] <= 8'h10 ;
			data[83159] <= 8'h10 ;
			data[83160] <= 8'h10 ;
			data[83161] <= 8'h10 ;
			data[83162] <= 8'h10 ;
			data[83163] <= 8'h10 ;
			data[83164] <= 8'h10 ;
			data[83165] <= 8'h10 ;
			data[83166] <= 8'h10 ;
			data[83167] <= 8'h10 ;
			data[83168] <= 8'h10 ;
			data[83169] <= 8'h10 ;
			data[83170] <= 8'h10 ;
			data[83171] <= 8'h10 ;
			data[83172] <= 8'h10 ;
			data[83173] <= 8'h10 ;
			data[83174] <= 8'h10 ;
			data[83175] <= 8'h10 ;
			data[83176] <= 8'h10 ;
			data[83177] <= 8'h10 ;
			data[83178] <= 8'h10 ;
			data[83179] <= 8'h10 ;
			data[83180] <= 8'h10 ;
			data[83181] <= 8'h10 ;
			data[83182] <= 8'h10 ;
			data[83183] <= 8'h10 ;
			data[83184] <= 8'h10 ;
			data[83185] <= 8'h10 ;
			data[83186] <= 8'h10 ;
			data[83187] <= 8'h10 ;
			data[83188] <= 8'h10 ;
			data[83189] <= 8'h10 ;
			data[83190] <= 8'h10 ;
			data[83191] <= 8'h10 ;
			data[83192] <= 8'h10 ;
			data[83193] <= 8'h10 ;
			data[83194] <= 8'h10 ;
			data[83195] <= 8'h10 ;
			data[83196] <= 8'h10 ;
			data[83197] <= 8'h10 ;
			data[83198] <= 8'h10 ;
			data[83199] <= 8'h10 ;
			data[83200] <= 8'h10 ;
			data[83201] <= 8'h10 ;
			data[83202] <= 8'h10 ;
			data[83203] <= 8'h10 ;
			data[83204] <= 8'h10 ;
			data[83205] <= 8'h10 ;
			data[83206] <= 8'h10 ;
			data[83207] <= 8'h10 ;
			data[83208] <= 8'h10 ;
			data[83209] <= 8'h10 ;
			data[83210] <= 8'h10 ;
			data[83211] <= 8'h10 ;
			data[83212] <= 8'h10 ;
			data[83213] <= 8'h10 ;
			data[83214] <= 8'h10 ;
			data[83215] <= 8'h10 ;
			data[83216] <= 8'h10 ;
			data[83217] <= 8'h10 ;
			data[83218] <= 8'h10 ;
			data[83219] <= 8'h10 ;
			data[83220] <= 8'h10 ;
			data[83221] <= 8'h10 ;
			data[83222] <= 8'h10 ;
			data[83223] <= 8'h10 ;
			data[83224] <= 8'h10 ;
			data[83225] <= 8'h10 ;
			data[83226] <= 8'h10 ;
			data[83227] <= 8'h10 ;
			data[83228] <= 8'h10 ;
			data[83229] <= 8'h10 ;
			data[83230] <= 8'h10 ;
			data[83231] <= 8'h10 ;
			data[83232] <= 8'h10 ;
			data[83233] <= 8'h10 ;
			data[83234] <= 8'h10 ;
			data[83235] <= 8'h10 ;
			data[83236] <= 8'h10 ;
			data[83237] <= 8'h10 ;
			data[83238] <= 8'h10 ;
			data[83239] <= 8'h10 ;
			data[83240] <= 8'h10 ;
			data[83241] <= 8'h10 ;
			data[83242] <= 8'h10 ;
			data[83243] <= 8'h10 ;
			data[83244] <= 8'h10 ;
			data[83245] <= 8'h10 ;
			data[83246] <= 8'h10 ;
			data[83247] <= 8'h10 ;
			data[83248] <= 8'h10 ;
			data[83249] <= 8'h10 ;
			data[83250] <= 8'h10 ;
			data[83251] <= 8'h10 ;
			data[83252] <= 8'h10 ;
			data[83253] <= 8'h10 ;
			data[83254] <= 8'h10 ;
			data[83255] <= 8'h10 ;
			data[83256] <= 8'h10 ;
			data[83257] <= 8'h10 ;
			data[83258] <= 8'h10 ;
			data[83259] <= 8'h10 ;
			data[83260] <= 8'h10 ;
			data[83261] <= 8'h10 ;
			data[83262] <= 8'h10 ;
			data[83263] <= 8'h10 ;
			data[83264] <= 8'h10 ;
			data[83265] <= 8'h10 ;
			data[83266] <= 8'h10 ;
			data[83267] <= 8'h10 ;
			data[83268] <= 8'h10 ;
			data[83269] <= 8'h10 ;
			data[83270] <= 8'h10 ;
			data[83271] <= 8'h10 ;
			data[83272] <= 8'h10 ;
			data[83273] <= 8'h10 ;
			data[83274] <= 8'h10 ;
			data[83275] <= 8'h10 ;
			data[83276] <= 8'h10 ;
			data[83277] <= 8'h10 ;
			data[83278] <= 8'h10 ;
			data[83279] <= 8'h10 ;
			data[83280] <= 8'h10 ;
			data[83281] <= 8'h10 ;
			data[83282] <= 8'h10 ;
			data[83283] <= 8'h10 ;
			data[83284] <= 8'h10 ;
			data[83285] <= 8'h10 ;
			data[83286] <= 8'h10 ;
			data[83287] <= 8'h10 ;
			data[83288] <= 8'h10 ;
			data[83289] <= 8'h10 ;
			data[83290] <= 8'h10 ;
			data[83291] <= 8'h10 ;
			data[83292] <= 8'h10 ;
			data[83293] <= 8'h10 ;
			data[83294] <= 8'h10 ;
			data[83295] <= 8'h10 ;
			data[83296] <= 8'h10 ;
			data[83297] <= 8'h10 ;
			data[83298] <= 8'h10 ;
			data[83299] <= 8'h10 ;
			data[83300] <= 8'h10 ;
			data[83301] <= 8'h10 ;
			data[83302] <= 8'h10 ;
			data[83303] <= 8'h10 ;
			data[83304] <= 8'h10 ;
			data[83305] <= 8'h10 ;
			data[83306] <= 8'h10 ;
			data[83307] <= 8'h10 ;
			data[83308] <= 8'h10 ;
			data[83309] <= 8'h10 ;
			data[83310] <= 8'h10 ;
			data[83311] <= 8'h10 ;
			data[83312] <= 8'h10 ;
			data[83313] <= 8'h10 ;
			data[83314] <= 8'h10 ;
			data[83315] <= 8'h10 ;
			data[83316] <= 8'h10 ;
			data[83317] <= 8'h10 ;
			data[83318] <= 8'h10 ;
			data[83319] <= 8'h10 ;
			data[83320] <= 8'h10 ;
			data[83321] <= 8'h10 ;
			data[83322] <= 8'h10 ;
			data[83323] <= 8'h10 ;
			data[83324] <= 8'h10 ;
			data[83325] <= 8'h10 ;
			data[83326] <= 8'h10 ;
			data[83327] <= 8'h10 ;
			data[83328] <= 8'h10 ;
			data[83329] <= 8'h10 ;
			data[83330] <= 8'h10 ;
			data[83331] <= 8'h10 ;
			data[83332] <= 8'h10 ;
			data[83333] <= 8'h10 ;
			data[83334] <= 8'h10 ;
			data[83335] <= 8'h10 ;
			data[83336] <= 8'h10 ;
			data[83337] <= 8'h10 ;
			data[83338] <= 8'h10 ;
			data[83339] <= 8'h10 ;
			data[83340] <= 8'h10 ;
			data[83341] <= 8'h10 ;
			data[83342] <= 8'h10 ;
			data[83343] <= 8'h10 ;
			data[83344] <= 8'h10 ;
			data[83345] <= 8'h10 ;
			data[83346] <= 8'h10 ;
			data[83347] <= 8'h10 ;
			data[83348] <= 8'h10 ;
			data[83349] <= 8'h10 ;
			data[83350] <= 8'h10 ;
			data[83351] <= 8'h10 ;
			data[83352] <= 8'h10 ;
			data[83353] <= 8'h10 ;
			data[83354] <= 8'h10 ;
			data[83355] <= 8'h10 ;
			data[83356] <= 8'h10 ;
			data[83357] <= 8'h10 ;
			data[83358] <= 8'h10 ;
			data[83359] <= 8'h10 ;
			data[83360] <= 8'h10 ;
			data[83361] <= 8'h10 ;
			data[83362] <= 8'h10 ;
			data[83363] <= 8'h10 ;
			data[83364] <= 8'h10 ;
			data[83365] <= 8'h10 ;
			data[83366] <= 8'h10 ;
			data[83367] <= 8'h10 ;
			data[83368] <= 8'h10 ;
			data[83369] <= 8'h10 ;
			data[83370] <= 8'h10 ;
			data[83371] <= 8'h10 ;
			data[83372] <= 8'h10 ;
			data[83373] <= 8'h10 ;
			data[83374] <= 8'h10 ;
			data[83375] <= 8'h10 ;
			data[83376] <= 8'h10 ;
			data[83377] <= 8'h10 ;
			data[83378] <= 8'h10 ;
			data[83379] <= 8'h10 ;
			data[83380] <= 8'h10 ;
			data[83381] <= 8'h10 ;
			data[83382] <= 8'h10 ;
			data[83383] <= 8'h10 ;
			data[83384] <= 8'h10 ;
			data[83385] <= 8'h10 ;
			data[83386] <= 8'h10 ;
			data[83387] <= 8'h10 ;
			data[83388] <= 8'h10 ;
			data[83389] <= 8'h10 ;
			data[83390] <= 8'h10 ;
			data[83391] <= 8'h10 ;
			data[83392] <= 8'h10 ;
			data[83393] <= 8'h10 ;
			data[83394] <= 8'h10 ;
			data[83395] <= 8'h10 ;
			data[83396] <= 8'h10 ;
			data[83397] <= 8'h10 ;
			data[83398] <= 8'h10 ;
			data[83399] <= 8'h10 ;
			data[83400] <= 8'h10 ;
			data[83401] <= 8'h10 ;
			data[83402] <= 8'h10 ;
			data[83403] <= 8'h10 ;
			data[83404] <= 8'h10 ;
			data[83405] <= 8'h10 ;
			data[83406] <= 8'h10 ;
			data[83407] <= 8'h10 ;
			data[83408] <= 8'h10 ;
			data[83409] <= 8'h10 ;
			data[83410] <= 8'h10 ;
			data[83411] <= 8'h10 ;
			data[83412] <= 8'h10 ;
			data[83413] <= 8'h10 ;
			data[83414] <= 8'h10 ;
			data[83415] <= 8'h10 ;
			data[83416] <= 8'h10 ;
			data[83417] <= 8'h10 ;
			data[83418] <= 8'h10 ;
			data[83419] <= 8'h10 ;
			data[83420] <= 8'h10 ;
			data[83421] <= 8'h10 ;
			data[83422] <= 8'h10 ;
			data[83423] <= 8'h10 ;
			data[83424] <= 8'h10 ;
			data[83425] <= 8'h10 ;
			data[83426] <= 8'h10 ;
			data[83427] <= 8'h10 ;
			data[83428] <= 8'h10 ;
			data[83429] <= 8'h10 ;
			data[83430] <= 8'h10 ;
			data[83431] <= 8'h10 ;
			data[83432] <= 8'h10 ;
			data[83433] <= 8'h10 ;
			data[83434] <= 8'h10 ;
			data[83435] <= 8'h10 ;
			data[83436] <= 8'h10 ;
			data[83437] <= 8'h10 ;
			data[83438] <= 8'h10 ;
			data[83439] <= 8'h10 ;
			data[83440] <= 8'h10 ;
			data[83441] <= 8'h10 ;
			data[83442] <= 8'h10 ;
			data[83443] <= 8'h10 ;
			data[83444] <= 8'h10 ;
			data[83445] <= 8'h10 ;
			data[83446] <= 8'h10 ;
			data[83447] <= 8'h10 ;
			data[83448] <= 8'h10 ;
			data[83449] <= 8'h10 ;
			data[83450] <= 8'h10 ;
			data[83451] <= 8'h10 ;
			data[83452] <= 8'h10 ;
			data[83453] <= 8'h10 ;
			data[83454] <= 8'h10 ;
			data[83455] <= 8'h10 ;
			data[83456] <= 8'h10 ;
			data[83457] <= 8'h10 ;
			data[83458] <= 8'h10 ;
			data[83459] <= 8'h10 ;
			data[83460] <= 8'h10 ;
			data[83461] <= 8'h10 ;
			data[83462] <= 8'h10 ;
			data[83463] <= 8'h10 ;
			data[83464] <= 8'h10 ;
			data[83465] <= 8'h10 ;
			data[83466] <= 8'h10 ;
			data[83467] <= 8'h10 ;
			data[83468] <= 8'h10 ;
			data[83469] <= 8'h10 ;
			data[83470] <= 8'h10 ;
			data[83471] <= 8'h10 ;
			data[83472] <= 8'h10 ;
			data[83473] <= 8'h10 ;
			data[83474] <= 8'h10 ;
			data[83475] <= 8'h10 ;
			data[83476] <= 8'h10 ;
			data[83477] <= 8'h10 ;
			data[83478] <= 8'h10 ;
			data[83479] <= 8'h10 ;
			data[83480] <= 8'h10 ;
			data[83481] <= 8'h10 ;
			data[83482] <= 8'h10 ;
			data[83483] <= 8'h10 ;
			data[83484] <= 8'h10 ;
			data[83485] <= 8'h10 ;
			data[83486] <= 8'h10 ;
			data[83487] <= 8'h10 ;
			data[83488] <= 8'h10 ;
			data[83489] <= 8'h10 ;
			data[83490] <= 8'h10 ;
			data[83491] <= 8'h10 ;
			data[83492] <= 8'h10 ;
			data[83493] <= 8'h10 ;
			data[83494] <= 8'h10 ;
			data[83495] <= 8'h10 ;
			data[83496] <= 8'h10 ;
			data[83497] <= 8'h10 ;
			data[83498] <= 8'h10 ;
			data[83499] <= 8'h10 ;
			data[83500] <= 8'h10 ;
			data[83501] <= 8'h10 ;
			data[83502] <= 8'h10 ;
			data[83503] <= 8'h10 ;
			data[83504] <= 8'h10 ;
			data[83505] <= 8'h10 ;
			data[83506] <= 8'h10 ;
			data[83507] <= 8'h10 ;
			data[83508] <= 8'h10 ;
			data[83509] <= 8'h10 ;
			data[83510] <= 8'h10 ;
			data[83511] <= 8'h10 ;
			data[83512] <= 8'h10 ;
			data[83513] <= 8'h10 ;
			data[83514] <= 8'h10 ;
			data[83515] <= 8'h10 ;
			data[83516] <= 8'h10 ;
			data[83517] <= 8'h10 ;
			data[83518] <= 8'h10 ;
			data[83519] <= 8'h10 ;
			data[83520] <= 8'h10 ;
			data[83521] <= 8'h10 ;
			data[83522] <= 8'h10 ;
			data[83523] <= 8'h10 ;
			data[83524] <= 8'h10 ;
			data[83525] <= 8'h10 ;
			data[83526] <= 8'h10 ;
			data[83527] <= 8'h10 ;
			data[83528] <= 8'h10 ;
			data[83529] <= 8'h10 ;
			data[83530] <= 8'h10 ;
			data[83531] <= 8'h10 ;
			data[83532] <= 8'h10 ;
			data[83533] <= 8'h10 ;
			data[83534] <= 8'h10 ;
			data[83535] <= 8'h10 ;
			data[83536] <= 8'h10 ;
			data[83537] <= 8'h10 ;
			data[83538] <= 8'h10 ;
			data[83539] <= 8'h10 ;
			data[83540] <= 8'h10 ;
			data[83541] <= 8'h10 ;
			data[83542] <= 8'h10 ;
			data[83543] <= 8'h10 ;
			data[83544] <= 8'h10 ;
			data[83545] <= 8'h10 ;
			data[83546] <= 8'h10 ;
			data[83547] <= 8'h10 ;
			data[83548] <= 8'h10 ;
			data[83549] <= 8'h10 ;
			data[83550] <= 8'h10 ;
			data[83551] <= 8'h10 ;
			data[83552] <= 8'h10 ;
			data[83553] <= 8'h10 ;
			data[83554] <= 8'h10 ;
			data[83555] <= 8'h10 ;
			data[83556] <= 8'h10 ;
			data[83557] <= 8'h10 ;
			data[83558] <= 8'h10 ;
			data[83559] <= 8'h10 ;
			data[83560] <= 8'h10 ;
			data[83561] <= 8'h10 ;
			data[83562] <= 8'h10 ;
			data[83563] <= 8'h10 ;
			data[83564] <= 8'h10 ;
			data[83565] <= 8'h10 ;
			data[83566] <= 8'h10 ;
			data[83567] <= 8'h10 ;
			data[83568] <= 8'h10 ;
			data[83569] <= 8'h10 ;
			data[83570] <= 8'h10 ;
			data[83571] <= 8'h10 ;
			data[83572] <= 8'h10 ;
			data[83573] <= 8'h10 ;
			data[83574] <= 8'h10 ;
			data[83575] <= 8'h10 ;
			data[83576] <= 8'h10 ;
			data[83577] <= 8'h10 ;
			data[83578] <= 8'h10 ;
			data[83579] <= 8'h10 ;
			data[83580] <= 8'h10 ;
			data[83581] <= 8'h10 ;
			data[83582] <= 8'h10 ;
			data[83583] <= 8'h10 ;
			data[83584] <= 8'h10 ;
			data[83585] <= 8'h10 ;
			data[83586] <= 8'h10 ;
			data[83587] <= 8'h10 ;
			data[83588] <= 8'h10 ;
			data[83589] <= 8'h10 ;
			data[83590] <= 8'h10 ;
			data[83591] <= 8'h10 ;
			data[83592] <= 8'h10 ;
			data[83593] <= 8'h10 ;
			data[83594] <= 8'h10 ;
			data[83595] <= 8'h10 ;
			data[83596] <= 8'h10 ;
			data[83597] <= 8'h10 ;
			data[83598] <= 8'h10 ;
			data[83599] <= 8'h10 ;
			data[83600] <= 8'h10 ;
			data[83601] <= 8'h10 ;
			data[83602] <= 8'h10 ;
			data[83603] <= 8'h10 ;
			data[83604] <= 8'h10 ;
			data[83605] <= 8'h10 ;
			data[83606] <= 8'h10 ;
			data[83607] <= 8'h10 ;
			data[83608] <= 8'h10 ;
			data[83609] <= 8'h10 ;
			data[83610] <= 8'h10 ;
			data[83611] <= 8'h10 ;
			data[83612] <= 8'h10 ;
			data[83613] <= 8'h10 ;
			data[83614] <= 8'h10 ;
			data[83615] <= 8'h10 ;
			data[83616] <= 8'h10 ;
			data[83617] <= 8'h10 ;
			data[83618] <= 8'h10 ;
			data[83619] <= 8'h10 ;
			data[83620] <= 8'h10 ;
			data[83621] <= 8'h10 ;
			data[83622] <= 8'h10 ;
			data[83623] <= 8'h10 ;
			data[83624] <= 8'h10 ;
			data[83625] <= 8'h10 ;
			data[83626] <= 8'h10 ;
			data[83627] <= 8'h10 ;
			data[83628] <= 8'h10 ;
			data[83629] <= 8'h10 ;
			data[83630] <= 8'h10 ;
			data[83631] <= 8'h10 ;
			data[83632] <= 8'h10 ;
			data[83633] <= 8'h10 ;
			data[83634] <= 8'h10 ;
			data[83635] <= 8'h10 ;
			data[83636] <= 8'h10 ;
			data[83637] <= 8'h10 ;
			data[83638] <= 8'h10 ;
			data[83639] <= 8'h10 ;
			data[83640] <= 8'h10 ;
			data[83641] <= 8'h10 ;
			data[83642] <= 8'h10 ;
			data[83643] <= 8'h10 ;
			data[83644] <= 8'h10 ;
			data[83645] <= 8'h10 ;
			data[83646] <= 8'h10 ;
			data[83647] <= 8'h10 ;
			data[83648] <= 8'h10 ;
			data[83649] <= 8'h10 ;
			data[83650] <= 8'h10 ;
			data[83651] <= 8'h10 ;
			data[83652] <= 8'h10 ;
			data[83653] <= 8'h10 ;
			data[83654] <= 8'h10 ;
			data[83655] <= 8'h10 ;
			data[83656] <= 8'h10 ;
			data[83657] <= 8'h10 ;
			data[83658] <= 8'h10 ;
			data[83659] <= 8'h10 ;
			data[83660] <= 8'h10 ;
			data[83661] <= 8'h10 ;
			data[83662] <= 8'h10 ;
			data[83663] <= 8'h10 ;
			data[83664] <= 8'h10 ;
			data[83665] <= 8'h10 ;
			data[83666] <= 8'h10 ;
			data[83667] <= 8'h10 ;
			data[83668] <= 8'h10 ;
			data[83669] <= 8'h10 ;
			data[83670] <= 8'h10 ;
			data[83671] <= 8'h10 ;
			data[83672] <= 8'h10 ;
			data[83673] <= 8'h10 ;
			data[83674] <= 8'h10 ;
			data[83675] <= 8'h10 ;
			data[83676] <= 8'h10 ;
			data[83677] <= 8'h10 ;
			data[83678] <= 8'h10 ;
			data[83679] <= 8'h10 ;
			data[83680] <= 8'h10 ;
			data[83681] <= 8'h10 ;
			data[83682] <= 8'h10 ;
			data[83683] <= 8'h10 ;
			data[83684] <= 8'h10 ;
			data[83685] <= 8'h10 ;
			data[83686] <= 8'h10 ;
			data[83687] <= 8'h10 ;
			data[83688] <= 8'h10 ;
			data[83689] <= 8'h10 ;
			data[83690] <= 8'h10 ;
			data[83691] <= 8'h10 ;
			data[83692] <= 8'h10 ;
			data[83693] <= 8'h10 ;
			data[83694] <= 8'h10 ;
			data[83695] <= 8'h10 ;
			data[83696] <= 8'h10 ;
			data[83697] <= 8'h10 ;
			data[83698] <= 8'h10 ;
			data[83699] <= 8'h10 ;
			data[83700] <= 8'h10 ;
			data[83701] <= 8'h10 ;
			data[83702] <= 8'h10 ;
			data[83703] <= 8'h10 ;
			data[83704] <= 8'h10 ;
			data[83705] <= 8'h10 ;
			data[83706] <= 8'h10 ;
			data[83707] <= 8'h10 ;
			data[83708] <= 8'h10 ;
			data[83709] <= 8'h10 ;
			data[83710] <= 8'h10 ;
			data[83711] <= 8'h10 ;
			data[83712] <= 8'h10 ;
			data[83713] <= 8'h10 ;
			data[83714] <= 8'h10 ;
			data[83715] <= 8'h10 ;
			data[83716] <= 8'h10 ;
			data[83717] <= 8'h10 ;
			data[83718] <= 8'h10 ;
			data[83719] <= 8'h10 ;
			data[83720] <= 8'h10 ;
			data[83721] <= 8'h10 ;
			data[83722] <= 8'h10 ;
			data[83723] <= 8'h10 ;
			data[83724] <= 8'h10 ;
			data[83725] <= 8'h10 ;
			data[83726] <= 8'h10 ;
			data[83727] <= 8'h10 ;
			data[83728] <= 8'h10 ;
			data[83729] <= 8'h10 ;
			data[83730] <= 8'h10 ;
			data[83731] <= 8'h10 ;
			data[83732] <= 8'h10 ;
			data[83733] <= 8'h10 ;
			data[83734] <= 8'h10 ;
			data[83735] <= 8'h10 ;
			data[83736] <= 8'h10 ;
			data[83737] <= 8'h10 ;
			data[83738] <= 8'h10 ;
			data[83739] <= 8'h10 ;
			data[83740] <= 8'h10 ;
			data[83741] <= 8'h10 ;
			data[83742] <= 8'h10 ;
			data[83743] <= 8'h10 ;
			data[83744] <= 8'h10 ;
			data[83745] <= 8'h10 ;
			data[83746] <= 8'h10 ;
			data[83747] <= 8'h10 ;
			data[83748] <= 8'h10 ;
			data[83749] <= 8'h10 ;
			data[83750] <= 8'h10 ;
			data[83751] <= 8'h10 ;
			data[83752] <= 8'h10 ;
			data[83753] <= 8'h10 ;
			data[83754] <= 8'h10 ;
			data[83755] <= 8'h10 ;
			data[83756] <= 8'h10 ;
			data[83757] <= 8'h10 ;
			data[83758] <= 8'h10 ;
			data[83759] <= 8'h10 ;
			data[83760] <= 8'h10 ;
			data[83761] <= 8'h10 ;
			data[83762] <= 8'h10 ;
			data[83763] <= 8'h10 ;
			data[83764] <= 8'h10 ;
			data[83765] <= 8'h10 ;
			data[83766] <= 8'h10 ;
			data[83767] <= 8'h10 ;
			data[83768] <= 8'h10 ;
			data[83769] <= 8'h10 ;
			data[83770] <= 8'h10 ;
			data[83771] <= 8'h10 ;
			data[83772] <= 8'h10 ;
			data[83773] <= 8'h10 ;
			data[83774] <= 8'h10 ;
			data[83775] <= 8'h10 ;
			data[83776] <= 8'h10 ;
			data[83777] <= 8'h10 ;
			data[83778] <= 8'h10 ;
			data[83779] <= 8'h10 ;
			data[83780] <= 8'h10 ;
			data[83781] <= 8'h10 ;
			data[83782] <= 8'h10 ;
			data[83783] <= 8'h10 ;
			data[83784] <= 8'h10 ;
			data[83785] <= 8'h10 ;
			data[83786] <= 8'h10 ;
			data[83787] <= 8'h10 ;
			data[83788] <= 8'h10 ;
			data[83789] <= 8'h10 ;
			data[83790] <= 8'h10 ;
			data[83791] <= 8'h10 ;
			data[83792] <= 8'h10 ;
			data[83793] <= 8'h10 ;
			data[83794] <= 8'h10 ;
			data[83795] <= 8'h10 ;
			data[83796] <= 8'h10 ;
			data[83797] <= 8'h10 ;
			data[83798] <= 8'h10 ;
			data[83799] <= 8'h10 ;
			data[83800] <= 8'h10 ;
			data[83801] <= 8'h10 ;
			data[83802] <= 8'h10 ;
			data[83803] <= 8'h10 ;
			data[83804] <= 8'h10 ;
			data[83805] <= 8'h10 ;
			data[83806] <= 8'h10 ;
			data[83807] <= 8'h10 ;
			data[83808] <= 8'h10 ;
			data[83809] <= 8'h10 ;
			data[83810] <= 8'h10 ;
			data[83811] <= 8'h10 ;
			data[83812] <= 8'h10 ;
			data[83813] <= 8'h10 ;
			data[83814] <= 8'h10 ;
			data[83815] <= 8'h10 ;
			data[83816] <= 8'h10 ;
			data[83817] <= 8'h10 ;
			data[83818] <= 8'h10 ;
			data[83819] <= 8'h10 ;
			data[83820] <= 8'h10 ;
			data[83821] <= 8'h10 ;
			data[83822] <= 8'h10 ;
			data[83823] <= 8'h10 ;
			data[83824] <= 8'h10 ;
			data[83825] <= 8'h10 ;
			data[83826] <= 8'h10 ;
			data[83827] <= 8'h10 ;
			data[83828] <= 8'h10 ;
			data[83829] <= 8'h10 ;
			data[83830] <= 8'h10 ;
			data[83831] <= 8'h10 ;
			data[83832] <= 8'h10 ;
			data[83833] <= 8'h10 ;
			data[83834] <= 8'h10 ;
			data[83835] <= 8'h10 ;
			data[83836] <= 8'h10 ;
			data[83837] <= 8'h10 ;
			data[83838] <= 8'h10 ;
			data[83839] <= 8'h10 ;
			data[83840] <= 8'h10 ;
			data[83841] <= 8'h10 ;
			data[83842] <= 8'h10 ;
			data[83843] <= 8'h10 ;
			data[83844] <= 8'h10 ;
			data[83845] <= 8'h10 ;
			data[83846] <= 8'h10 ;
			data[83847] <= 8'h10 ;
			data[83848] <= 8'h10 ;
			data[83849] <= 8'h10 ;
			data[83850] <= 8'h10 ;
			data[83851] <= 8'h10 ;
			data[83852] <= 8'h10 ;
			data[83853] <= 8'h10 ;
			data[83854] <= 8'h10 ;
			data[83855] <= 8'h10 ;
			data[83856] <= 8'h10 ;
			data[83857] <= 8'h10 ;
			data[83858] <= 8'h10 ;
			data[83859] <= 8'h10 ;
			data[83860] <= 8'h10 ;
			data[83861] <= 8'h10 ;
			data[83862] <= 8'h10 ;
			data[83863] <= 8'h10 ;
			data[83864] <= 8'h10 ;
			data[83865] <= 8'h10 ;
			data[83866] <= 8'h10 ;
			data[83867] <= 8'h10 ;
			data[83868] <= 8'h10 ;
			data[83869] <= 8'h10 ;
			data[83870] <= 8'h10 ;
			data[83871] <= 8'h10 ;
			data[83872] <= 8'h10 ;
			data[83873] <= 8'h10 ;
			data[83874] <= 8'h10 ;
			data[83875] <= 8'h10 ;
			data[83876] <= 8'h10 ;
			data[83877] <= 8'h10 ;
			data[83878] <= 8'h10 ;
			data[83879] <= 8'h10 ;
			data[83880] <= 8'h10 ;
			data[83881] <= 8'h10 ;
			data[83882] <= 8'h10 ;
			data[83883] <= 8'h10 ;
			data[83884] <= 8'h10 ;
			data[83885] <= 8'h10 ;
			data[83886] <= 8'h10 ;
			data[83887] <= 8'h10 ;
			data[83888] <= 8'h10 ;
			data[83889] <= 8'h10 ;
			data[83890] <= 8'h10 ;
			data[83891] <= 8'h10 ;
			data[83892] <= 8'h10 ;
			data[83893] <= 8'h10 ;
			data[83894] <= 8'h10 ;
			data[83895] <= 8'h10 ;
			data[83896] <= 8'h10 ;
			data[83897] <= 8'h10 ;
			data[83898] <= 8'h10 ;
			data[83899] <= 8'h10 ;
			data[83900] <= 8'h10 ;
			data[83901] <= 8'h10 ;
			data[83902] <= 8'h10 ;
			data[83903] <= 8'h10 ;
			data[83904] <= 8'h10 ;
			data[83905] <= 8'h10 ;
			data[83906] <= 8'h10 ;
			data[83907] <= 8'h10 ;
			data[83908] <= 8'h10 ;
			data[83909] <= 8'h10 ;
			data[83910] <= 8'h10 ;
			data[83911] <= 8'h10 ;
			data[83912] <= 8'h10 ;
			data[83913] <= 8'h10 ;
			data[83914] <= 8'h10 ;
			data[83915] <= 8'h10 ;
			data[83916] <= 8'h10 ;
			data[83917] <= 8'h10 ;
			data[83918] <= 8'h10 ;
			data[83919] <= 8'h10 ;
			data[83920] <= 8'h10 ;
			data[83921] <= 8'h10 ;
			data[83922] <= 8'h10 ;
			data[83923] <= 8'h10 ;
			data[83924] <= 8'h10 ;
			data[83925] <= 8'h10 ;
			data[83926] <= 8'h10 ;
			data[83927] <= 8'h10 ;
			data[83928] <= 8'h10 ;
			data[83929] <= 8'h10 ;
			data[83930] <= 8'h10 ;
			data[83931] <= 8'h10 ;
			data[83932] <= 8'h10 ;
			data[83933] <= 8'h10 ;
			data[83934] <= 8'h10 ;
			data[83935] <= 8'h10 ;
			data[83936] <= 8'h10 ;
			data[83937] <= 8'h10 ;
			data[83938] <= 8'h10 ;
			data[83939] <= 8'h10 ;
			data[83940] <= 8'h10 ;
			data[83941] <= 8'h10 ;
			data[83942] <= 8'h10 ;
			data[83943] <= 8'h10 ;
			data[83944] <= 8'h10 ;
			data[83945] <= 8'h10 ;
			data[83946] <= 8'h10 ;
			data[83947] <= 8'h10 ;
			data[83948] <= 8'h10 ;
			data[83949] <= 8'h10 ;
			data[83950] <= 8'h10 ;
			data[83951] <= 8'h10 ;
			data[83952] <= 8'h10 ;
			data[83953] <= 8'h10 ;
			data[83954] <= 8'h10 ;
			data[83955] <= 8'h10 ;
			data[83956] <= 8'h10 ;
			data[83957] <= 8'h10 ;
			data[83958] <= 8'h10 ;
			data[83959] <= 8'h10 ;
			data[83960] <= 8'h10 ;
			data[83961] <= 8'h10 ;
			data[83962] <= 8'h10 ;
			data[83963] <= 8'h10 ;
			data[83964] <= 8'h10 ;
			data[83965] <= 8'h10 ;
			data[83966] <= 8'h10 ;
			data[83967] <= 8'h10 ;
			data[83968] <= 8'h10 ;
			data[83969] <= 8'h10 ;
			data[83970] <= 8'h10 ;
			data[83971] <= 8'h10 ;
			data[83972] <= 8'h10 ;
			data[83973] <= 8'h10 ;
			data[83974] <= 8'h10 ;
			data[83975] <= 8'h10 ;
			data[83976] <= 8'h10 ;
			data[83977] <= 8'h10 ;
			data[83978] <= 8'h10 ;
			data[83979] <= 8'h10 ;
			data[83980] <= 8'h10 ;
			data[83981] <= 8'h10 ;
			data[83982] <= 8'h10 ;
			data[83983] <= 8'h10 ;
			data[83984] <= 8'h10 ;
			data[83985] <= 8'h10 ;
			data[83986] <= 8'h10 ;
			data[83987] <= 8'h10 ;
			data[83988] <= 8'h10 ;
			data[83989] <= 8'h10 ;
			data[83990] <= 8'h10 ;
			data[83991] <= 8'h10 ;
			data[83992] <= 8'h10 ;
			data[83993] <= 8'h10 ;
			data[83994] <= 8'h10 ;
			data[83995] <= 8'h10 ;
			data[83996] <= 8'h10 ;
			data[83997] <= 8'h10 ;
			data[83998] <= 8'h10 ;
			data[83999] <= 8'h10 ;
			data[84000] <= 8'h10 ;
			data[84001] <= 8'h10 ;
			data[84002] <= 8'h10 ;
			data[84003] <= 8'h10 ;
			data[84004] <= 8'h10 ;
			data[84005] <= 8'h10 ;
			data[84006] <= 8'h10 ;
			data[84007] <= 8'h10 ;
			data[84008] <= 8'h10 ;
			data[84009] <= 8'h10 ;
			data[84010] <= 8'h10 ;
			data[84011] <= 8'h10 ;
			data[84012] <= 8'h10 ;
			data[84013] <= 8'h10 ;
			data[84014] <= 8'h10 ;
			data[84015] <= 8'h10 ;
			data[84016] <= 8'h10 ;
			data[84017] <= 8'h10 ;
			data[84018] <= 8'h10 ;
			data[84019] <= 8'h10 ;
			data[84020] <= 8'h10 ;
			data[84021] <= 8'h10 ;
			data[84022] <= 8'h10 ;
			data[84023] <= 8'h10 ;
			data[84024] <= 8'h10 ;
			data[84025] <= 8'h10 ;
			data[84026] <= 8'h10 ;
			data[84027] <= 8'h10 ;
			data[84028] <= 8'h10 ;
			data[84029] <= 8'h10 ;
			data[84030] <= 8'h10 ;
			data[84031] <= 8'h10 ;
			data[84032] <= 8'h10 ;
			data[84033] <= 8'h10 ;
			data[84034] <= 8'h10 ;
			data[84035] <= 8'h10 ;
			data[84036] <= 8'h10 ;
			data[84037] <= 8'h10 ;
			data[84038] <= 8'h10 ;
			data[84039] <= 8'h10 ;
			data[84040] <= 8'h10 ;
			data[84041] <= 8'h10 ;
			data[84042] <= 8'h10 ;
			data[84043] <= 8'h10 ;
			data[84044] <= 8'h10 ;
			data[84045] <= 8'h10 ;
			data[84046] <= 8'h10 ;
			data[84047] <= 8'h10 ;
			data[84048] <= 8'h10 ;
			data[84049] <= 8'h10 ;
			data[84050] <= 8'h10 ;
			data[84051] <= 8'h10 ;
			data[84052] <= 8'h10 ;
			data[84053] <= 8'h10 ;
			data[84054] <= 8'h10 ;
			data[84055] <= 8'h10 ;
			data[84056] <= 8'h10 ;
			data[84057] <= 8'h10 ;
			data[84058] <= 8'h10 ;
			data[84059] <= 8'h10 ;
			data[84060] <= 8'h10 ;
			data[84061] <= 8'h10 ;
			data[84062] <= 8'h10 ;
			data[84063] <= 8'h10 ;
			data[84064] <= 8'h10 ;
			data[84065] <= 8'h10 ;
			data[84066] <= 8'h10 ;
			data[84067] <= 8'h10 ;
			data[84068] <= 8'h10 ;
			data[84069] <= 8'h10 ;
			data[84070] <= 8'h10 ;
			data[84071] <= 8'h10 ;
			data[84072] <= 8'h10 ;
			data[84073] <= 8'h10 ;
			data[84074] <= 8'h10 ;
			data[84075] <= 8'h10 ;
			data[84076] <= 8'h10 ;
			data[84077] <= 8'h10 ;
			data[84078] <= 8'h10 ;
			data[84079] <= 8'h10 ;
			data[84080] <= 8'h10 ;
			data[84081] <= 8'h10 ;
			data[84082] <= 8'h10 ;
			data[84083] <= 8'h10 ;
			data[84084] <= 8'h10 ;
			data[84085] <= 8'h10 ;
			data[84086] <= 8'h10 ;
			data[84087] <= 8'h10 ;
			data[84088] <= 8'h10 ;
			data[84089] <= 8'h10 ;
			data[84090] <= 8'h10 ;
			data[84091] <= 8'h10 ;
			data[84092] <= 8'h10 ;
			data[84093] <= 8'h10 ;
			data[84094] <= 8'h10 ;
			data[84095] <= 8'h10 ;
			data[84096] <= 8'h10 ;
			data[84097] <= 8'h10 ;
			data[84098] <= 8'h10 ;
			data[84099] <= 8'h10 ;
			data[84100] <= 8'h10 ;
			data[84101] <= 8'h10 ;
			data[84102] <= 8'h10 ;
			data[84103] <= 8'h10 ;
			data[84104] <= 8'h10 ;
			data[84105] <= 8'h10 ;
			data[84106] <= 8'h10 ;
			data[84107] <= 8'h10 ;
			data[84108] <= 8'h10 ;
			data[84109] <= 8'h10 ;
			data[84110] <= 8'h10 ;
			data[84111] <= 8'h10 ;
			data[84112] <= 8'h10 ;
			data[84113] <= 8'h10 ;
			data[84114] <= 8'h10 ;
			data[84115] <= 8'h10 ;
			data[84116] <= 8'h10 ;
			data[84117] <= 8'h10 ;
			data[84118] <= 8'h10 ;
			data[84119] <= 8'h10 ;
			data[84120] <= 8'h10 ;
			data[84121] <= 8'h10 ;
			data[84122] <= 8'h10 ;
			data[84123] <= 8'h10 ;
			data[84124] <= 8'h10 ;
			data[84125] <= 8'h10 ;
			data[84126] <= 8'h10 ;
			data[84127] <= 8'h10 ;
			data[84128] <= 8'h10 ;
			data[84129] <= 8'h10 ;
			data[84130] <= 8'h10 ;
			data[84131] <= 8'h10 ;
			data[84132] <= 8'h10 ;
			data[84133] <= 8'h10 ;
			data[84134] <= 8'h10 ;
			data[84135] <= 8'h10 ;
			data[84136] <= 8'h10 ;
			data[84137] <= 8'h10 ;
			data[84138] <= 8'h10 ;
			data[84139] <= 8'h10 ;
			data[84140] <= 8'h10 ;
			data[84141] <= 8'h10 ;
			data[84142] <= 8'h10 ;
			data[84143] <= 8'h10 ;
			data[84144] <= 8'h10 ;
			data[84145] <= 8'h10 ;
			data[84146] <= 8'h10 ;
			data[84147] <= 8'h10 ;
			data[84148] <= 8'h10 ;
			data[84149] <= 8'h10 ;
			data[84150] <= 8'h10 ;
			data[84151] <= 8'h10 ;
			data[84152] <= 8'h10 ;
			data[84153] <= 8'h10 ;
			data[84154] <= 8'h10 ;
			data[84155] <= 8'h10 ;
			data[84156] <= 8'h10 ;
			data[84157] <= 8'h10 ;
			data[84158] <= 8'h10 ;
			data[84159] <= 8'h10 ;
			data[84160] <= 8'h10 ;
			data[84161] <= 8'h10 ;
			data[84162] <= 8'h10 ;
			data[84163] <= 8'h10 ;
			data[84164] <= 8'h10 ;
			data[84165] <= 8'h10 ;
			data[84166] <= 8'h10 ;
			data[84167] <= 8'h10 ;
			data[84168] <= 8'h10 ;
			data[84169] <= 8'h10 ;
			data[84170] <= 8'h10 ;
			data[84171] <= 8'h10 ;
			data[84172] <= 8'h10 ;
			data[84173] <= 8'h10 ;
			data[84174] <= 8'h10 ;
			data[84175] <= 8'h10 ;
			data[84176] <= 8'h10 ;
			data[84177] <= 8'h10 ;
			data[84178] <= 8'h10 ;
			data[84179] <= 8'h10 ;
			data[84180] <= 8'h10 ;
			data[84181] <= 8'h10 ;
			data[84182] <= 8'h10 ;
			data[84183] <= 8'h10 ;
			data[84184] <= 8'h10 ;
			data[84185] <= 8'h10 ;
			data[84186] <= 8'h10 ;
			data[84187] <= 8'h10 ;
			data[84188] <= 8'h10 ;
			data[84189] <= 8'h10 ;
			data[84190] <= 8'h10 ;
			data[84191] <= 8'h10 ;
			data[84192] <= 8'h10 ;
			data[84193] <= 8'h10 ;
			data[84194] <= 8'h10 ;
			data[84195] <= 8'h10 ;
			data[84196] <= 8'h10 ;
			data[84197] <= 8'h10 ;
			data[84198] <= 8'h10 ;
			data[84199] <= 8'h10 ;
			data[84200] <= 8'h10 ;
			data[84201] <= 8'h10 ;
			data[84202] <= 8'h10 ;
			data[84203] <= 8'h10 ;
			data[84204] <= 8'h10 ;
			data[84205] <= 8'h10 ;
			data[84206] <= 8'h10 ;
			data[84207] <= 8'h10 ;
			data[84208] <= 8'h10 ;
			data[84209] <= 8'h10 ;
			data[84210] <= 8'h10 ;
			data[84211] <= 8'h10 ;
			data[84212] <= 8'h10 ;
			data[84213] <= 8'h10 ;
			data[84214] <= 8'h10 ;
			data[84215] <= 8'h10 ;
			data[84216] <= 8'h10 ;
			data[84217] <= 8'h10 ;
			data[84218] <= 8'h10 ;
			data[84219] <= 8'h10 ;
			data[84220] <= 8'h10 ;
			data[84221] <= 8'h10 ;
			data[84222] <= 8'h10 ;
			data[84223] <= 8'h10 ;
			data[84224] <= 8'h10 ;
			data[84225] <= 8'h10 ;
			data[84226] <= 8'h10 ;
			data[84227] <= 8'h10 ;
			data[84228] <= 8'h10 ;
			data[84229] <= 8'h10 ;
			data[84230] <= 8'h10 ;
			data[84231] <= 8'h10 ;
			data[84232] <= 8'h10 ;
			data[84233] <= 8'h10 ;
			data[84234] <= 8'h10 ;
			data[84235] <= 8'h10 ;
			data[84236] <= 8'h10 ;
			data[84237] <= 8'h10 ;
			data[84238] <= 8'h10 ;
			data[84239] <= 8'h10 ;
			data[84240] <= 8'h10 ;
			data[84241] <= 8'h10 ;
			data[84242] <= 8'h10 ;
			data[84243] <= 8'h10 ;
			data[84244] <= 8'h10 ;
			data[84245] <= 8'h10 ;
			data[84246] <= 8'h10 ;
			data[84247] <= 8'h10 ;
			data[84248] <= 8'h10 ;
			data[84249] <= 8'h10 ;
			data[84250] <= 8'h10 ;
			data[84251] <= 8'h10 ;
			data[84252] <= 8'h10 ;
			data[84253] <= 8'h10 ;
			data[84254] <= 8'h10 ;
			data[84255] <= 8'h10 ;
			data[84256] <= 8'h10 ;
			data[84257] <= 8'h10 ;
			data[84258] <= 8'h10 ;
			data[84259] <= 8'h10 ;
			data[84260] <= 8'h10 ;
			data[84261] <= 8'h10 ;
			data[84262] <= 8'h10 ;
			data[84263] <= 8'h10 ;
			data[84264] <= 8'h10 ;
			data[84265] <= 8'h10 ;
			data[84266] <= 8'h10 ;
			data[84267] <= 8'h10 ;
			data[84268] <= 8'h10 ;
			data[84269] <= 8'h10 ;
			data[84270] <= 8'h10 ;
			data[84271] <= 8'h10 ;
			data[84272] <= 8'h10 ;
			data[84273] <= 8'h10 ;
			data[84274] <= 8'h10 ;
			data[84275] <= 8'h10 ;
			data[84276] <= 8'h10 ;
			data[84277] <= 8'h10 ;
			data[84278] <= 8'h10 ;
			data[84279] <= 8'h10 ;
			data[84280] <= 8'h10 ;
			data[84281] <= 8'h10 ;
			data[84282] <= 8'h10 ;
			data[84283] <= 8'h10 ;
			data[84284] <= 8'h10 ;
			data[84285] <= 8'h10 ;
			data[84286] <= 8'h10 ;
			data[84287] <= 8'h10 ;
			data[84288] <= 8'h10 ;
			data[84289] <= 8'h10 ;
			data[84290] <= 8'h10 ;
			data[84291] <= 8'h10 ;
			data[84292] <= 8'h10 ;
			data[84293] <= 8'h10 ;
			data[84294] <= 8'h10 ;
			data[84295] <= 8'h10 ;
			data[84296] <= 8'h10 ;
			data[84297] <= 8'h10 ;
			data[84298] <= 8'h10 ;
			data[84299] <= 8'h10 ;
			data[84300] <= 8'h10 ;
			data[84301] <= 8'h10 ;
			data[84302] <= 8'h10 ;
			data[84303] <= 8'h10 ;
			data[84304] <= 8'h10 ;
			data[84305] <= 8'h10 ;
			data[84306] <= 8'h10 ;
			data[84307] <= 8'h10 ;
			data[84308] <= 8'h10 ;
			data[84309] <= 8'h10 ;
			data[84310] <= 8'h10 ;
			data[84311] <= 8'h10 ;
			data[84312] <= 8'h10 ;
			data[84313] <= 8'h10 ;
			data[84314] <= 8'h10 ;
			data[84315] <= 8'h10 ;
			data[84316] <= 8'h10 ;
			data[84317] <= 8'h10 ;
			data[84318] <= 8'h10 ;
			data[84319] <= 8'h10 ;
			data[84320] <= 8'h10 ;
			data[84321] <= 8'h10 ;
			data[84322] <= 8'h10 ;
			data[84323] <= 8'h10 ;
			data[84324] <= 8'h10 ;
			data[84325] <= 8'h10 ;
			data[84326] <= 8'h10 ;
			data[84327] <= 8'h10 ;
			data[84328] <= 8'h10 ;
			data[84329] <= 8'h10 ;
			data[84330] <= 8'h10 ;
			data[84331] <= 8'h10 ;
			data[84332] <= 8'h10 ;
			data[84333] <= 8'h10 ;
			data[84334] <= 8'h10 ;
			data[84335] <= 8'h10 ;
			data[84336] <= 8'h10 ;
			data[84337] <= 8'h10 ;
			data[84338] <= 8'h10 ;
			data[84339] <= 8'h10 ;
			data[84340] <= 8'h10 ;
			data[84341] <= 8'h10 ;
			data[84342] <= 8'h10 ;
			data[84343] <= 8'h10 ;
			data[84344] <= 8'h10 ;
			data[84345] <= 8'h10 ;
			data[84346] <= 8'h10 ;
			data[84347] <= 8'h10 ;
			data[84348] <= 8'h10 ;
			data[84349] <= 8'h10 ;
			data[84350] <= 8'h10 ;
			data[84351] <= 8'h10 ;
			data[84352] <= 8'h10 ;
			data[84353] <= 8'h10 ;
			data[84354] <= 8'h10 ;
			data[84355] <= 8'h10 ;
			data[84356] <= 8'h10 ;
			data[84357] <= 8'h10 ;
			data[84358] <= 8'h10 ;
			data[84359] <= 8'h10 ;
			data[84360] <= 8'h10 ;
			data[84361] <= 8'h10 ;
			data[84362] <= 8'h10 ;
			data[84363] <= 8'h10 ;
			data[84364] <= 8'h10 ;
			data[84365] <= 8'h10 ;
			data[84366] <= 8'h10 ;
			data[84367] <= 8'h10 ;
			data[84368] <= 8'h10 ;
			data[84369] <= 8'h10 ;
			data[84370] <= 8'h10 ;
			data[84371] <= 8'h10 ;
			data[84372] <= 8'h10 ;
			data[84373] <= 8'h10 ;
			data[84374] <= 8'h10 ;
			data[84375] <= 8'h10 ;
			data[84376] <= 8'h10 ;
			data[84377] <= 8'h10 ;
			data[84378] <= 8'h10 ;
			data[84379] <= 8'h10 ;
			data[84380] <= 8'h10 ;
			data[84381] <= 8'h10 ;
			data[84382] <= 8'h10 ;
			data[84383] <= 8'h10 ;
			data[84384] <= 8'h10 ;
			data[84385] <= 8'h10 ;
			data[84386] <= 8'h10 ;
			data[84387] <= 8'h10 ;
			data[84388] <= 8'h10 ;
			data[84389] <= 8'h10 ;
			data[84390] <= 8'h10 ;
			data[84391] <= 8'h10 ;
			data[84392] <= 8'h10 ;
			data[84393] <= 8'h10 ;
			data[84394] <= 8'h10 ;
			data[84395] <= 8'h10 ;
			data[84396] <= 8'h10 ;
			data[84397] <= 8'h10 ;
			data[84398] <= 8'h10 ;
			data[84399] <= 8'h10 ;
			data[84400] <= 8'h10 ;
			data[84401] <= 8'h10 ;
			data[84402] <= 8'h10 ;
			data[84403] <= 8'h10 ;
			data[84404] <= 8'h10 ;
			data[84405] <= 8'h10 ;
			data[84406] <= 8'h10 ;
			data[84407] <= 8'h10 ;
			data[84408] <= 8'h10 ;
			data[84409] <= 8'h10 ;
			data[84410] <= 8'h10 ;
			data[84411] <= 8'h10 ;
			data[84412] <= 8'h10 ;
			data[84413] <= 8'h10 ;
			data[84414] <= 8'h10 ;
			data[84415] <= 8'h10 ;
			data[84416] <= 8'h10 ;
			data[84417] <= 8'h10 ;
			data[84418] <= 8'h10 ;
			data[84419] <= 8'h10 ;
			data[84420] <= 8'h10 ;
			data[84421] <= 8'h10 ;
			data[84422] <= 8'h10 ;
			data[84423] <= 8'h10 ;
			data[84424] <= 8'h10 ;
			data[84425] <= 8'h10 ;
			data[84426] <= 8'h10 ;
			data[84427] <= 8'h10 ;
			data[84428] <= 8'h10 ;
			data[84429] <= 8'h10 ;
			data[84430] <= 8'h10 ;
			data[84431] <= 8'h10 ;
			data[84432] <= 8'h10 ;
			data[84433] <= 8'h10 ;
			data[84434] <= 8'h10 ;
			data[84435] <= 8'h10 ;
			data[84436] <= 8'h10 ;
			data[84437] <= 8'h10 ;
			data[84438] <= 8'h10 ;
			data[84439] <= 8'h10 ;
			data[84440] <= 8'h10 ;
			data[84441] <= 8'h10 ;
			data[84442] <= 8'h10 ;
			data[84443] <= 8'h10 ;
			data[84444] <= 8'h10 ;
			data[84445] <= 8'h10 ;
			data[84446] <= 8'h10 ;
			data[84447] <= 8'h10 ;
			data[84448] <= 8'h10 ;
			data[84449] <= 8'h10 ;
			data[84450] <= 8'h10 ;
			data[84451] <= 8'h10 ;
			data[84452] <= 8'h10 ;
			data[84453] <= 8'h10 ;
			data[84454] <= 8'h10 ;
			data[84455] <= 8'h10 ;
			data[84456] <= 8'h10 ;
			data[84457] <= 8'h10 ;
			data[84458] <= 8'h10 ;
			data[84459] <= 8'h10 ;
			data[84460] <= 8'h10 ;
			data[84461] <= 8'h10 ;
			data[84462] <= 8'h10 ;
			data[84463] <= 8'h10 ;
			data[84464] <= 8'h10 ;
			data[84465] <= 8'h10 ;
			data[84466] <= 8'h10 ;
			data[84467] <= 8'h10 ;
			data[84468] <= 8'h10 ;
			data[84469] <= 8'h10 ;
			data[84470] <= 8'h10 ;
			data[84471] <= 8'h10 ;
			data[84472] <= 8'h10 ;
			data[84473] <= 8'h10 ;
			data[84474] <= 8'h10 ;
			data[84475] <= 8'h10 ;
			data[84476] <= 8'h10 ;
			data[84477] <= 8'h10 ;
			data[84478] <= 8'h10 ;
			data[84479] <= 8'h10 ;
			data[84480] <= 8'h10 ;
			data[84481] <= 8'h10 ;
			data[84482] <= 8'h10 ;
			data[84483] <= 8'h10 ;
			data[84484] <= 8'h10 ;
			data[84485] <= 8'h10 ;
			data[84486] <= 8'h10 ;
			data[84487] <= 8'h10 ;
			data[84488] <= 8'h10 ;
			data[84489] <= 8'h10 ;
			data[84490] <= 8'h10 ;
			data[84491] <= 8'h10 ;
			data[84492] <= 8'h10 ;
			data[84493] <= 8'h10 ;
			data[84494] <= 8'h10 ;
			data[84495] <= 8'h10 ;
			data[84496] <= 8'h10 ;
			data[84497] <= 8'h10 ;
			data[84498] <= 8'h10 ;
			data[84499] <= 8'h10 ;
			data[84500] <= 8'h10 ;
			data[84501] <= 8'h10 ;
			data[84502] <= 8'h10 ;
			data[84503] <= 8'h10 ;
			data[84504] <= 8'h10 ;
			data[84505] <= 8'h10 ;
			data[84506] <= 8'h10 ;
			data[84507] <= 8'h10 ;
			data[84508] <= 8'h10 ;
			data[84509] <= 8'h10 ;
			data[84510] <= 8'h10 ;
			data[84511] <= 8'h10 ;
			data[84512] <= 8'h10 ;
			data[84513] <= 8'h10 ;
			data[84514] <= 8'h10 ;
			data[84515] <= 8'h10 ;
			data[84516] <= 8'h10 ;
			data[84517] <= 8'h10 ;
			data[84518] <= 8'h10 ;
			data[84519] <= 8'h10 ;
			data[84520] <= 8'h10 ;
			data[84521] <= 8'h10 ;
			data[84522] <= 8'h10 ;
			data[84523] <= 8'h10 ;
			data[84524] <= 8'h10 ;
			data[84525] <= 8'h10 ;
			data[84526] <= 8'h10 ;
			data[84527] <= 8'h10 ;
			data[84528] <= 8'h10 ;
			data[84529] <= 8'h10 ;
			data[84530] <= 8'h10 ;
			data[84531] <= 8'h10 ;
			data[84532] <= 8'h10 ;
			data[84533] <= 8'h10 ;
			data[84534] <= 8'h10 ;
			data[84535] <= 8'h10 ;
			data[84536] <= 8'h10 ;
			data[84537] <= 8'h10 ;
			data[84538] <= 8'h10 ;
			data[84539] <= 8'h10 ;
			data[84540] <= 8'h10 ;
			data[84541] <= 8'h10 ;
			data[84542] <= 8'h10 ;
			data[84543] <= 8'h10 ;
			data[84544] <= 8'h10 ;
			data[84545] <= 8'h10 ;
			data[84546] <= 8'h10 ;
			data[84547] <= 8'h10 ;
			data[84548] <= 8'h10 ;
			data[84549] <= 8'h10 ;
			data[84550] <= 8'h10 ;
			data[84551] <= 8'h10 ;
			data[84552] <= 8'h10 ;
			data[84553] <= 8'h10 ;
			data[84554] <= 8'h10 ;
			data[84555] <= 8'h10 ;
			data[84556] <= 8'h10 ;
			data[84557] <= 8'h10 ;
			data[84558] <= 8'h10 ;
			data[84559] <= 8'h10 ;
			data[84560] <= 8'h10 ;
			data[84561] <= 8'h10 ;
			data[84562] <= 8'h10 ;
			data[84563] <= 8'h10 ;
			data[84564] <= 8'h10 ;
			data[84565] <= 8'h10 ;
			data[84566] <= 8'h10 ;
			data[84567] <= 8'h10 ;
			data[84568] <= 8'h10 ;
			data[84569] <= 8'h10 ;
			data[84570] <= 8'h10 ;
			data[84571] <= 8'h10 ;
			data[84572] <= 8'h10 ;
			data[84573] <= 8'h10 ;
			data[84574] <= 8'h10 ;
			data[84575] <= 8'h10 ;
			data[84576] <= 8'h10 ;
			data[84577] <= 8'h10 ;
			data[84578] <= 8'h10 ;
			data[84579] <= 8'h10 ;
			data[84580] <= 8'h10 ;
			data[84581] <= 8'h10 ;
			data[84582] <= 8'h10 ;
			data[84583] <= 8'h10 ;
			data[84584] <= 8'h10 ;
			data[84585] <= 8'h10 ;
			data[84586] <= 8'h10 ;
			data[84587] <= 8'h10 ;
			data[84588] <= 8'h10 ;
			data[84589] <= 8'h10 ;
			data[84590] <= 8'h10 ;
			data[84591] <= 8'h10 ;
			data[84592] <= 8'h10 ;
			data[84593] <= 8'h10 ;
			data[84594] <= 8'h10 ;
			data[84595] <= 8'h10 ;
			data[84596] <= 8'h10 ;
			data[84597] <= 8'h10 ;
			data[84598] <= 8'h10 ;
			data[84599] <= 8'h10 ;
			data[84600] <= 8'h10 ;
			data[84601] <= 8'h10 ;
			data[84602] <= 8'h10 ;
			data[84603] <= 8'h10 ;
			data[84604] <= 8'h10 ;
			data[84605] <= 8'h10 ;
			data[84606] <= 8'h10 ;
			data[84607] <= 8'h10 ;
			data[84608] <= 8'h10 ;
			data[84609] <= 8'h10 ;
			data[84610] <= 8'h10 ;
			data[84611] <= 8'h10 ;
			data[84612] <= 8'h10 ;
			data[84613] <= 8'h10 ;
			data[84614] <= 8'h10 ;
			data[84615] <= 8'h10 ;
			data[84616] <= 8'h10 ;
			data[84617] <= 8'h10 ;
			data[84618] <= 8'h10 ;
			data[84619] <= 8'h10 ;
			data[84620] <= 8'h10 ;
			data[84621] <= 8'h10 ;
			data[84622] <= 8'h10 ;
			data[84623] <= 8'h10 ;
			data[84624] <= 8'h10 ;
			data[84625] <= 8'h10 ;
			data[84626] <= 8'h10 ;
			data[84627] <= 8'h10 ;
			data[84628] <= 8'h10 ;
			data[84629] <= 8'h10 ;
			data[84630] <= 8'h10 ;
			data[84631] <= 8'h10 ;
			data[84632] <= 8'h10 ;
			data[84633] <= 8'h10 ;
			data[84634] <= 8'h10 ;
			data[84635] <= 8'h10 ;
			data[84636] <= 8'h10 ;
			data[84637] <= 8'h10 ;
			data[84638] <= 8'h10 ;
			data[84639] <= 8'h10 ;
			data[84640] <= 8'h10 ;
			data[84641] <= 8'h10 ;
			data[84642] <= 8'h10 ;
			data[84643] <= 8'h10 ;
			data[84644] <= 8'h10 ;
			data[84645] <= 8'h10 ;
			data[84646] <= 8'h10 ;
			data[84647] <= 8'h10 ;
			data[84648] <= 8'h10 ;
			data[84649] <= 8'h10 ;
			data[84650] <= 8'h10 ;
			data[84651] <= 8'h10 ;
			data[84652] <= 8'h10 ;
			data[84653] <= 8'h10 ;
			data[84654] <= 8'h10 ;
			data[84655] <= 8'h10 ;
			data[84656] <= 8'h10 ;
			data[84657] <= 8'h10 ;
			data[84658] <= 8'h10 ;
			data[84659] <= 8'h10 ;
			data[84660] <= 8'h10 ;
			data[84661] <= 8'h10 ;
			data[84662] <= 8'h10 ;
			data[84663] <= 8'h10 ;
			data[84664] <= 8'h10 ;
			data[84665] <= 8'h10 ;
			data[84666] <= 8'h10 ;
			data[84667] <= 8'h10 ;
			data[84668] <= 8'h10 ;
			data[84669] <= 8'h10 ;
			data[84670] <= 8'h10 ;
			data[84671] <= 8'h10 ;
			data[84672] <= 8'h10 ;
			data[84673] <= 8'h10 ;
			data[84674] <= 8'h10 ;
			data[84675] <= 8'h10 ;
			data[84676] <= 8'h10 ;
			data[84677] <= 8'h10 ;
			data[84678] <= 8'h10 ;
			data[84679] <= 8'h10 ;
			data[84680] <= 8'h10 ;
			data[84681] <= 8'h10 ;
			data[84682] <= 8'h10 ;
			data[84683] <= 8'h10 ;
			data[84684] <= 8'h10 ;
			data[84685] <= 8'h10 ;
			data[84686] <= 8'h10 ;
			data[84687] <= 8'h10 ;
			data[84688] <= 8'h10 ;
			data[84689] <= 8'h10 ;
			data[84690] <= 8'h10 ;
			data[84691] <= 8'h10 ;
			data[84692] <= 8'h10 ;
			data[84693] <= 8'h10 ;
			data[84694] <= 8'h10 ;
			data[84695] <= 8'h10 ;
			data[84696] <= 8'h10 ;
			data[84697] <= 8'h10 ;
			data[84698] <= 8'h10 ;
			data[84699] <= 8'h10 ;
			data[84700] <= 8'h10 ;
			data[84701] <= 8'h10 ;
			data[84702] <= 8'h10 ;
			data[84703] <= 8'h10 ;
			data[84704] <= 8'h10 ;
			data[84705] <= 8'h10 ;
			data[84706] <= 8'h10 ;
			data[84707] <= 8'h10 ;
			data[84708] <= 8'h10 ;
			data[84709] <= 8'h10 ;
			data[84710] <= 8'h10 ;
			data[84711] <= 8'h10 ;
			data[84712] <= 8'h10 ;
			data[84713] <= 8'h10 ;
			data[84714] <= 8'h10 ;
			data[84715] <= 8'h10 ;
			data[84716] <= 8'h10 ;
			data[84717] <= 8'h10 ;
			data[84718] <= 8'h10 ;
			data[84719] <= 8'h10 ;
			data[84720] <= 8'h10 ;
			data[84721] <= 8'h10 ;
			data[84722] <= 8'h10 ;
			data[84723] <= 8'h10 ;
			data[84724] <= 8'h10 ;
			data[84725] <= 8'h10 ;
			data[84726] <= 8'h10 ;
			data[84727] <= 8'h10 ;
			data[84728] <= 8'h10 ;
			data[84729] <= 8'h10 ;
			data[84730] <= 8'h10 ;
			data[84731] <= 8'h10 ;
			data[84732] <= 8'h10 ;
			data[84733] <= 8'h10 ;
			data[84734] <= 8'h10 ;
			data[84735] <= 8'h10 ;
			data[84736] <= 8'h10 ;
			data[84737] <= 8'h10 ;
			data[84738] <= 8'h10 ;
			data[84739] <= 8'h10 ;
			data[84740] <= 8'h10 ;
			data[84741] <= 8'h10 ;
			data[84742] <= 8'h10 ;
			data[84743] <= 8'h10 ;
			data[84744] <= 8'h10 ;
			data[84745] <= 8'h10 ;
			data[84746] <= 8'h10 ;
			data[84747] <= 8'h10 ;
			data[84748] <= 8'h10 ;
			data[84749] <= 8'h10 ;
			data[84750] <= 8'h10 ;
			data[84751] <= 8'h10 ;
			data[84752] <= 8'h10 ;
			data[84753] <= 8'h10 ;
			data[84754] <= 8'h10 ;
			data[84755] <= 8'h10 ;
			data[84756] <= 8'h10 ;
			data[84757] <= 8'h10 ;
			data[84758] <= 8'h10 ;
			data[84759] <= 8'h10 ;
			data[84760] <= 8'h10 ;
			data[84761] <= 8'h10 ;
			data[84762] <= 8'h10 ;
			data[84763] <= 8'h10 ;
			data[84764] <= 8'h10 ;
			data[84765] <= 8'h10 ;
			data[84766] <= 8'h10 ;
			data[84767] <= 8'h10 ;
			data[84768] <= 8'h10 ;
			data[84769] <= 8'h10 ;
			data[84770] <= 8'h10 ;
			data[84771] <= 8'h10 ;
			data[84772] <= 8'h10 ;
			data[84773] <= 8'h10 ;
			data[84774] <= 8'h10 ;
			data[84775] <= 8'h10 ;
			data[84776] <= 8'h10 ;
			data[84777] <= 8'h10 ;
			data[84778] <= 8'h10 ;
			data[84779] <= 8'h10 ;
			data[84780] <= 8'h10 ;
			data[84781] <= 8'h10 ;
			data[84782] <= 8'h10 ;
			data[84783] <= 8'h10 ;
			data[84784] <= 8'h10 ;
			data[84785] <= 8'h10 ;
			data[84786] <= 8'h10 ;
			data[84787] <= 8'h10 ;
			data[84788] <= 8'h10 ;
			data[84789] <= 8'h10 ;
			data[84790] <= 8'h10 ;
			data[84791] <= 8'h10 ;
			data[84792] <= 8'h10 ;
			data[84793] <= 8'h10 ;
			data[84794] <= 8'h10 ;
			data[84795] <= 8'h10 ;
			data[84796] <= 8'h10 ;
			data[84797] <= 8'h10 ;
			data[84798] <= 8'h10 ;
			data[84799] <= 8'h10 ;
			data[84800] <= 8'h10 ;
			data[84801] <= 8'h10 ;
			data[84802] <= 8'h10 ;
			data[84803] <= 8'h10 ;
			data[84804] <= 8'h10 ;
			data[84805] <= 8'h10 ;
			data[84806] <= 8'h10 ;
			data[84807] <= 8'h10 ;
			data[84808] <= 8'h10 ;
			data[84809] <= 8'h10 ;
			data[84810] <= 8'h10 ;
			data[84811] <= 8'h10 ;
			data[84812] <= 8'h10 ;
			data[84813] <= 8'h10 ;
			data[84814] <= 8'h10 ;
			data[84815] <= 8'h10 ;
			data[84816] <= 8'h10 ;
			data[84817] <= 8'h10 ;
			data[84818] <= 8'h10 ;
			data[84819] <= 8'h10 ;
			data[84820] <= 8'h10 ;
			data[84821] <= 8'h10 ;
			data[84822] <= 8'h10 ;
			data[84823] <= 8'h10 ;
			data[84824] <= 8'h10 ;
			data[84825] <= 8'h10 ;
			data[84826] <= 8'h10 ;
			data[84827] <= 8'h10 ;
			data[84828] <= 8'h10 ;
			data[84829] <= 8'h10 ;
			data[84830] <= 8'h10 ;
			data[84831] <= 8'h10 ;
			data[84832] <= 8'h10 ;
			data[84833] <= 8'h10 ;
			data[84834] <= 8'h10 ;
			data[84835] <= 8'h10 ;
			data[84836] <= 8'h10 ;
			data[84837] <= 8'h10 ;
			data[84838] <= 8'h10 ;
			data[84839] <= 8'h10 ;
			data[84840] <= 8'h10 ;
			data[84841] <= 8'h10 ;
			data[84842] <= 8'h10 ;
			data[84843] <= 8'h10 ;
			data[84844] <= 8'h10 ;
			data[84845] <= 8'h10 ;
			data[84846] <= 8'h10 ;
			data[84847] <= 8'h10 ;
			data[84848] <= 8'h10 ;
			data[84849] <= 8'h10 ;
			data[84850] <= 8'h10 ;
			data[84851] <= 8'h10 ;
			data[84852] <= 8'h10 ;
			data[84853] <= 8'h10 ;
			data[84854] <= 8'h10 ;
			data[84855] <= 8'h10 ;
			data[84856] <= 8'h10 ;
			data[84857] <= 8'h10 ;
			data[84858] <= 8'h10 ;
			data[84859] <= 8'h10 ;
			data[84860] <= 8'h10 ;
			data[84861] <= 8'h10 ;
			data[84862] <= 8'h10 ;
			data[84863] <= 8'h10 ;
			data[84864] <= 8'h10 ;
			data[84865] <= 8'h10 ;
			data[84866] <= 8'h10 ;
			data[84867] <= 8'h10 ;
			data[84868] <= 8'h10 ;
			data[84869] <= 8'h10 ;
			data[84870] <= 8'h10 ;
			data[84871] <= 8'h10 ;
			data[84872] <= 8'h10 ;
			data[84873] <= 8'h10 ;
			data[84874] <= 8'h10 ;
			data[84875] <= 8'h10 ;
			data[84876] <= 8'h10 ;
			data[84877] <= 8'h10 ;
			data[84878] <= 8'h10 ;
			data[84879] <= 8'h10 ;
			data[84880] <= 8'h10 ;
			data[84881] <= 8'h10 ;
			data[84882] <= 8'h10 ;
			data[84883] <= 8'h10 ;
			data[84884] <= 8'h10 ;
			data[84885] <= 8'h10 ;
			data[84886] <= 8'h10 ;
			data[84887] <= 8'h10 ;
			data[84888] <= 8'h10 ;
			data[84889] <= 8'h10 ;
			data[84890] <= 8'h10 ;
			data[84891] <= 8'h10 ;
			data[84892] <= 8'h10 ;
			data[84893] <= 8'h10 ;
			data[84894] <= 8'h10 ;
			data[84895] <= 8'h10 ;
			data[84896] <= 8'h10 ;
			data[84897] <= 8'h10 ;
			data[84898] <= 8'h10 ;
			data[84899] <= 8'h10 ;
			data[84900] <= 8'h10 ;
			data[84901] <= 8'h10 ;
			data[84902] <= 8'h10 ;
			data[84903] <= 8'h10 ;
			data[84904] <= 8'h10 ;
			data[84905] <= 8'h10 ;
			data[84906] <= 8'h10 ;
			data[84907] <= 8'h10 ;
			data[84908] <= 8'h10 ;
			data[84909] <= 8'h10 ;
			data[84910] <= 8'h10 ;
			data[84911] <= 8'h10 ;
			data[84912] <= 8'h10 ;
			data[84913] <= 8'h10 ;
			data[84914] <= 8'h10 ;
			data[84915] <= 8'h10 ;
			data[84916] <= 8'h10 ;
			data[84917] <= 8'h10 ;
			data[84918] <= 8'h10 ;
			data[84919] <= 8'h10 ;
			data[84920] <= 8'h10 ;
			data[84921] <= 8'h10 ;
			data[84922] <= 8'h10 ;
			data[84923] <= 8'h10 ;
			data[84924] <= 8'h10 ;
			data[84925] <= 8'h10 ;
			data[84926] <= 8'h10 ;
			data[84927] <= 8'h10 ;
			data[84928] <= 8'h10 ;
			data[84929] <= 8'h10 ;
			data[84930] <= 8'h10 ;
			data[84931] <= 8'h10 ;
			data[84932] <= 8'h10 ;
			data[84933] <= 8'h10 ;
			data[84934] <= 8'h10 ;
			data[84935] <= 8'h10 ;
			data[84936] <= 8'h10 ;
			data[84937] <= 8'h10 ;
			data[84938] <= 8'h10 ;
			data[84939] <= 8'h10 ;
			data[84940] <= 8'h10 ;
			data[84941] <= 8'h10 ;
			data[84942] <= 8'h10 ;
			data[84943] <= 8'h10 ;
			data[84944] <= 8'h10 ;
			data[84945] <= 8'h10 ;
			data[84946] <= 8'h10 ;
			data[84947] <= 8'h10 ;
			data[84948] <= 8'h10 ;
			data[84949] <= 8'h10 ;
			data[84950] <= 8'h10 ;
			data[84951] <= 8'h10 ;
			data[84952] <= 8'h10 ;
			data[84953] <= 8'h10 ;
			data[84954] <= 8'h10 ;
			data[84955] <= 8'h10 ;
			data[84956] <= 8'h10 ;
			data[84957] <= 8'h10 ;
			data[84958] <= 8'h10 ;
			data[84959] <= 8'h10 ;
			data[84960] <= 8'h10 ;
			data[84961] <= 8'h10 ;
			data[84962] <= 8'h10 ;
			data[84963] <= 8'h10 ;
			data[84964] <= 8'h10 ;
			data[84965] <= 8'h10 ;
			data[84966] <= 8'h10 ;
			data[84967] <= 8'h10 ;
			data[84968] <= 8'h10 ;
			data[84969] <= 8'h10 ;
			data[84970] <= 8'h10 ;
			data[84971] <= 8'h10 ;
			data[84972] <= 8'h10 ;
			data[84973] <= 8'h10 ;
			data[84974] <= 8'h10 ;
			data[84975] <= 8'h10 ;
			data[84976] <= 8'h10 ;
			data[84977] <= 8'h10 ;
			data[84978] <= 8'h10 ;
			data[84979] <= 8'h10 ;
			data[84980] <= 8'h10 ;
			data[84981] <= 8'h10 ;
			data[84982] <= 8'h10 ;
			data[84983] <= 8'h10 ;
			data[84984] <= 8'h10 ;
			data[84985] <= 8'h10 ;
			data[84986] <= 8'h10 ;
			data[84987] <= 8'h10 ;
			data[84988] <= 8'h10 ;
			data[84989] <= 8'h10 ;
			data[84990] <= 8'h10 ;
			data[84991] <= 8'h10 ;
			data[84992] <= 8'h10 ;
			data[84993] <= 8'h10 ;
			data[84994] <= 8'h10 ;
			data[84995] <= 8'h10 ;
			data[84996] <= 8'h10 ;
			data[84997] <= 8'h10 ;
			data[84998] <= 8'h10 ;
			data[84999] <= 8'h10 ;
			data[85000] <= 8'h10 ;
			data[85001] <= 8'h10 ;
			data[85002] <= 8'h10 ;
			data[85003] <= 8'h10 ;
			data[85004] <= 8'h10 ;
			data[85005] <= 8'h10 ;
			data[85006] <= 8'h10 ;
			data[85007] <= 8'h10 ;
			data[85008] <= 8'h10 ;
			data[85009] <= 8'h10 ;
			data[85010] <= 8'h10 ;
			data[85011] <= 8'h10 ;
			data[85012] <= 8'h10 ;
			data[85013] <= 8'h10 ;
			data[85014] <= 8'h10 ;
			data[85015] <= 8'h10 ;
			data[85016] <= 8'h10 ;
			data[85017] <= 8'h10 ;
			data[85018] <= 8'h10 ;
			data[85019] <= 8'h10 ;
			data[85020] <= 8'h10 ;
			data[85021] <= 8'h10 ;
			data[85022] <= 8'h10 ;
			data[85023] <= 8'h10 ;
			data[85024] <= 8'h10 ;
			data[85025] <= 8'h10 ;
			data[85026] <= 8'h10 ;
			data[85027] <= 8'h10 ;
			data[85028] <= 8'h10 ;
			data[85029] <= 8'h10 ;
			data[85030] <= 8'h10 ;
			data[85031] <= 8'h10 ;
			data[85032] <= 8'h10 ;
			data[85033] <= 8'h10 ;
			data[85034] <= 8'h10 ;
			data[85035] <= 8'h10 ;
			data[85036] <= 8'h10 ;
			data[85037] <= 8'h10 ;
			data[85038] <= 8'h10 ;
			data[85039] <= 8'h10 ;
			data[85040] <= 8'h10 ;
			data[85041] <= 8'h10 ;
			data[85042] <= 8'h10 ;
			data[85043] <= 8'h10 ;
			data[85044] <= 8'h10 ;
			data[85045] <= 8'h10 ;
			data[85046] <= 8'h10 ;
			data[85047] <= 8'h10 ;
			data[85048] <= 8'h10 ;
			data[85049] <= 8'h10 ;
			data[85050] <= 8'h10 ;
			data[85051] <= 8'h10 ;
			data[85052] <= 8'h10 ;
			data[85053] <= 8'h10 ;
			data[85054] <= 8'h10 ;
			data[85055] <= 8'h10 ;
			data[85056] <= 8'h10 ;
			data[85057] <= 8'h10 ;
			data[85058] <= 8'h10 ;
			data[85059] <= 8'h10 ;
			data[85060] <= 8'h10 ;
			data[85061] <= 8'h10 ;
			data[85062] <= 8'h10 ;
			data[85063] <= 8'h10 ;
			data[85064] <= 8'h10 ;
			data[85065] <= 8'h10 ;
			data[85066] <= 8'h10 ;
			data[85067] <= 8'h10 ;
			data[85068] <= 8'h10 ;
			data[85069] <= 8'h10 ;
			data[85070] <= 8'h10 ;
			data[85071] <= 8'h10 ;
			data[85072] <= 8'h10 ;
			data[85073] <= 8'h10 ;
			data[85074] <= 8'h10 ;
			data[85075] <= 8'h10 ;
			data[85076] <= 8'h10 ;
			data[85077] <= 8'h10 ;
			data[85078] <= 8'h10 ;
			data[85079] <= 8'h10 ;
			data[85080] <= 8'h10 ;
			data[85081] <= 8'h10 ;
			data[85082] <= 8'h10 ;
			data[85083] <= 8'h10 ;
			data[85084] <= 8'h10 ;
			data[85085] <= 8'h10 ;
			data[85086] <= 8'h10 ;
			data[85087] <= 8'h10 ;
			data[85088] <= 8'h10 ;
			data[85089] <= 8'h10 ;
			data[85090] <= 8'h10 ;
			data[85091] <= 8'h10 ;
			data[85092] <= 8'h10 ;
			data[85093] <= 8'h10 ;
			data[85094] <= 8'h10 ;
			data[85095] <= 8'h10 ;
			data[85096] <= 8'h10 ;
			data[85097] <= 8'h10 ;
			data[85098] <= 8'h10 ;
			data[85099] <= 8'h10 ;
			data[85100] <= 8'h10 ;
			data[85101] <= 8'h10 ;
			data[85102] <= 8'h10 ;
			data[85103] <= 8'h10 ;
			data[85104] <= 8'h10 ;
			data[85105] <= 8'h10 ;
			data[85106] <= 8'h10 ;
			data[85107] <= 8'h10 ;
			data[85108] <= 8'h10 ;
			data[85109] <= 8'h10 ;
			data[85110] <= 8'h10 ;
			data[85111] <= 8'h10 ;
			data[85112] <= 8'h10 ;
			data[85113] <= 8'h10 ;
			data[85114] <= 8'h10 ;
			data[85115] <= 8'h10 ;
			data[85116] <= 8'h10 ;
			data[85117] <= 8'h10 ;
			data[85118] <= 8'h10 ;
			data[85119] <= 8'h10 ;
			data[85120] <= 8'h10 ;
			data[85121] <= 8'h10 ;
			data[85122] <= 8'h10 ;
			data[85123] <= 8'h10 ;
			data[85124] <= 8'h10 ;
			data[85125] <= 8'h10 ;
			data[85126] <= 8'h10 ;
			data[85127] <= 8'h10 ;
			data[85128] <= 8'h10 ;
			data[85129] <= 8'h10 ;
			data[85130] <= 8'h10 ;
			data[85131] <= 8'h10 ;
			data[85132] <= 8'h10 ;
			data[85133] <= 8'h10 ;
			data[85134] <= 8'h10 ;
			data[85135] <= 8'h10 ;
			data[85136] <= 8'h10 ;
			data[85137] <= 8'h10 ;
			data[85138] <= 8'h10 ;
			data[85139] <= 8'h10 ;
			data[85140] <= 8'h10 ;
			data[85141] <= 8'h10 ;
			data[85142] <= 8'h10 ;
			data[85143] <= 8'h10 ;
			data[85144] <= 8'h10 ;
			data[85145] <= 8'h10 ;
			data[85146] <= 8'h10 ;
			data[85147] <= 8'h10 ;
			data[85148] <= 8'h10 ;
			data[85149] <= 8'h10 ;
			data[85150] <= 8'h10 ;
			data[85151] <= 8'h10 ;
			data[85152] <= 8'h10 ;
			data[85153] <= 8'h10 ;
			data[85154] <= 8'h10 ;
			data[85155] <= 8'h10 ;
			data[85156] <= 8'h10 ;
			data[85157] <= 8'h10 ;
			data[85158] <= 8'h10 ;
			data[85159] <= 8'h10 ;
			data[85160] <= 8'h10 ;
			data[85161] <= 8'h10 ;
			data[85162] <= 8'h10 ;
			data[85163] <= 8'h10 ;
			data[85164] <= 8'h10 ;
			data[85165] <= 8'h10 ;
			data[85166] <= 8'h10 ;
			data[85167] <= 8'h10 ;
			data[85168] <= 8'h10 ;
			data[85169] <= 8'h10 ;
			data[85170] <= 8'h10 ;
			data[85171] <= 8'h10 ;
			data[85172] <= 8'h10 ;
			data[85173] <= 8'h10 ;
			data[85174] <= 8'h10 ;
			data[85175] <= 8'h10 ;
			data[85176] <= 8'h10 ;
			data[85177] <= 8'h10 ;
			data[85178] <= 8'h10 ;
			data[85179] <= 8'h10 ;
			data[85180] <= 8'h10 ;
			data[85181] <= 8'h10 ;
			data[85182] <= 8'h10 ;
			data[85183] <= 8'h10 ;
			data[85184] <= 8'h10 ;
			data[85185] <= 8'h10 ;
			data[85186] <= 8'h10 ;
			data[85187] <= 8'h10 ;
			data[85188] <= 8'h10 ;
			data[85189] <= 8'h10 ;
			data[85190] <= 8'h10 ;
			data[85191] <= 8'h10 ;
			data[85192] <= 8'h10 ;
			data[85193] <= 8'h10 ;
			data[85194] <= 8'h10 ;
			data[85195] <= 8'h10 ;
			data[85196] <= 8'h10 ;
			data[85197] <= 8'h10 ;
			data[85198] <= 8'h10 ;
			data[85199] <= 8'h10 ;
			data[85200] <= 8'h10 ;
			data[85201] <= 8'h10 ;
			data[85202] <= 8'h10 ;
			data[85203] <= 8'h10 ;
			data[85204] <= 8'h10 ;
			data[85205] <= 8'h10 ;
			data[85206] <= 8'h10 ;
			data[85207] <= 8'h10 ;
			data[85208] <= 8'h10 ;
			data[85209] <= 8'h10 ;
			data[85210] <= 8'h10 ;
			data[85211] <= 8'h10 ;
			data[85212] <= 8'h10 ;
			data[85213] <= 8'h10 ;
			data[85214] <= 8'h10 ;
			data[85215] <= 8'h10 ;
			data[85216] <= 8'h10 ;
			data[85217] <= 8'h10 ;
			data[85218] <= 8'h10 ;
			data[85219] <= 8'h10 ;
			data[85220] <= 8'h10 ;
			data[85221] <= 8'h10 ;
			data[85222] <= 8'h10 ;
			data[85223] <= 8'h10 ;
			data[85224] <= 8'h10 ;
			data[85225] <= 8'h10 ;
			data[85226] <= 8'h10 ;
			data[85227] <= 8'h10 ;
			data[85228] <= 8'h10 ;
			data[85229] <= 8'h10 ;
			data[85230] <= 8'h10 ;
			data[85231] <= 8'h10 ;
			data[85232] <= 8'h10 ;
			data[85233] <= 8'h10 ;
			data[85234] <= 8'h10 ;
			data[85235] <= 8'h10 ;
			data[85236] <= 8'h10 ;
			data[85237] <= 8'h10 ;
			data[85238] <= 8'h10 ;
			data[85239] <= 8'h10 ;
			data[85240] <= 8'h10 ;
			data[85241] <= 8'h10 ;
			data[85242] <= 8'h10 ;
			data[85243] <= 8'h10 ;
			data[85244] <= 8'h10 ;
			data[85245] <= 8'h10 ;
			data[85246] <= 8'h10 ;
			data[85247] <= 8'h10 ;
			data[85248] <= 8'h10 ;
			data[85249] <= 8'h10 ;
			data[85250] <= 8'h10 ;
			data[85251] <= 8'h10 ;
			data[85252] <= 8'h10 ;
			data[85253] <= 8'h10 ;
			data[85254] <= 8'h10 ;
			data[85255] <= 8'h10 ;
			data[85256] <= 8'h10 ;
			data[85257] <= 8'h10 ;
			data[85258] <= 8'h10 ;
			data[85259] <= 8'h10 ;
			data[85260] <= 8'h10 ;
			data[85261] <= 8'h10 ;
			data[85262] <= 8'h10 ;
			data[85263] <= 8'h10 ;
			data[85264] <= 8'h10 ;
			data[85265] <= 8'h10 ;
			data[85266] <= 8'h10 ;
			data[85267] <= 8'h10 ;
			data[85268] <= 8'h10 ;
			data[85269] <= 8'h10 ;
			data[85270] <= 8'h10 ;
			data[85271] <= 8'h10 ;
			data[85272] <= 8'h10 ;
			data[85273] <= 8'h10 ;
			data[85274] <= 8'h10 ;
			data[85275] <= 8'h10 ;
			data[85276] <= 8'h10 ;
			data[85277] <= 8'h10 ;
			data[85278] <= 8'h10 ;
			data[85279] <= 8'h10 ;
			data[85280] <= 8'h10 ;
			data[85281] <= 8'h10 ;
			data[85282] <= 8'h10 ;
			data[85283] <= 8'h10 ;
			data[85284] <= 8'h10 ;
			data[85285] <= 8'h10 ;
			data[85286] <= 8'h10 ;
			data[85287] <= 8'h10 ;
			data[85288] <= 8'h10 ;
			data[85289] <= 8'h10 ;
			data[85290] <= 8'h10 ;
			data[85291] <= 8'h10 ;
			data[85292] <= 8'h10 ;
			data[85293] <= 8'h10 ;
			data[85294] <= 8'h10 ;
			data[85295] <= 8'h10 ;
			data[85296] <= 8'h10 ;
			data[85297] <= 8'h10 ;
			data[85298] <= 8'h10 ;
			data[85299] <= 8'h10 ;
			data[85300] <= 8'h10 ;
			data[85301] <= 8'h10 ;
			data[85302] <= 8'h10 ;
			data[85303] <= 8'h10 ;
			data[85304] <= 8'h10 ;
			data[85305] <= 8'h10 ;
			data[85306] <= 8'h10 ;
			data[85307] <= 8'h10 ;
			data[85308] <= 8'h10 ;
			data[85309] <= 8'h10 ;
			data[85310] <= 8'h10 ;
			data[85311] <= 8'h10 ;
			data[85312] <= 8'h10 ;
			data[85313] <= 8'h10 ;
			data[85314] <= 8'h10 ;
			data[85315] <= 8'h10 ;
			data[85316] <= 8'h10 ;
			data[85317] <= 8'h10 ;
			data[85318] <= 8'h10 ;
			data[85319] <= 8'h10 ;
			data[85320] <= 8'h10 ;
			data[85321] <= 8'h10 ;
			data[85322] <= 8'h10 ;
			data[85323] <= 8'h10 ;
			data[85324] <= 8'h10 ;
			data[85325] <= 8'h10 ;
			data[85326] <= 8'h10 ;
			data[85327] <= 8'h10 ;
			data[85328] <= 8'h10 ;
			data[85329] <= 8'h10 ;
			data[85330] <= 8'h10 ;
			data[85331] <= 8'h10 ;
			data[85332] <= 8'h10 ;
			data[85333] <= 8'h10 ;
			data[85334] <= 8'h10 ;
			data[85335] <= 8'h10 ;
			data[85336] <= 8'h10 ;
			data[85337] <= 8'h10 ;
			data[85338] <= 8'h10 ;
			data[85339] <= 8'h10 ;
			data[85340] <= 8'h10 ;
			data[85341] <= 8'h10 ;
			data[85342] <= 8'h10 ;
			data[85343] <= 8'h10 ;
			data[85344] <= 8'h10 ;
			data[85345] <= 8'h10 ;
			data[85346] <= 8'h10 ;
			data[85347] <= 8'h10 ;
			data[85348] <= 8'h10 ;
			data[85349] <= 8'h10 ;
			data[85350] <= 8'h10 ;
			data[85351] <= 8'h10 ;
			data[85352] <= 8'h10 ;
			data[85353] <= 8'h10 ;
			data[85354] <= 8'h10 ;
			data[85355] <= 8'h10 ;
			data[85356] <= 8'h10 ;
			data[85357] <= 8'h10 ;
			data[85358] <= 8'h10 ;
			data[85359] <= 8'h10 ;
			data[85360] <= 8'h10 ;
			data[85361] <= 8'h10 ;
			data[85362] <= 8'h10 ;
			data[85363] <= 8'h10 ;
			data[85364] <= 8'h10 ;
			data[85365] <= 8'h10 ;
			data[85366] <= 8'h10 ;
			data[85367] <= 8'h10 ;
			data[85368] <= 8'h10 ;
			data[85369] <= 8'h10 ;
			data[85370] <= 8'h10 ;
			data[85371] <= 8'h10 ;
			data[85372] <= 8'h10 ;
			data[85373] <= 8'h10 ;
			data[85374] <= 8'h10 ;
			data[85375] <= 8'h10 ;
			data[85376] <= 8'h10 ;
			data[85377] <= 8'h10 ;
			data[85378] <= 8'h10 ;
			data[85379] <= 8'h10 ;
			data[85380] <= 8'h10 ;
			data[85381] <= 8'h10 ;
			data[85382] <= 8'h10 ;
			data[85383] <= 8'h10 ;
			data[85384] <= 8'h10 ;
			data[85385] <= 8'h10 ;
			data[85386] <= 8'h10 ;
			data[85387] <= 8'h10 ;
			data[85388] <= 8'h10 ;
			data[85389] <= 8'h10 ;
			data[85390] <= 8'h10 ;
			data[85391] <= 8'h10 ;
			data[85392] <= 8'h10 ;
			data[85393] <= 8'h10 ;
			data[85394] <= 8'h10 ;
			data[85395] <= 8'h10 ;
			data[85396] <= 8'h10 ;
			data[85397] <= 8'h10 ;
			data[85398] <= 8'h10 ;
			data[85399] <= 8'h10 ;
			data[85400] <= 8'h10 ;
			data[85401] <= 8'h10 ;
			data[85402] <= 8'h10 ;
			data[85403] <= 8'h10 ;
			data[85404] <= 8'h10 ;
			data[85405] <= 8'h10 ;
			data[85406] <= 8'h10 ;
			data[85407] <= 8'h10 ;
			data[85408] <= 8'h10 ;
			data[85409] <= 8'h10 ;
			data[85410] <= 8'h10 ;
			data[85411] <= 8'h10 ;
			data[85412] <= 8'h10 ;
			data[85413] <= 8'h10 ;
			data[85414] <= 8'h10 ;
			data[85415] <= 8'h10 ;
			data[85416] <= 8'h10 ;
			data[85417] <= 8'h10 ;
			data[85418] <= 8'h10 ;
			data[85419] <= 8'h10 ;
			data[85420] <= 8'h10 ;
			data[85421] <= 8'h10 ;
			data[85422] <= 8'h10 ;
			data[85423] <= 8'h10 ;
			data[85424] <= 8'h10 ;
			data[85425] <= 8'h10 ;
			data[85426] <= 8'h10 ;
			data[85427] <= 8'h10 ;
			data[85428] <= 8'h10 ;
			data[85429] <= 8'h10 ;
			data[85430] <= 8'h10 ;
			data[85431] <= 8'h10 ;
			data[85432] <= 8'h10 ;
			data[85433] <= 8'h10 ;
			data[85434] <= 8'h10 ;
			data[85435] <= 8'h10 ;
			data[85436] <= 8'h10 ;
			data[85437] <= 8'h10 ;
			data[85438] <= 8'h10 ;
			data[85439] <= 8'h10 ;
			data[85440] <= 8'h10 ;
			data[85441] <= 8'h10 ;
			data[85442] <= 8'h10 ;
			data[85443] <= 8'h10 ;
			data[85444] <= 8'h10 ;
			data[85445] <= 8'h10 ;
			data[85446] <= 8'h10 ;
			data[85447] <= 8'h10 ;
			data[85448] <= 8'h10 ;
			data[85449] <= 8'h10 ;
			data[85450] <= 8'h10 ;
			data[85451] <= 8'h10 ;
			data[85452] <= 8'h10 ;
			data[85453] <= 8'h10 ;
			data[85454] <= 8'h10 ;
			data[85455] <= 8'h10 ;
			data[85456] <= 8'h10 ;
			data[85457] <= 8'h10 ;
			data[85458] <= 8'h10 ;
			data[85459] <= 8'h10 ;
			data[85460] <= 8'h10 ;
			data[85461] <= 8'h10 ;
			data[85462] <= 8'h10 ;
			data[85463] <= 8'h10 ;
			data[85464] <= 8'h10 ;
			data[85465] <= 8'h10 ;
			data[85466] <= 8'h10 ;
			data[85467] <= 8'h10 ;
			data[85468] <= 8'h10 ;
			data[85469] <= 8'h10 ;
			data[85470] <= 8'h10 ;
			data[85471] <= 8'h10 ;
			data[85472] <= 8'h10 ;
			data[85473] <= 8'h10 ;
			data[85474] <= 8'h10 ;
			data[85475] <= 8'h10 ;
			data[85476] <= 8'h10 ;
			data[85477] <= 8'h10 ;
			data[85478] <= 8'h10 ;
			data[85479] <= 8'h10 ;
			data[85480] <= 8'h10 ;
			data[85481] <= 8'h10 ;
			data[85482] <= 8'h10 ;
			data[85483] <= 8'h10 ;
			data[85484] <= 8'h10 ;
			data[85485] <= 8'h10 ;
			data[85486] <= 8'h10 ;
			data[85487] <= 8'h10 ;
			data[85488] <= 8'h10 ;
			data[85489] <= 8'h10 ;
			data[85490] <= 8'h10 ;
			data[85491] <= 8'h10 ;
			data[85492] <= 8'h10 ;
			data[85493] <= 8'h10 ;
			data[85494] <= 8'h10 ;
			data[85495] <= 8'h10 ;
			data[85496] <= 8'h10 ;
			data[85497] <= 8'h10 ;
			data[85498] <= 8'h10 ;
			data[85499] <= 8'h10 ;
			data[85500] <= 8'h10 ;
			data[85501] <= 8'h10 ;
			data[85502] <= 8'h10 ;
			data[85503] <= 8'h10 ;
			data[85504] <= 8'h10 ;
			data[85505] <= 8'h10 ;
			data[85506] <= 8'h10 ;
			data[85507] <= 8'h10 ;
			data[85508] <= 8'h10 ;
			data[85509] <= 8'h10 ;
			data[85510] <= 8'h10 ;
			data[85511] <= 8'h10 ;
			data[85512] <= 8'h10 ;
			data[85513] <= 8'h10 ;
			data[85514] <= 8'h10 ;
			data[85515] <= 8'h10 ;
			data[85516] <= 8'h10 ;
			data[85517] <= 8'h10 ;
			data[85518] <= 8'h10 ;
			data[85519] <= 8'h10 ;
			data[85520] <= 8'h10 ;
			data[85521] <= 8'h10 ;
			data[85522] <= 8'h10 ;
			data[85523] <= 8'h10 ;
			data[85524] <= 8'h10 ;
			data[85525] <= 8'h10 ;
			data[85526] <= 8'h10 ;
			data[85527] <= 8'h10 ;
			data[85528] <= 8'h10 ;
			data[85529] <= 8'h10 ;
			data[85530] <= 8'h10 ;
			data[85531] <= 8'h10 ;
			data[85532] <= 8'h10 ;
			data[85533] <= 8'h10 ;
			data[85534] <= 8'h10 ;
			data[85535] <= 8'h10 ;
			data[85536] <= 8'h10 ;
			data[85537] <= 8'h10 ;
			data[85538] <= 8'h10 ;
			data[85539] <= 8'h10 ;
			data[85540] <= 8'h10 ;
			data[85541] <= 8'h10 ;
			data[85542] <= 8'h10 ;
			data[85543] <= 8'h10 ;
			data[85544] <= 8'h10 ;
			data[85545] <= 8'h10 ;
			data[85546] <= 8'h10 ;
			data[85547] <= 8'h10 ;
			data[85548] <= 8'h10 ;
			data[85549] <= 8'h10 ;
			data[85550] <= 8'h10 ;
			data[85551] <= 8'h10 ;
			data[85552] <= 8'h10 ;
			data[85553] <= 8'h10 ;
			data[85554] <= 8'h10 ;
			data[85555] <= 8'h10 ;
			data[85556] <= 8'h10 ;
			data[85557] <= 8'h10 ;
			data[85558] <= 8'h10 ;
			data[85559] <= 8'h10 ;
			data[85560] <= 8'h10 ;
			data[85561] <= 8'h10 ;
			data[85562] <= 8'h10 ;
			data[85563] <= 8'h10 ;
			data[85564] <= 8'h10 ;
			data[85565] <= 8'h10 ;
			data[85566] <= 8'h10 ;
			data[85567] <= 8'h10 ;
			data[85568] <= 8'h10 ;
			data[85569] <= 8'h10 ;
			data[85570] <= 8'h10 ;
			data[85571] <= 8'h10 ;
			data[85572] <= 8'h10 ;
			data[85573] <= 8'h10 ;
			data[85574] <= 8'h10 ;
			data[85575] <= 8'h10 ;
			data[85576] <= 8'h10 ;
			data[85577] <= 8'h10 ;
			data[85578] <= 8'h10 ;
			data[85579] <= 8'h10 ;
			data[85580] <= 8'h10 ;
			data[85581] <= 8'h10 ;
			data[85582] <= 8'h10 ;
			data[85583] <= 8'h10 ;
			data[85584] <= 8'h10 ;
			data[85585] <= 8'h10 ;
			data[85586] <= 8'h10 ;
			data[85587] <= 8'h10 ;
			data[85588] <= 8'h10 ;
			data[85589] <= 8'h10 ;
			data[85590] <= 8'h10 ;
			data[85591] <= 8'h10 ;
			data[85592] <= 8'h10 ;
			data[85593] <= 8'h10 ;
			data[85594] <= 8'h10 ;
			data[85595] <= 8'h10 ;
			data[85596] <= 8'h10 ;
			data[85597] <= 8'h10 ;
			data[85598] <= 8'h10 ;
			data[85599] <= 8'h10 ;
			data[85600] <= 8'h10 ;
			data[85601] <= 8'h10 ;
			data[85602] <= 8'h10 ;
			data[85603] <= 8'h10 ;
			data[85604] <= 8'h10 ;
			data[85605] <= 8'h10 ;
			data[85606] <= 8'h10 ;
			data[85607] <= 8'h10 ;
			data[85608] <= 8'h10 ;
			data[85609] <= 8'h10 ;
			data[85610] <= 8'h10 ;
			data[85611] <= 8'h10 ;
			data[85612] <= 8'h10 ;
			data[85613] <= 8'h10 ;
			data[85614] <= 8'h10 ;
			data[85615] <= 8'h10 ;
			data[85616] <= 8'h10 ;
			data[85617] <= 8'h10 ;
			data[85618] <= 8'h10 ;
			data[85619] <= 8'h10 ;
			data[85620] <= 8'h10 ;
			data[85621] <= 8'h10 ;
			data[85622] <= 8'h10 ;
			data[85623] <= 8'h10 ;
			data[85624] <= 8'h10 ;
			data[85625] <= 8'h10 ;
			data[85626] <= 8'h10 ;
			data[85627] <= 8'h10 ;
			data[85628] <= 8'h10 ;
			data[85629] <= 8'h10 ;
			data[85630] <= 8'h10 ;
			data[85631] <= 8'h10 ;
			data[85632] <= 8'h10 ;
			data[85633] <= 8'h10 ;
			data[85634] <= 8'h10 ;
			data[85635] <= 8'h10 ;
			data[85636] <= 8'h10 ;
			data[85637] <= 8'h10 ;
			data[85638] <= 8'h10 ;
			data[85639] <= 8'h10 ;
			data[85640] <= 8'h10 ;
			data[85641] <= 8'h10 ;
			data[85642] <= 8'h10 ;
			data[85643] <= 8'h10 ;
			data[85644] <= 8'h10 ;
			data[85645] <= 8'h10 ;
			data[85646] <= 8'h10 ;
			data[85647] <= 8'h10 ;
			data[85648] <= 8'h10 ;
			data[85649] <= 8'h10 ;
			data[85650] <= 8'h10 ;
			data[85651] <= 8'h10 ;
			data[85652] <= 8'h10 ;
			data[85653] <= 8'h10 ;
			data[85654] <= 8'h10 ;
			data[85655] <= 8'h10 ;
			data[85656] <= 8'h10 ;
			data[85657] <= 8'h10 ;
			data[85658] <= 8'h10 ;
			data[85659] <= 8'h10 ;
			data[85660] <= 8'h10 ;
			data[85661] <= 8'h10 ;
			data[85662] <= 8'h10 ;
			data[85663] <= 8'h10 ;
			data[85664] <= 8'h10 ;
			data[85665] <= 8'h10 ;
			data[85666] <= 8'h10 ;
			data[85667] <= 8'h10 ;
			data[85668] <= 8'h10 ;
			data[85669] <= 8'h10 ;
			data[85670] <= 8'h10 ;
			data[85671] <= 8'h10 ;
			data[85672] <= 8'h10 ;
			data[85673] <= 8'h10 ;
			data[85674] <= 8'h10 ;
			data[85675] <= 8'h10 ;
			data[85676] <= 8'h10 ;
			data[85677] <= 8'h10 ;
			data[85678] <= 8'h10 ;
			data[85679] <= 8'h10 ;
			data[85680] <= 8'h10 ;
			data[85681] <= 8'h10 ;
			data[85682] <= 8'h10 ;
			data[85683] <= 8'h10 ;
			data[85684] <= 8'h10 ;
			data[85685] <= 8'h10 ;
			data[85686] <= 8'h10 ;
			data[85687] <= 8'h10 ;
			data[85688] <= 8'h10 ;
			data[85689] <= 8'h10 ;
			data[85690] <= 8'h10 ;
			data[85691] <= 8'h10 ;
			data[85692] <= 8'h10 ;
			data[85693] <= 8'h10 ;
			data[85694] <= 8'h10 ;
			data[85695] <= 8'h10 ;
			data[85696] <= 8'h10 ;
			data[85697] <= 8'h10 ;
			data[85698] <= 8'h10 ;
			data[85699] <= 8'h10 ;
			data[85700] <= 8'h10 ;
			data[85701] <= 8'h10 ;
			data[85702] <= 8'h10 ;
			data[85703] <= 8'h10 ;
			data[85704] <= 8'h10 ;
			data[85705] <= 8'h10 ;
			data[85706] <= 8'h10 ;
			data[85707] <= 8'h10 ;
			data[85708] <= 8'h10 ;
			data[85709] <= 8'h10 ;
			data[85710] <= 8'h10 ;
			data[85711] <= 8'h10 ;
			data[85712] <= 8'h10 ;
			data[85713] <= 8'h10 ;
			data[85714] <= 8'h10 ;
			data[85715] <= 8'h10 ;
			data[85716] <= 8'h10 ;
			data[85717] <= 8'h10 ;
			data[85718] <= 8'h10 ;
			data[85719] <= 8'h10 ;
			data[85720] <= 8'h10 ;
			data[85721] <= 8'h10 ;
			data[85722] <= 8'h10 ;
			data[85723] <= 8'h10 ;
			data[85724] <= 8'h10 ;
			data[85725] <= 8'h10 ;
			data[85726] <= 8'h10 ;
			data[85727] <= 8'h10 ;
			data[85728] <= 8'h10 ;
			data[85729] <= 8'h10 ;
			data[85730] <= 8'h10 ;
			data[85731] <= 8'h10 ;
			data[85732] <= 8'h10 ;
			data[85733] <= 8'h10 ;
			data[85734] <= 8'h10 ;
			data[85735] <= 8'h10 ;
			data[85736] <= 8'h10 ;
			data[85737] <= 8'h10 ;
			data[85738] <= 8'h10 ;
			data[85739] <= 8'h10 ;
			data[85740] <= 8'h10 ;
			data[85741] <= 8'h10 ;
			data[85742] <= 8'h10 ;
			data[85743] <= 8'h10 ;
			data[85744] <= 8'h10 ;
			data[85745] <= 8'h10 ;
			data[85746] <= 8'h10 ;
			data[85747] <= 8'h10 ;
			data[85748] <= 8'h10 ;
			data[85749] <= 8'h10 ;
			data[85750] <= 8'h10 ;
			data[85751] <= 8'h10 ;
			data[85752] <= 8'h10 ;
			data[85753] <= 8'h10 ;
			data[85754] <= 8'h10 ;
			data[85755] <= 8'h10 ;
			data[85756] <= 8'h10 ;
			data[85757] <= 8'h10 ;
			data[85758] <= 8'h10 ;
			data[85759] <= 8'h10 ;
			data[85760] <= 8'h10 ;
			data[85761] <= 8'h10 ;
			data[85762] <= 8'h10 ;
			data[85763] <= 8'h10 ;
			data[85764] <= 8'h10 ;
			data[85765] <= 8'h10 ;
			data[85766] <= 8'h10 ;
			data[85767] <= 8'h10 ;
			data[85768] <= 8'h10 ;
			data[85769] <= 8'h10 ;
			data[85770] <= 8'h10 ;
			data[85771] <= 8'h10 ;
			data[85772] <= 8'h10 ;
			data[85773] <= 8'h10 ;
			data[85774] <= 8'h10 ;
			data[85775] <= 8'h10 ;
			data[85776] <= 8'h10 ;
			data[85777] <= 8'h10 ;
			data[85778] <= 8'h10 ;
			data[85779] <= 8'h10 ;
			data[85780] <= 8'h10 ;
			data[85781] <= 8'h10 ;
			data[85782] <= 8'h10 ;
			data[85783] <= 8'h10 ;
			data[85784] <= 8'h10 ;
			data[85785] <= 8'h10 ;
			data[85786] <= 8'h10 ;
			data[85787] <= 8'h10 ;
			data[85788] <= 8'h10 ;
			data[85789] <= 8'h10 ;
			data[85790] <= 8'h10 ;
			data[85791] <= 8'h10 ;
			data[85792] <= 8'h10 ;
			data[85793] <= 8'h10 ;
			data[85794] <= 8'h10 ;
			data[85795] <= 8'h10 ;
			data[85796] <= 8'h10 ;
			data[85797] <= 8'h10 ;
			data[85798] <= 8'h10 ;
			data[85799] <= 8'h10 ;
			data[85800] <= 8'h10 ;
			data[85801] <= 8'h10 ;
			data[85802] <= 8'h10 ;
			data[85803] <= 8'h10 ;
			data[85804] <= 8'h10 ;
			data[85805] <= 8'h10 ;
			data[85806] <= 8'h10 ;
			data[85807] <= 8'h10 ;
			data[85808] <= 8'h10 ;
			data[85809] <= 8'h10 ;
			data[85810] <= 8'h10 ;
			data[85811] <= 8'h10 ;
			data[85812] <= 8'h10 ;
			data[85813] <= 8'h10 ;
			data[85814] <= 8'h10 ;
			data[85815] <= 8'h10 ;
			data[85816] <= 8'h10 ;
			data[85817] <= 8'h10 ;
			data[85818] <= 8'h10 ;
			data[85819] <= 8'h10 ;
			data[85820] <= 8'h10 ;
			data[85821] <= 8'h10 ;
			data[85822] <= 8'h10 ;
			data[85823] <= 8'h10 ;
			data[85824] <= 8'h10 ;
			data[85825] <= 8'h10 ;
			data[85826] <= 8'h10 ;
			data[85827] <= 8'h10 ;
			data[85828] <= 8'h10 ;
			data[85829] <= 8'h10 ;
			data[85830] <= 8'h10 ;
			data[85831] <= 8'h10 ;
			data[85832] <= 8'h10 ;
			data[85833] <= 8'h10 ;
			data[85834] <= 8'h10 ;
			data[85835] <= 8'h10 ;
			data[85836] <= 8'h10 ;
			data[85837] <= 8'h10 ;
			data[85838] <= 8'h10 ;
			data[85839] <= 8'h10 ;
			data[85840] <= 8'h10 ;
			data[85841] <= 8'h10 ;
			data[85842] <= 8'h10 ;
			data[85843] <= 8'h10 ;
			data[85844] <= 8'h10 ;
			data[85845] <= 8'h10 ;
			data[85846] <= 8'h10 ;
			data[85847] <= 8'h10 ;
			data[85848] <= 8'h10 ;
			data[85849] <= 8'h10 ;
			data[85850] <= 8'h10 ;
			data[85851] <= 8'h10 ;
			data[85852] <= 8'h10 ;
			data[85853] <= 8'h10 ;
			data[85854] <= 8'h10 ;
			data[85855] <= 8'h10 ;
			data[85856] <= 8'h10 ;
			data[85857] <= 8'h10 ;
			data[85858] <= 8'h10 ;
			data[85859] <= 8'h10 ;
			data[85860] <= 8'h10 ;
			data[85861] <= 8'h10 ;
			data[85862] <= 8'h10 ;
			data[85863] <= 8'h10 ;
			data[85864] <= 8'h10 ;
			data[85865] <= 8'h10 ;
			data[85866] <= 8'h10 ;
			data[85867] <= 8'h10 ;
			data[85868] <= 8'h10 ;
			data[85869] <= 8'h10 ;
			data[85870] <= 8'h10 ;
			data[85871] <= 8'h10 ;
			data[85872] <= 8'h10 ;
			data[85873] <= 8'h10 ;
			data[85874] <= 8'h10 ;
			data[85875] <= 8'h10 ;
			data[85876] <= 8'h10 ;
			data[85877] <= 8'h10 ;
			data[85878] <= 8'h10 ;
			data[85879] <= 8'h10 ;
			data[85880] <= 8'h10 ;
			data[85881] <= 8'h10 ;
			data[85882] <= 8'h10 ;
			data[85883] <= 8'h10 ;
			data[85884] <= 8'h10 ;
			data[85885] <= 8'h10 ;
			data[85886] <= 8'h10 ;
			data[85887] <= 8'h10 ;
			data[85888] <= 8'h10 ;
			data[85889] <= 8'h10 ;
			data[85890] <= 8'h10 ;
			data[85891] <= 8'h10 ;
			data[85892] <= 8'h10 ;
			data[85893] <= 8'h10 ;
			data[85894] <= 8'h10 ;
			data[85895] <= 8'h10 ;
			data[85896] <= 8'h10 ;
			data[85897] <= 8'h10 ;
			data[85898] <= 8'h10 ;
			data[85899] <= 8'h10 ;
			data[85900] <= 8'h10 ;
			data[85901] <= 8'h10 ;
			data[85902] <= 8'h10 ;
			data[85903] <= 8'h10 ;
			data[85904] <= 8'h10 ;
			data[85905] <= 8'h10 ;
			data[85906] <= 8'h10 ;
			data[85907] <= 8'h10 ;
			data[85908] <= 8'h10 ;
			data[85909] <= 8'h10 ;
			data[85910] <= 8'h10 ;
			data[85911] <= 8'h10 ;
			data[85912] <= 8'h10 ;
			data[85913] <= 8'h10 ;
			data[85914] <= 8'h10 ;
			data[85915] <= 8'h10 ;
			data[85916] <= 8'h10 ;
			data[85917] <= 8'h10 ;
			data[85918] <= 8'h10 ;
			data[85919] <= 8'h10 ;
			data[85920] <= 8'h10 ;
			data[85921] <= 8'h10 ;
			data[85922] <= 8'h10 ;
			data[85923] <= 8'h10 ;
			data[85924] <= 8'h10 ;
			data[85925] <= 8'h10 ;
			data[85926] <= 8'h10 ;
			data[85927] <= 8'h10 ;
			data[85928] <= 8'h10 ;
			data[85929] <= 8'h10 ;
			data[85930] <= 8'h10 ;
			data[85931] <= 8'h10 ;
			data[85932] <= 8'h10 ;
			data[85933] <= 8'h10 ;
			data[85934] <= 8'h10 ;
			data[85935] <= 8'h10 ;
			data[85936] <= 8'h10 ;
			data[85937] <= 8'h10 ;
			data[85938] <= 8'h10 ;
			data[85939] <= 8'h10 ;
			data[85940] <= 8'h10 ;
			data[85941] <= 8'h10 ;
			data[85942] <= 8'h10 ;
			data[85943] <= 8'h10 ;
			data[85944] <= 8'h10 ;
			data[85945] <= 8'h10 ;
			data[85946] <= 8'h10 ;
			data[85947] <= 8'h10 ;
			data[85948] <= 8'h10 ;
			data[85949] <= 8'h10 ;
			data[85950] <= 8'h10 ;
			data[85951] <= 8'h10 ;
			data[85952] <= 8'h10 ;
			data[85953] <= 8'h10 ;
			data[85954] <= 8'h10 ;
			data[85955] <= 8'h10 ;
			data[85956] <= 8'h10 ;
			data[85957] <= 8'h10 ;
			data[85958] <= 8'h10 ;
			data[85959] <= 8'h10 ;
			data[85960] <= 8'h10 ;
			data[85961] <= 8'h10 ;
			data[85962] <= 8'h10 ;
			data[85963] <= 8'h10 ;
			data[85964] <= 8'h10 ;
			data[85965] <= 8'h10 ;
			data[85966] <= 8'h10 ;
			data[85967] <= 8'h10 ;
			data[85968] <= 8'h10 ;
			data[85969] <= 8'h10 ;
			data[85970] <= 8'h10 ;
			data[85971] <= 8'h10 ;
			data[85972] <= 8'h10 ;
			data[85973] <= 8'h10 ;
			data[85974] <= 8'h10 ;
			data[85975] <= 8'h10 ;
			data[85976] <= 8'h10 ;
			data[85977] <= 8'h10 ;
			data[85978] <= 8'h10 ;
			data[85979] <= 8'h10 ;
			data[85980] <= 8'h10 ;
			data[85981] <= 8'h10 ;
			data[85982] <= 8'h10 ;
			data[85983] <= 8'h10 ;
			data[85984] <= 8'h10 ;
			data[85985] <= 8'h10 ;
			data[85986] <= 8'h10 ;
			data[85987] <= 8'h10 ;
			data[85988] <= 8'h10 ;
			data[85989] <= 8'h10 ;
			data[85990] <= 8'h10 ;
			data[85991] <= 8'h10 ;
			data[85992] <= 8'h10 ;
			data[85993] <= 8'h10 ;
			data[85994] <= 8'h10 ;
			data[85995] <= 8'h10 ;
			data[85996] <= 8'h10 ;
			data[85997] <= 8'h10 ;
			data[85998] <= 8'h10 ;
			data[85999] <= 8'h10 ;
			data[86000] <= 8'h10 ;
			data[86001] <= 8'h10 ;
			data[86002] <= 8'h10 ;
			data[86003] <= 8'h10 ;
			data[86004] <= 8'h10 ;
			data[86005] <= 8'h10 ;
			data[86006] <= 8'h10 ;
			data[86007] <= 8'h10 ;
			data[86008] <= 8'h10 ;
			data[86009] <= 8'h10 ;
			data[86010] <= 8'h10 ;
			data[86011] <= 8'h10 ;
			data[86012] <= 8'h10 ;
			data[86013] <= 8'h10 ;
			data[86014] <= 8'h10 ;
			data[86015] <= 8'h10 ;
			data[86016] <= 8'h10 ;
			data[86017] <= 8'h10 ;
			data[86018] <= 8'h10 ;
			data[86019] <= 8'h10 ;
			data[86020] <= 8'h10 ;
			data[86021] <= 8'h10 ;
			data[86022] <= 8'h10 ;
			data[86023] <= 8'h10 ;
			data[86024] <= 8'h10 ;
			data[86025] <= 8'h10 ;
			data[86026] <= 8'h10 ;
			data[86027] <= 8'h10 ;
			data[86028] <= 8'h10 ;
			data[86029] <= 8'h10 ;
			data[86030] <= 8'h10 ;
			data[86031] <= 8'h10 ;
			data[86032] <= 8'h10 ;
			data[86033] <= 8'h10 ;
			data[86034] <= 8'h10 ;
			data[86035] <= 8'h10 ;
			data[86036] <= 8'h10 ;
			data[86037] <= 8'h10 ;
			data[86038] <= 8'h10 ;
			data[86039] <= 8'h10 ;
			data[86040] <= 8'h10 ;
			data[86041] <= 8'h10 ;
			data[86042] <= 8'h10 ;
			data[86043] <= 8'h10 ;
			data[86044] <= 8'h10 ;
			data[86045] <= 8'h10 ;
			data[86046] <= 8'h10 ;
			data[86047] <= 8'h10 ;
			data[86048] <= 8'h10 ;
			data[86049] <= 8'h10 ;
			data[86050] <= 8'h10 ;
			data[86051] <= 8'h10 ;
			data[86052] <= 8'h10 ;
			data[86053] <= 8'h10 ;
			data[86054] <= 8'h10 ;
			data[86055] <= 8'h10 ;
			data[86056] <= 8'h10 ;
			data[86057] <= 8'h10 ;
			data[86058] <= 8'h10 ;
			data[86059] <= 8'h10 ;
			data[86060] <= 8'h10 ;
			data[86061] <= 8'h10 ;
			data[86062] <= 8'h10 ;
			data[86063] <= 8'h10 ;
			data[86064] <= 8'h10 ;
			data[86065] <= 8'h10 ;
			data[86066] <= 8'h10 ;
			data[86067] <= 8'h10 ;
			data[86068] <= 8'h10 ;
			data[86069] <= 8'h10 ;
			data[86070] <= 8'h10 ;
			data[86071] <= 8'h10 ;
			data[86072] <= 8'h10 ;
			data[86073] <= 8'h10 ;
			data[86074] <= 8'h10 ;
			data[86075] <= 8'h10 ;
			data[86076] <= 8'h10 ;
			data[86077] <= 8'h10 ;
			data[86078] <= 8'h10 ;
			data[86079] <= 8'h10 ;
			data[86080] <= 8'h10 ;
			data[86081] <= 8'h10 ;
			data[86082] <= 8'h10 ;
			data[86083] <= 8'h10 ;
			data[86084] <= 8'h10 ;
			data[86085] <= 8'h10 ;
			data[86086] <= 8'h10 ;
			data[86087] <= 8'h10 ;
			data[86088] <= 8'h10 ;
			data[86089] <= 8'h10 ;
			data[86090] <= 8'h10 ;
			data[86091] <= 8'h10 ;
			data[86092] <= 8'h10 ;
			data[86093] <= 8'h10 ;
			data[86094] <= 8'h10 ;
			data[86095] <= 8'h10 ;
			data[86096] <= 8'h10 ;
			data[86097] <= 8'h10 ;
			data[86098] <= 8'h10 ;
			data[86099] <= 8'h10 ;
			data[86100] <= 8'h10 ;
			data[86101] <= 8'h10 ;
			data[86102] <= 8'h10 ;
			data[86103] <= 8'h10 ;
			data[86104] <= 8'h10 ;
			data[86105] <= 8'h10 ;
			data[86106] <= 8'h10 ;
			data[86107] <= 8'h10 ;
			data[86108] <= 8'h10 ;
			data[86109] <= 8'h10 ;
			data[86110] <= 8'h10 ;
			data[86111] <= 8'h10 ;
			data[86112] <= 8'h10 ;
			data[86113] <= 8'h10 ;
			data[86114] <= 8'h10 ;
			data[86115] <= 8'h10 ;
			data[86116] <= 8'h10 ;
			data[86117] <= 8'h10 ;
			data[86118] <= 8'h10 ;
			data[86119] <= 8'h10 ;
			data[86120] <= 8'h10 ;
			data[86121] <= 8'h10 ;
			data[86122] <= 8'h10 ;
			data[86123] <= 8'h10 ;
			data[86124] <= 8'h10 ;
			data[86125] <= 8'h10 ;
			data[86126] <= 8'h10 ;
			data[86127] <= 8'h10 ;
			data[86128] <= 8'h10 ;
			data[86129] <= 8'h10 ;
			data[86130] <= 8'h10 ;
			data[86131] <= 8'h10 ;
			data[86132] <= 8'h10 ;
			data[86133] <= 8'h10 ;
			data[86134] <= 8'h10 ;
			data[86135] <= 8'h10 ;
			data[86136] <= 8'h10 ;
			data[86137] <= 8'h10 ;
			data[86138] <= 8'h10 ;
			data[86139] <= 8'h10 ;
			data[86140] <= 8'h10 ;
			data[86141] <= 8'h10 ;
			data[86142] <= 8'h10 ;
			data[86143] <= 8'h10 ;
			data[86144] <= 8'h10 ;
			data[86145] <= 8'h10 ;
			data[86146] <= 8'h10 ;
			data[86147] <= 8'h10 ;
			data[86148] <= 8'h10 ;
			data[86149] <= 8'h10 ;
			data[86150] <= 8'h10 ;
			data[86151] <= 8'h10 ;
			data[86152] <= 8'h10 ;
			data[86153] <= 8'h10 ;
			data[86154] <= 8'h10 ;
			data[86155] <= 8'h10 ;
			data[86156] <= 8'h10 ;
			data[86157] <= 8'h10 ;
			data[86158] <= 8'h10 ;
			data[86159] <= 8'h10 ;
			data[86160] <= 8'h10 ;
			data[86161] <= 8'h10 ;
			data[86162] <= 8'h10 ;
			data[86163] <= 8'h10 ;
			data[86164] <= 8'h10 ;
			data[86165] <= 8'h10 ;
			data[86166] <= 8'h10 ;
			data[86167] <= 8'h10 ;
			data[86168] <= 8'h10 ;
			data[86169] <= 8'h10 ;
			data[86170] <= 8'h10 ;
			data[86171] <= 8'h10 ;
			data[86172] <= 8'h10 ;
			data[86173] <= 8'h10 ;
			data[86174] <= 8'h10 ;
			data[86175] <= 8'h10 ;
			data[86176] <= 8'h10 ;
			data[86177] <= 8'h10 ;
			data[86178] <= 8'h10 ;
			data[86179] <= 8'h10 ;
			data[86180] <= 8'h10 ;
			data[86181] <= 8'h10 ;
			data[86182] <= 8'h10 ;
			data[86183] <= 8'h10 ;
			data[86184] <= 8'h10 ;
			data[86185] <= 8'h10 ;
			data[86186] <= 8'h10 ;
			data[86187] <= 8'h10 ;
			data[86188] <= 8'h10 ;
			data[86189] <= 8'h10 ;
			data[86190] <= 8'h10 ;
			data[86191] <= 8'h10 ;
			data[86192] <= 8'h10 ;
			data[86193] <= 8'h10 ;
			data[86194] <= 8'h10 ;
			data[86195] <= 8'h10 ;
			data[86196] <= 8'h10 ;
			data[86197] <= 8'h10 ;
			data[86198] <= 8'h10 ;
			data[86199] <= 8'h10 ;
			data[86200] <= 8'h10 ;
			data[86201] <= 8'h10 ;
			data[86202] <= 8'h10 ;
			data[86203] <= 8'h10 ;
			data[86204] <= 8'h10 ;
			data[86205] <= 8'h10 ;
			data[86206] <= 8'h10 ;
			data[86207] <= 8'h10 ;
			data[86208] <= 8'h10 ;
			data[86209] <= 8'h10 ;
			data[86210] <= 8'h10 ;
			data[86211] <= 8'h10 ;
			data[86212] <= 8'h10 ;
			data[86213] <= 8'h10 ;
			data[86214] <= 8'h10 ;
			data[86215] <= 8'h10 ;
			data[86216] <= 8'h10 ;
			data[86217] <= 8'h10 ;
			data[86218] <= 8'h10 ;
			data[86219] <= 8'h10 ;
			data[86220] <= 8'h10 ;
			data[86221] <= 8'h10 ;
			data[86222] <= 8'h10 ;
			data[86223] <= 8'h10 ;
			data[86224] <= 8'h10 ;
			data[86225] <= 8'h10 ;
			data[86226] <= 8'h10 ;
			data[86227] <= 8'h10 ;
			data[86228] <= 8'h10 ;
			data[86229] <= 8'h10 ;
			data[86230] <= 8'h10 ;
			data[86231] <= 8'h10 ;
			data[86232] <= 8'h10 ;
			data[86233] <= 8'h10 ;
			data[86234] <= 8'h10 ;
			data[86235] <= 8'h10 ;
			data[86236] <= 8'h10 ;
			data[86237] <= 8'h10 ;
			data[86238] <= 8'h10 ;
			data[86239] <= 8'h10 ;
			data[86240] <= 8'h10 ;
			data[86241] <= 8'h10 ;
			data[86242] <= 8'h10 ;
			data[86243] <= 8'h10 ;
			data[86244] <= 8'h10 ;
			data[86245] <= 8'h10 ;
			data[86246] <= 8'h10 ;
			data[86247] <= 8'h10 ;
			data[86248] <= 8'h10 ;
			data[86249] <= 8'h10 ;
			data[86250] <= 8'h10 ;
			data[86251] <= 8'h10 ;
			data[86252] <= 8'h10 ;
			data[86253] <= 8'h10 ;
			data[86254] <= 8'h10 ;
			data[86255] <= 8'h10 ;
			data[86256] <= 8'h10 ;
			data[86257] <= 8'h10 ;
			data[86258] <= 8'h10 ;
			data[86259] <= 8'h10 ;
			data[86260] <= 8'h10 ;
			data[86261] <= 8'h10 ;
			data[86262] <= 8'h10 ;
			data[86263] <= 8'h10 ;
			data[86264] <= 8'h10 ;
			data[86265] <= 8'h10 ;
			data[86266] <= 8'h10 ;
			data[86267] <= 8'h10 ;
			data[86268] <= 8'h10 ;
			data[86269] <= 8'h10 ;
			data[86270] <= 8'h10 ;
			data[86271] <= 8'h10 ;
			data[86272] <= 8'h10 ;
			data[86273] <= 8'h10 ;
			data[86274] <= 8'h10 ;
			data[86275] <= 8'h10 ;
			data[86276] <= 8'h10 ;
			data[86277] <= 8'h10 ;
			data[86278] <= 8'h10 ;
			data[86279] <= 8'h10 ;
			data[86280] <= 8'h10 ;
			data[86281] <= 8'h10 ;
			data[86282] <= 8'h10 ;
			data[86283] <= 8'h10 ;
			data[86284] <= 8'h10 ;
			data[86285] <= 8'h10 ;
			data[86286] <= 8'h10 ;
			data[86287] <= 8'h10 ;
			data[86288] <= 8'h10 ;
			data[86289] <= 8'h10 ;
			data[86290] <= 8'h10 ;
			data[86291] <= 8'h10 ;
			data[86292] <= 8'h10 ;
			data[86293] <= 8'h10 ;
			data[86294] <= 8'h10 ;
			data[86295] <= 8'h10 ;
			data[86296] <= 8'h10 ;
			data[86297] <= 8'h10 ;
			data[86298] <= 8'h10 ;
			data[86299] <= 8'h10 ;
			data[86300] <= 8'h10 ;
			data[86301] <= 8'h10 ;
			data[86302] <= 8'h10 ;
			data[86303] <= 8'h10 ;
			data[86304] <= 8'h10 ;
			data[86305] <= 8'h10 ;
			data[86306] <= 8'h10 ;
			data[86307] <= 8'h10 ;
			data[86308] <= 8'h10 ;
			data[86309] <= 8'h10 ;
			data[86310] <= 8'h10 ;
			data[86311] <= 8'h10 ;
			data[86312] <= 8'h10 ;
			data[86313] <= 8'h10 ;
			data[86314] <= 8'h10 ;
			data[86315] <= 8'h10 ;
			data[86316] <= 8'h10 ;
			data[86317] <= 8'h10 ;
			data[86318] <= 8'h10 ;
			data[86319] <= 8'h10 ;
			data[86320] <= 8'h10 ;
			data[86321] <= 8'h10 ;
			data[86322] <= 8'h10 ;
			data[86323] <= 8'h10 ;
			data[86324] <= 8'h10 ;
			data[86325] <= 8'h10 ;
			data[86326] <= 8'h10 ;
			data[86327] <= 8'h10 ;
			data[86328] <= 8'h10 ;
			data[86329] <= 8'h10 ;
			data[86330] <= 8'h10 ;
			data[86331] <= 8'h10 ;
			data[86332] <= 8'h10 ;
			data[86333] <= 8'h10 ;
			data[86334] <= 8'h10 ;
			data[86335] <= 8'h10 ;
			data[86336] <= 8'h10 ;
			data[86337] <= 8'h10 ;
			data[86338] <= 8'h10 ;
			data[86339] <= 8'h10 ;
			data[86340] <= 8'h10 ;
			data[86341] <= 8'h10 ;
			data[86342] <= 8'h10 ;
			data[86343] <= 8'h10 ;
			data[86344] <= 8'h10 ;
			data[86345] <= 8'h10 ;
			data[86346] <= 8'h10 ;
			data[86347] <= 8'h10 ;
			data[86348] <= 8'h10 ;
			data[86349] <= 8'h10 ;
			data[86350] <= 8'h10 ;
			data[86351] <= 8'h10 ;
			data[86352] <= 8'h10 ;
			data[86353] <= 8'h10 ;
			data[86354] <= 8'h10 ;
			data[86355] <= 8'h10 ;
			data[86356] <= 8'h10 ;
			data[86357] <= 8'h10 ;
			data[86358] <= 8'h10 ;
			data[86359] <= 8'h10 ;
			data[86360] <= 8'h10 ;
			data[86361] <= 8'h10 ;
			data[86362] <= 8'h10 ;
			data[86363] <= 8'h10 ;
			data[86364] <= 8'h10 ;
			data[86365] <= 8'h10 ;
			data[86366] <= 8'h10 ;
			data[86367] <= 8'h10 ;
			data[86368] <= 8'h10 ;
			data[86369] <= 8'h10 ;
			data[86370] <= 8'h10 ;
			data[86371] <= 8'h10 ;
			data[86372] <= 8'h10 ;
			data[86373] <= 8'h10 ;
			data[86374] <= 8'h10 ;
			data[86375] <= 8'h10 ;
			data[86376] <= 8'h10 ;
			data[86377] <= 8'h10 ;
			data[86378] <= 8'h10 ;
			data[86379] <= 8'h10 ;
			data[86380] <= 8'h10 ;
			data[86381] <= 8'h10 ;
			data[86382] <= 8'h10 ;
			data[86383] <= 8'h10 ;
			data[86384] <= 8'h10 ;
			data[86385] <= 8'h10 ;
			data[86386] <= 8'h10 ;
			data[86387] <= 8'h10 ;
			data[86388] <= 8'h10 ;
			data[86389] <= 8'h10 ;
			data[86390] <= 8'h10 ;
			data[86391] <= 8'h10 ;
			data[86392] <= 8'h10 ;
			data[86393] <= 8'h10 ;
			data[86394] <= 8'h10 ;
			data[86395] <= 8'h10 ;
			data[86396] <= 8'h10 ;
			data[86397] <= 8'h10 ;
			data[86398] <= 8'h10 ;
			data[86399] <= 8'h10 ;
			data[86400] <= 8'h10 ;
			data[86401] <= 8'h10 ;
			data[86402] <= 8'h10 ;
			data[86403] <= 8'h10 ;
			data[86404] <= 8'h10 ;
			data[86405] <= 8'h10 ;
			data[86406] <= 8'h10 ;
			data[86407] <= 8'h10 ;
			data[86408] <= 8'h10 ;
			data[86409] <= 8'h10 ;
			data[86410] <= 8'h10 ;
			data[86411] <= 8'h10 ;
			data[86412] <= 8'h10 ;
			data[86413] <= 8'h10 ;
			data[86414] <= 8'h10 ;
			data[86415] <= 8'h10 ;
			data[86416] <= 8'h10 ;
			data[86417] <= 8'h10 ;
			data[86418] <= 8'h10 ;
			data[86419] <= 8'h10 ;
			data[86420] <= 8'h10 ;
			data[86421] <= 8'h10 ;
			data[86422] <= 8'h10 ;
			data[86423] <= 8'h10 ;
			data[86424] <= 8'h10 ;
			data[86425] <= 8'h10 ;
			data[86426] <= 8'h10 ;
			data[86427] <= 8'h10 ;
			data[86428] <= 8'h10 ;
			data[86429] <= 8'h10 ;
			data[86430] <= 8'h10 ;
			data[86431] <= 8'h10 ;
			data[86432] <= 8'h10 ;
			data[86433] <= 8'h10 ;
			data[86434] <= 8'h10 ;
			data[86435] <= 8'h10 ;
			data[86436] <= 8'h10 ;
			data[86437] <= 8'h10 ;
			data[86438] <= 8'h10 ;
			data[86439] <= 8'h10 ;
			data[86440] <= 8'h10 ;
			data[86441] <= 8'h10 ;
			data[86442] <= 8'h10 ;
			data[86443] <= 8'h10 ;
			data[86444] <= 8'h10 ;
			data[86445] <= 8'h10 ;
			data[86446] <= 8'h10 ;
			data[86447] <= 8'h10 ;
			data[86448] <= 8'h10 ;
			data[86449] <= 8'h10 ;
			data[86450] <= 8'h10 ;
			data[86451] <= 8'h10 ;
			data[86452] <= 8'h10 ;
			data[86453] <= 8'h10 ;
			data[86454] <= 8'h10 ;
			data[86455] <= 8'h10 ;
			data[86456] <= 8'h10 ;
			data[86457] <= 8'h10 ;
			data[86458] <= 8'h10 ;
			data[86459] <= 8'h10 ;
			data[86460] <= 8'h10 ;
			data[86461] <= 8'h10 ;
			data[86462] <= 8'h10 ;
			data[86463] <= 8'h10 ;
			data[86464] <= 8'h10 ;
			data[86465] <= 8'h10 ;
			data[86466] <= 8'h10 ;
			data[86467] <= 8'h10 ;
			data[86468] <= 8'h10 ;
			data[86469] <= 8'h10 ;
			data[86470] <= 8'h10 ;
			data[86471] <= 8'h10 ;
			data[86472] <= 8'h10 ;
			data[86473] <= 8'h10 ;
			data[86474] <= 8'h10 ;
			data[86475] <= 8'h10 ;
			data[86476] <= 8'h10 ;
			data[86477] <= 8'h10 ;
			data[86478] <= 8'h10 ;
			data[86479] <= 8'h10 ;
			data[86480] <= 8'h10 ;
			data[86481] <= 8'h10 ;
			data[86482] <= 8'h10 ;
			data[86483] <= 8'h10 ;
			data[86484] <= 8'h10 ;
			data[86485] <= 8'h10 ;
			data[86486] <= 8'h10 ;
			data[86487] <= 8'h10 ;
			data[86488] <= 8'h10 ;
			data[86489] <= 8'h10 ;
			data[86490] <= 8'h10 ;
			data[86491] <= 8'h10 ;
			data[86492] <= 8'h10 ;
			data[86493] <= 8'h10 ;
			data[86494] <= 8'h10 ;
			data[86495] <= 8'h10 ;
			data[86496] <= 8'h10 ;
			data[86497] <= 8'h10 ;
			data[86498] <= 8'h10 ;
			data[86499] <= 8'h10 ;
			data[86500] <= 8'h10 ;
			data[86501] <= 8'h10 ;
			data[86502] <= 8'h10 ;
			data[86503] <= 8'h10 ;
			data[86504] <= 8'h10 ;
			data[86505] <= 8'h10 ;
			data[86506] <= 8'h10 ;
			data[86507] <= 8'h10 ;
			data[86508] <= 8'h10 ;
			data[86509] <= 8'h10 ;
			data[86510] <= 8'h10 ;
			data[86511] <= 8'h10 ;
			data[86512] <= 8'h10 ;
			data[86513] <= 8'h10 ;
			data[86514] <= 8'h10 ;
			data[86515] <= 8'h10 ;
			data[86516] <= 8'h10 ;
			data[86517] <= 8'h10 ;
			data[86518] <= 8'h10 ;
			data[86519] <= 8'h10 ;
			data[86520] <= 8'h10 ;
			data[86521] <= 8'h10 ;
			data[86522] <= 8'h10 ;
			data[86523] <= 8'h10 ;
			data[86524] <= 8'h10 ;
			data[86525] <= 8'h10 ;
			data[86526] <= 8'h10 ;
			data[86527] <= 8'h10 ;
			data[86528] <= 8'h10 ;
			data[86529] <= 8'h10 ;
			data[86530] <= 8'h10 ;
			data[86531] <= 8'h10 ;
			data[86532] <= 8'h10 ;
			data[86533] <= 8'h10 ;
			data[86534] <= 8'h10 ;
			data[86535] <= 8'h10 ;
			data[86536] <= 8'h10 ;
			data[86537] <= 8'h10 ;
			data[86538] <= 8'h10 ;
			data[86539] <= 8'h10 ;
			data[86540] <= 8'h10 ;
			data[86541] <= 8'h10 ;
			data[86542] <= 8'h10 ;
			data[86543] <= 8'h10 ;
			data[86544] <= 8'h10 ;
			data[86545] <= 8'h10 ;
			data[86546] <= 8'h10 ;
			data[86547] <= 8'h10 ;
			data[86548] <= 8'h10 ;
			data[86549] <= 8'h10 ;
			data[86550] <= 8'h10 ;
			data[86551] <= 8'h10 ;
			data[86552] <= 8'h10 ;
			data[86553] <= 8'h10 ;
			data[86554] <= 8'h10 ;
			data[86555] <= 8'h10 ;
			data[86556] <= 8'h10 ;
			data[86557] <= 8'h10 ;
			data[86558] <= 8'h10 ;
			data[86559] <= 8'h10 ;
			data[86560] <= 8'h10 ;
			data[86561] <= 8'h10 ;
			data[86562] <= 8'h10 ;
			data[86563] <= 8'h10 ;
			data[86564] <= 8'h10 ;
			data[86565] <= 8'h10 ;
			data[86566] <= 8'h10 ;
			data[86567] <= 8'h10 ;
			data[86568] <= 8'h10 ;
			data[86569] <= 8'h10 ;
			data[86570] <= 8'h10 ;
			data[86571] <= 8'h10 ;
			data[86572] <= 8'h10 ;
			data[86573] <= 8'h10 ;
			data[86574] <= 8'h10 ;
			data[86575] <= 8'h10 ;
			data[86576] <= 8'h10 ;
			data[86577] <= 8'h10 ;
			data[86578] <= 8'h10 ;
			data[86579] <= 8'h10 ;
			data[86580] <= 8'h10 ;
			data[86581] <= 8'h10 ;
			data[86582] <= 8'h10 ;
			data[86583] <= 8'h10 ;
			data[86584] <= 8'h10 ;
			data[86585] <= 8'h10 ;
			data[86586] <= 8'h10 ;
			data[86587] <= 8'h10 ;
			data[86588] <= 8'h10 ;
			data[86589] <= 8'h10 ;
			data[86590] <= 8'h10 ;
			data[86591] <= 8'h10 ;
			data[86592] <= 8'h10 ;
			data[86593] <= 8'h10 ;
			data[86594] <= 8'h10 ;
			data[86595] <= 8'h10 ;
			data[86596] <= 8'h10 ;
			data[86597] <= 8'h10 ;
			data[86598] <= 8'h10 ;
			data[86599] <= 8'h10 ;
			data[86600] <= 8'h10 ;
			data[86601] <= 8'h10 ;
			data[86602] <= 8'h10 ;
			data[86603] <= 8'h10 ;
			data[86604] <= 8'h10 ;
			data[86605] <= 8'h10 ;
			data[86606] <= 8'h10 ;
			data[86607] <= 8'h10 ;
			data[86608] <= 8'h10 ;
			data[86609] <= 8'h10 ;
			data[86610] <= 8'h10 ;
			data[86611] <= 8'h10 ;
			data[86612] <= 8'h10 ;
			data[86613] <= 8'h10 ;
			data[86614] <= 8'h10 ;
			data[86615] <= 8'h10 ;
			data[86616] <= 8'h10 ;
			data[86617] <= 8'h10 ;
			data[86618] <= 8'h10 ;
			data[86619] <= 8'h10 ;
			data[86620] <= 8'h10 ;
			data[86621] <= 8'h10 ;
			data[86622] <= 8'h10 ;
			data[86623] <= 8'h10 ;
			data[86624] <= 8'h10 ;
			data[86625] <= 8'h10 ;
			data[86626] <= 8'h10 ;
			data[86627] <= 8'h10 ;
			data[86628] <= 8'h10 ;
			data[86629] <= 8'h10 ;
			data[86630] <= 8'h10 ;
			data[86631] <= 8'h10 ;
			data[86632] <= 8'h10 ;
			data[86633] <= 8'h10 ;
			data[86634] <= 8'h10 ;
			data[86635] <= 8'h10 ;
			data[86636] <= 8'h10 ;
			data[86637] <= 8'h10 ;
			data[86638] <= 8'h10 ;
			data[86639] <= 8'h10 ;
			data[86640] <= 8'h10 ;
			data[86641] <= 8'h10 ;
			data[86642] <= 8'h10 ;
			data[86643] <= 8'h10 ;
			data[86644] <= 8'h10 ;
			data[86645] <= 8'h10 ;
			data[86646] <= 8'h10 ;
			data[86647] <= 8'h10 ;
			data[86648] <= 8'h10 ;
			data[86649] <= 8'h10 ;
			data[86650] <= 8'h10 ;
			data[86651] <= 8'h10 ;
			data[86652] <= 8'h10 ;
			data[86653] <= 8'h10 ;
			data[86654] <= 8'h10 ;
			data[86655] <= 8'h10 ;
			data[86656] <= 8'h10 ;
			data[86657] <= 8'h10 ;
			data[86658] <= 8'h10 ;
			data[86659] <= 8'h10 ;
			data[86660] <= 8'h10 ;
			data[86661] <= 8'h10 ;
			data[86662] <= 8'h10 ;
			data[86663] <= 8'h10 ;
			data[86664] <= 8'h10 ;
			data[86665] <= 8'h10 ;
			data[86666] <= 8'h10 ;
			data[86667] <= 8'h10 ;
			data[86668] <= 8'h10 ;
			data[86669] <= 8'h10 ;
			data[86670] <= 8'h10 ;
			data[86671] <= 8'h10 ;
			data[86672] <= 8'h10 ;
			data[86673] <= 8'h10 ;
			data[86674] <= 8'h10 ;
			data[86675] <= 8'h10 ;
			data[86676] <= 8'h10 ;
			data[86677] <= 8'h10 ;
			data[86678] <= 8'h10 ;
			data[86679] <= 8'h10 ;
			data[86680] <= 8'h10 ;
			data[86681] <= 8'h10 ;
			data[86682] <= 8'h10 ;
			data[86683] <= 8'h10 ;
			data[86684] <= 8'h10 ;
			data[86685] <= 8'h10 ;
			data[86686] <= 8'h10 ;
			data[86687] <= 8'h10 ;
			data[86688] <= 8'h10 ;
			data[86689] <= 8'h10 ;
			data[86690] <= 8'h10 ;
			data[86691] <= 8'h10 ;
			data[86692] <= 8'h10 ;
			data[86693] <= 8'h10 ;
			data[86694] <= 8'h10 ;
			data[86695] <= 8'h10 ;
			data[86696] <= 8'h10 ;
			data[86697] <= 8'h10 ;
			data[86698] <= 8'h10 ;
			data[86699] <= 8'h10 ;
			data[86700] <= 8'h10 ;
			data[86701] <= 8'h10 ;
			data[86702] <= 8'h10 ;
			data[86703] <= 8'h10 ;
			data[86704] <= 8'h10 ;
			data[86705] <= 8'h10 ;
			data[86706] <= 8'h10 ;
			data[86707] <= 8'h10 ;
			data[86708] <= 8'h10 ;
			data[86709] <= 8'h10 ;
			data[86710] <= 8'h10 ;
			data[86711] <= 8'h10 ;
			data[86712] <= 8'h10 ;
			data[86713] <= 8'h10 ;
			data[86714] <= 8'h10 ;
			data[86715] <= 8'h10 ;
			data[86716] <= 8'h10 ;
			data[86717] <= 8'h10 ;
			data[86718] <= 8'h10 ;
			data[86719] <= 8'h10 ;
			data[86720] <= 8'h10 ;
			data[86721] <= 8'h10 ;
			data[86722] <= 8'h10 ;
			data[86723] <= 8'h10 ;
			data[86724] <= 8'h10 ;
			data[86725] <= 8'h10 ;
			data[86726] <= 8'h10 ;
			data[86727] <= 8'h10 ;
			data[86728] <= 8'h10 ;
			data[86729] <= 8'h10 ;
			data[86730] <= 8'h10 ;
			data[86731] <= 8'h10 ;
			data[86732] <= 8'h10 ;
			data[86733] <= 8'h10 ;
			data[86734] <= 8'h10 ;
			data[86735] <= 8'h10 ;
			data[86736] <= 8'h10 ;
			data[86737] <= 8'h10 ;
			data[86738] <= 8'h10 ;
			data[86739] <= 8'h10 ;
			data[86740] <= 8'h10 ;
			data[86741] <= 8'h10 ;
			data[86742] <= 8'h10 ;
			data[86743] <= 8'h10 ;
			data[86744] <= 8'h10 ;
			data[86745] <= 8'h10 ;
			data[86746] <= 8'h10 ;
			data[86747] <= 8'h10 ;
			data[86748] <= 8'h10 ;
			data[86749] <= 8'h10 ;
			data[86750] <= 8'h10 ;
			data[86751] <= 8'h10 ;
			data[86752] <= 8'h10 ;
			data[86753] <= 8'h10 ;
			data[86754] <= 8'h10 ;
			data[86755] <= 8'h10 ;
			data[86756] <= 8'h10 ;
			data[86757] <= 8'h10 ;
			data[86758] <= 8'h10 ;
			data[86759] <= 8'h10 ;
			data[86760] <= 8'h10 ;
			data[86761] <= 8'h10 ;
			data[86762] <= 8'h10 ;
			data[86763] <= 8'h10 ;
			data[86764] <= 8'h10 ;
			data[86765] <= 8'h10 ;
			data[86766] <= 8'h10 ;
			data[86767] <= 8'h10 ;
			data[86768] <= 8'h10 ;
			data[86769] <= 8'h10 ;
			data[86770] <= 8'h10 ;
			data[86771] <= 8'h10 ;
			data[86772] <= 8'h10 ;
			data[86773] <= 8'h10 ;
			data[86774] <= 8'h10 ;
			data[86775] <= 8'h10 ;
			data[86776] <= 8'h10 ;
			data[86777] <= 8'h10 ;
			data[86778] <= 8'h10 ;
			data[86779] <= 8'h10 ;
			data[86780] <= 8'h10 ;
			data[86781] <= 8'h10 ;
			data[86782] <= 8'h10 ;
			data[86783] <= 8'h10 ;
			data[86784] <= 8'h10 ;
			data[86785] <= 8'h10 ;
			data[86786] <= 8'h10 ;
			data[86787] <= 8'h10 ;
			data[86788] <= 8'h10 ;
			data[86789] <= 8'h10 ;
			data[86790] <= 8'h10 ;
			data[86791] <= 8'h10 ;
			data[86792] <= 8'h10 ;
			data[86793] <= 8'h10 ;
			data[86794] <= 8'h10 ;
			data[86795] <= 8'h10 ;
			data[86796] <= 8'h10 ;
			data[86797] <= 8'h10 ;
			data[86798] <= 8'h10 ;
			data[86799] <= 8'h10 ;
			data[86800] <= 8'h10 ;
			data[86801] <= 8'h10 ;
			data[86802] <= 8'h10 ;
			data[86803] <= 8'h10 ;
			data[86804] <= 8'h10 ;
			data[86805] <= 8'h10 ;
			data[86806] <= 8'h10 ;
			data[86807] <= 8'h10 ;
			data[86808] <= 8'h10 ;
			data[86809] <= 8'h10 ;
			data[86810] <= 8'h10 ;
			data[86811] <= 8'h10 ;
			data[86812] <= 8'h10 ;
			data[86813] <= 8'h10 ;
			data[86814] <= 8'h10 ;
			data[86815] <= 8'h10 ;
			data[86816] <= 8'h10 ;
			data[86817] <= 8'h10 ;
			data[86818] <= 8'h10 ;
			data[86819] <= 8'h10 ;
			data[86820] <= 8'h10 ;
			data[86821] <= 8'h10 ;
			data[86822] <= 8'h10 ;
			data[86823] <= 8'h10 ;
			data[86824] <= 8'h10 ;
			data[86825] <= 8'h10 ;
			data[86826] <= 8'h10 ;
			data[86827] <= 8'h10 ;
			data[86828] <= 8'h10 ;
			data[86829] <= 8'h10 ;
			data[86830] <= 8'h10 ;
			data[86831] <= 8'h10 ;
			data[86832] <= 8'h10 ;
			data[86833] <= 8'h10 ;
			data[86834] <= 8'h10 ;
			data[86835] <= 8'h10 ;
			data[86836] <= 8'h10 ;
			data[86837] <= 8'h10 ;
			data[86838] <= 8'h10 ;
			data[86839] <= 8'h10 ;
			data[86840] <= 8'h10 ;
			data[86841] <= 8'h10 ;
			data[86842] <= 8'h10 ;
			data[86843] <= 8'h10 ;
			data[86844] <= 8'h10 ;
			data[86845] <= 8'h10 ;
			data[86846] <= 8'h10 ;
			data[86847] <= 8'h10 ;
			data[86848] <= 8'h10 ;
			data[86849] <= 8'h10 ;
			data[86850] <= 8'h10 ;
			data[86851] <= 8'h10 ;
			data[86852] <= 8'h10 ;
			data[86853] <= 8'h10 ;
			data[86854] <= 8'h10 ;
			data[86855] <= 8'h10 ;
			data[86856] <= 8'h10 ;
			data[86857] <= 8'h10 ;
			data[86858] <= 8'h10 ;
			data[86859] <= 8'h10 ;
			data[86860] <= 8'h10 ;
			data[86861] <= 8'h10 ;
			data[86862] <= 8'h10 ;
			data[86863] <= 8'h10 ;
			data[86864] <= 8'h10 ;
			data[86865] <= 8'h10 ;
			data[86866] <= 8'h10 ;
			data[86867] <= 8'h10 ;
			data[86868] <= 8'h10 ;
			data[86869] <= 8'h10 ;
			data[86870] <= 8'h10 ;
			data[86871] <= 8'h10 ;
			data[86872] <= 8'h10 ;
			data[86873] <= 8'h10 ;
			data[86874] <= 8'h10 ;
			data[86875] <= 8'h10 ;
			data[86876] <= 8'h10 ;
			data[86877] <= 8'h10 ;
			data[86878] <= 8'h10 ;
			data[86879] <= 8'h10 ;
			data[86880] <= 8'h10 ;
			data[86881] <= 8'h10 ;
			data[86882] <= 8'h10 ;
			data[86883] <= 8'h10 ;
			data[86884] <= 8'h10 ;
			data[86885] <= 8'h10 ;
			data[86886] <= 8'h10 ;
			data[86887] <= 8'h10 ;
			data[86888] <= 8'h10 ;
			data[86889] <= 8'h10 ;
			data[86890] <= 8'h10 ;
			data[86891] <= 8'h10 ;
			data[86892] <= 8'h10 ;
			data[86893] <= 8'h10 ;
			data[86894] <= 8'h10 ;
			data[86895] <= 8'h10 ;
			data[86896] <= 8'h10 ;
			data[86897] <= 8'h10 ;
			data[86898] <= 8'h10 ;
			data[86899] <= 8'h10 ;
			data[86900] <= 8'h10 ;
			data[86901] <= 8'h10 ;
			data[86902] <= 8'h10 ;
			data[86903] <= 8'h10 ;
			data[86904] <= 8'h10 ;
			data[86905] <= 8'h10 ;
			data[86906] <= 8'h10 ;
			data[86907] <= 8'h10 ;
			data[86908] <= 8'h10 ;
			data[86909] <= 8'h10 ;
			data[86910] <= 8'h10 ;
			data[86911] <= 8'h10 ;
			data[86912] <= 8'h10 ;
			data[86913] <= 8'h10 ;
			data[86914] <= 8'h10 ;
			data[86915] <= 8'h10 ;
			data[86916] <= 8'h10 ;
			data[86917] <= 8'h10 ;
			data[86918] <= 8'h10 ;
			data[86919] <= 8'h10 ;
			data[86920] <= 8'h10 ;
			data[86921] <= 8'h10 ;
			data[86922] <= 8'h10 ;
			data[86923] <= 8'h10 ;
			data[86924] <= 8'h10 ;
			data[86925] <= 8'h10 ;
			data[86926] <= 8'h10 ;
			data[86927] <= 8'h10 ;
			data[86928] <= 8'h10 ;
			data[86929] <= 8'h10 ;
			data[86930] <= 8'h10 ;
			data[86931] <= 8'h10 ;
			data[86932] <= 8'h10 ;
			data[86933] <= 8'h10 ;
			data[86934] <= 8'h10 ;
			data[86935] <= 8'h10 ;
			data[86936] <= 8'h10 ;
			data[86937] <= 8'h10 ;
			data[86938] <= 8'h10 ;
			data[86939] <= 8'h10 ;
			data[86940] <= 8'h10 ;
			data[86941] <= 8'h10 ;
			data[86942] <= 8'h10 ;
			data[86943] <= 8'h10 ;
			data[86944] <= 8'h10 ;
			data[86945] <= 8'h10 ;
			data[86946] <= 8'h10 ;
			data[86947] <= 8'h10 ;
			data[86948] <= 8'h10 ;
			data[86949] <= 8'h10 ;
			data[86950] <= 8'h10 ;
			data[86951] <= 8'h10 ;
			data[86952] <= 8'h10 ;
			data[86953] <= 8'h10 ;
			data[86954] <= 8'h10 ;
			data[86955] <= 8'h10 ;
			data[86956] <= 8'h10 ;
			data[86957] <= 8'h10 ;
			data[86958] <= 8'h10 ;
			data[86959] <= 8'h10 ;
			data[86960] <= 8'h10 ;
			data[86961] <= 8'h10 ;
			data[86962] <= 8'h10 ;
			data[86963] <= 8'h10 ;
			data[86964] <= 8'h10 ;
			data[86965] <= 8'h10 ;
			data[86966] <= 8'h10 ;
			data[86967] <= 8'h10 ;
			data[86968] <= 8'h10 ;
			data[86969] <= 8'h10 ;
			data[86970] <= 8'h10 ;
			data[86971] <= 8'h10 ;
			data[86972] <= 8'h10 ;
			data[86973] <= 8'h10 ;
			data[86974] <= 8'h10 ;
			data[86975] <= 8'h10 ;
			data[86976] <= 8'h10 ;
			data[86977] <= 8'h10 ;
			data[86978] <= 8'h10 ;
			data[86979] <= 8'h10 ;
			data[86980] <= 8'h10 ;
			data[86981] <= 8'h10 ;
			data[86982] <= 8'h10 ;
			data[86983] <= 8'h10 ;
			data[86984] <= 8'h10 ;
			data[86985] <= 8'h10 ;
			data[86986] <= 8'h10 ;
			data[86987] <= 8'h10 ;
			data[86988] <= 8'h10 ;
			data[86989] <= 8'h10 ;
			data[86990] <= 8'h10 ;
			data[86991] <= 8'h10 ;
			data[86992] <= 8'h10 ;
			data[86993] <= 8'h10 ;
			data[86994] <= 8'h10 ;
			data[86995] <= 8'h10 ;
			data[86996] <= 8'h10 ;
			data[86997] <= 8'h10 ;
			data[86998] <= 8'h10 ;
			data[86999] <= 8'h10 ;
			data[87000] <= 8'h10 ;
			data[87001] <= 8'h10 ;
			data[87002] <= 8'h10 ;
			data[87003] <= 8'h10 ;
			data[87004] <= 8'h10 ;
			data[87005] <= 8'h10 ;
			data[87006] <= 8'h10 ;
			data[87007] <= 8'h10 ;
			data[87008] <= 8'h10 ;
			data[87009] <= 8'h10 ;
			data[87010] <= 8'h10 ;
			data[87011] <= 8'h10 ;
			data[87012] <= 8'h10 ;
			data[87013] <= 8'h10 ;
			data[87014] <= 8'h10 ;
			data[87015] <= 8'h10 ;
			data[87016] <= 8'h10 ;
			data[87017] <= 8'h10 ;
			data[87018] <= 8'h10 ;
			data[87019] <= 8'h10 ;
			data[87020] <= 8'h10 ;
			data[87021] <= 8'h10 ;
			data[87022] <= 8'h10 ;
			data[87023] <= 8'h10 ;
			data[87024] <= 8'h10 ;
			data[87025] <= 8'h10 ;
			data[87026] <= 8'h10 ;
			data[87027] <= 8'h10 ;
			data[87028] <= 8'h10 ;
			data[87029] <= 8'h10 ;
			data[87030] <= 8'h10 ;
			data[87031] <= 8'h10 ;
			data[87032] <= 8'h10 ;
			data[87033] <= 8'h10 ;
			data[87034] <= 8'h10 ;
			data[87035] <= 8'h10 ;
			data[87036] <= 8'h10 ;
			data[87037] <= 8'h10 ;
			data[87038] <= 8'h10 ;
			data[87039] <= 8'h10 ;
			data[87040] <= 8'h10 ;
			data[87041] <= 8'h10 ;
			data[87042] <= 8'h10 ;
			data[87043] <= 8'h10 ;
			data[87044] <= 8'h10 ;
			data[87045] <= 8'h10 ;
			data[87046] <= 8'h10 ;
			data[87047] <= 8'h10 ;
			data[87048] <= 8'h10 ;
			data[87049] <= 8'h10 ;
			data[87050] <= 8'h10 ;
			data[87051] <= 8'h10 ;
			data[87052] <= 8'h10 ;
			data[87053] <= 8'h10 ;
			data[87054] <= 8'h10 ;
			data[87055] <= 8'h10 ;
			data[87056] <= 8'h10 ;
			data[87057] <= 8'h10 ;
			data[87058] <= 8'h10 ;
			data[87059] <= 8'h10 ;
			data[87060] <= 8'h10 ;
			data[87061] <= 8'h10 ;
			data[87062] <= 8'h10 ;
			data[87063] <= 8'h10 ;
			data[87064] <= 8'h10 ;
			data[87065] <= 8'h10 ;
			data[87066] <= 8'h10 ;
			data[87067] <= 8'h10 ;
			data[87068] <= 8'h10 ;
			data[87069] <= 8'h10 ;
			data[87070] <= 8'h10 ;
			data[87071] <= 8'h10 ;
			data[87072] <= 8'h10 ;
			data[87073] <= 8'h10 ;
			data[87074] <= 8'h10 ;
			data[87075] <= 8'h10 ;
			data[87076] <= 8'h10 ;
			data[87077] <= 8'h10 ;
			data[87078] <= 8'h10 ;
			data[87079] <= 8'h10 ;
			data[87080] <= 8'h10 ;
			data[87081] <= 8'h10 ;
			data[87082] <= 8'h10 ;
			data[87083] <= 8'h10 ;
			data[87084] <= 8'h10 ;
			data[87085] <= 8'h10 ;
			data[87086] <= 8'h10 ;
			data[87087] <= 8'h10 ;
			data[87088] <= 8'h10 ;
			data[87089] <= 8'h10 ;
			data[87090] <= 8'h10 ;
			data[87091] <= 8'h10 ;
			data[87092] <= 8'h10 ;
			data[87093] <= 8'h10 ;
			data[87094] <= 8'h10 ;
			data[87095] <= 8'h10 ;
			data[87096] <= 8'h10 ;
			data[87097] <= 8'h10 ;
			data[87098] <= 8'h10 ;
			data[87099] <= 8'h10 ;
			data[87100] <= 8'h10 ;
			data[87101] <= 8'h10 ;
			data[87102] <= 8'h10 ;
			data[87103] <= 8'h10 ;
			data[87104] <= 8'h10 ;
			data[87105] <= 8'h10 ;
			data[87106] <= 8'h10 ;
			data[87107] <= 8'h10 ;
			data[87108] <= 8'h10 ;
			data[87109] <= 8'h10 ;
			data[87110] <= 8'h10 ;
			data[87111] <= 8'h10 ;
			data[87112] <= 8'h10 ;
			data[87113] <= 8'h10 ;
			data[87114] <= 8'h10 ;
			data[87115] <= 8'h10 ;
			data[87116] <= 8'h10 ;
			data[87117] <= 8'h10 ;
			data[87118] <= 8'h10 ;
			data[87119] <= 8'h10 ;
			data[87120] <= 8'h10 ;
			data[87121] <= 8'h10 ;
			data[87122] <= 8'h10 ;
			data[87123] <= 8'h10 ;
			data[87124] <= 8'h10 ;
			data[87125] <= 8'h10 ;
			data[87126] <= 8'h10 ;
			data[87127] <= 8'h10 ;
			data[87128] <= 8'h10 ;
			data[87129] <= 8'h10 ;
			data[87130] <= 8'h10 ;
			data[87131] <= 8'h10 ;
			data[87132] <= 8'h10 ;
			data[87133] <= 8'h10 ;
			data[87134] <= 8'h10 ;
			data[87135] <= 8'h10 ;
			data[87136] <= 8'h10 ;
			data[87137] <= 8'h10 ;
			data[87138] <= 8'h10 ;
			data[87139] <= 8'h10 ;
			data[87140] <= 8'h10 ;
			data[87141] <= 8'h10 ;
			data[87142] <= 8'h10 ;
			data[87143] <= 8'h10 ;
			data[87144] <= 8'h10 ;
			data[87145] <= 8'h10 ;
			data[87146] <= 8'h10 ;
			data[87147] <= 8'h10 ;
			data[87148] <= 8'h10 ;
			data[87149] <= 8'h10 ;
			data[87150] <= 8'h10 ;
			data[87151] <= 8'h10 ;
			data[87152] <= 8'h10 ;
			data[87153] <= 8'h10 ;
			data[87154] <= 8'h10 ;
			data[87155] <= 8'h10 ;
			data[87156] <= 8'h10 ;
			data[87157] <= 8'h10 ;
			data[87158] <= 8'h10 ;
			data[87159] <= 8'h10 ;
			data[87160] <= 8'h10 ;
			data[87161] <= 8'h10 ;
			data[87162] <= 8'h10 ;
			data[87163] <= 8'h10 ;
			data[87164] <= 8'h10 ;
			data[87165] <= 8'h10 ;
			data[87166] <= 8'h10 ;
			data[87167] <= 8'h10 ;
			data[87168] <= 8'h10 ;
			data[87169] <= 8'h10 ;
			data[87170] <= 8'h10 ;
			data[87171] <= 8'h10 ;
			data[87172] <= 8'h10 ;
			data[87173] <= 8'h10 ;
			data[87174] <= 8'h10 ;
			data[87175] <= 8'h10 ;
			data[87176] <= 8'h10 ;
			data[87177] <= 8'h10 ;
			data[87178] <= 8'h10 ;
			data[87179] <= 8'h10 ;
			data[87180] <= 8'h10 ;
			data[87181] <= 8'h10 ;
			data[87182] <= 8'h10 ;
			data[87183] <= 8'h10 ;
			data[87184] <= 8'h10 ;
			data[87185] <= 8'h10 ;
			data[87186] <= 8'h10 ;
			data[87187] <= 8'h10 ;
			data[87188] <= 8'h10 ;
			data[87189] <= 8'h10 ;
			data[87190] <= 8'h10 ;
			data[87191] <= 8'h10 ;
			data[87192] <= 8'h10 ;
			data[87193] <= 8'h10 ;
			data[87194] <= 8'h10 ;
			data[87195] <= 8'h10 ;
			data[87196] <= 8'h10 ;
			data[87197] <= 8'h10 ;
			data[87198] <= 8'h10 ;
			data[87199] <= 8'h10 ;
			data[87200] <= 8'h10 ;
			data[87201] <= 8'h10 ;
			data[87202] <= 8'h10 ;
			data[87203] <= 8'h10 ;
			data[87204] <= 8'h10 ;
			data[87205] <= 8'h10 ;
			data[87206] <= 8'h10 ;
			data[87207] <= 8'h10 ;
			data[87208] <= 8'h10 ;
			data[87209] <= 8'h10 ;
			data[87210] <= 8'h10 ;
			data[87211] <= 8'h10 ;
			data[87212] <= 8'h10 ;
			data[87213] <= 8'h10 ;
			data[87214] <= 8'h10 ;
			data[87215] <= 8'h10 ;
			data[87216] <= 8'h10 ;
			data[87217] <= 8'h10 ;
			data[87218] <= 8'h10 ;
			data[87219] <= 8'h10 ;
			data[87220] <= 8'h10 ;
			data[87221] <= 8'h10 ;
			data[87222] <= 8'h10 ;
			data[87223] <= 8'h10 ;
			data[87224] <= 8'h10 ;
			data[87225] <= 8'h10 ;
			data[87226] <= 8'h10 ;
			data[87227] <= 8'h10 ;
			data[87228] <= 8'h10 ;
			data[87229] <= 8'h10 ;
			data[87230] <= 8'h10 ;
			data[87231] <= 8'h10 ;
			data[87232] <= 8'h10 ;
			data[87233] <= 8'h10 ;
			data[87234] <= 8'h10 ;
			data[87235] <= 8'h10 ;
			data[87236] <= 8'h10 ;
			data[87237] <= 8'h10 ;
			data[87238] <= 8'h10 ;
			data[87239] <= 8'h10 ;
			data[87240] <= 8'h10 ;
			data[87241] <= 8'h10 ;
			data[87242] <= 8'h10 ;
			data[87243] <= 8'h10 ;
			data[87244] <= 8'h10 ;
			data[87245] <= 8'h10 ;
			data[87246] <= 8'h10 ;
			data[87247] <= 8'h10 ;
			data[87248] <= 8'h10 ;
			data[87249] <= 8'h10 ;
			data[87250] <= 8'h10 ;
			data[87251] <= 8'h10 ;
			data[87252] <= 8'h10 ;
			data[87253] <= 8'h10 ;
			data[87254] <= 8'h10 ;
			data[87255] <= 8'h10 ;
			data[87256] <= 8'h10 ;
			data[87257] <= 8'h10 ;
			data[87258] <= 8'h10 ;
			data[87259] <= 8'h10 ;
			data[87260] <= 8'h10 ;
			data[87261] <= 8'h10 ;
			data[87262] <= 8'h10 ;
			data[87263] <= 8'h10 ;
			data[87264] <= 8'h10 ;
			data[87265] <= 8'h10 ;
			data[87266] <= 8'h10 ;
			data[87267] <= 8'h10 ;
			data[87268] <= 8'h10 ;
			data[87269] <= 8'h10 ;
			data[87270] <= 8'h10 ;
			data[87271] <= 8'h10 ;
			data[87272] <= 8'h10 ;
			data[87273] <= 8'h10 ;
			data[87274] <= 8'h10 ;
			data[87275] <= 8'h10 ;
			data[87276] <= 8'h10 ;
			data[87277] <= 8'h10 ;
			data[87278] <= 8'h10 ;
			data[87279] <= 8'h10 ;
			data[87280] <= 8'h10 ;
			data[87281] <= 8'h10 ;
			data[87282] <= 8'h10 ;
			data[87283] <= 8'h10 ;
			data[87284] <= 8'h10 ;
			data[87285] <= 8'h10 ;
			data[87286] <= 8'h10 ;
			data[87287] <= 8'h10 ;
			data[87288] <= 8'h10 ;
			data[87289] <= 8'h10 ;
			data[87290] <= 8'h10 ;
			data[87291] <= 8'h10 ;
			data[87292] <= 8'h10 ;
			data[87293] <= 8'h10 ;
			data[87294] <= 8'h10 ;
			data[87295] <= 8'h10 ;
			data[87296] <= 8'h10 ;
			data[87297] <= 8'h10 ;
			data[87298] <= 8'h10 ;
			data[87299] <= 8'h10 ;
			data[87300] <= 8'h10 ;
			data[87301] <= 8'h10 ;
			data[87302] <= 8'h10 ;
			data[87303] <= 8'h10 ;
			data[87304] <= 8'h10 ;
			data[87305] <= 8'h10 ;
			data[87306] <= 8'h10 ;
			data[87307] <= 8'h10 ;
			data[87308] <= 8'h10 ;
			data[87309] <= 8'h10 ;
			data[87310] <= 8'h10 ;
			data[87311] <= 8'h10 ;
			data[87312] <= 8'h10 ;
			data[87313] <= 8'h10 ;
			data[87314] <= 8'h10 ;
			data[87315] <= 8'h10 ;
			data[87316] <= 8'h10 ;
			data[87317] <= 8'h10 ;
			data[87318] <= 8'h10 ;
			data[87319] <= 8'h10 ;
			data[87320] <= 8'h10 ;
			data[87321] <= 8'h10 ;
			data[87322] <= 8'h10 ;
			data[87323] <= 8'h10 ;
			data[87324] <= 8'h10 ;
			data[87325] <= 8'h10 ;
			data[87326] <= 8'h10 ;
			data[87327] <= 8'h10 ;
			data[87328] <= 8'h10 ;
			data[87329] <= 8'h10 ;
			data[87330] <= 8'h10 ;
			data[87331] <= 8'h10 ;
			data[87332] <= 8'h10 ;
			data[87333] <= 8'h10 ;
			data[87334] <= 8'h10 ;
			data[87335] <= 8'h10 ;
			data[87336] <= 8'h10 ;
			data[87337] <= 8'h10 ;
			data[87338] <= 8'h10 ;
			data[87339] <= 8'h10 ;
			data[87340] <= 8'h10 ;
			data[87341] <= 8'h10 ;
			data[87342] <= 8'h10 ;
			data[87343] <= 8'h10 ;
			data[87344] <= 8'h10 ;
			data[87345] <= 8'h10 ;
			data[87346] <= 8'h10 ;
			data[87347] <= 8'h10 ;
			data[87348] <= 8'h10 ;
			data[87349] <= 8'h10 ;
			data[87350] <= 8'h10 ;
			data[87351] <= 8'h10 ;
			data[87352] <= 8'h10 ;
			data[87353] <= 8'h10 ;
			data[87354] <= 8'h10 ;
			data[87355] <= 8'h10 ;
			data[87356] <= 8'h10 ;
			data[87357] <= 8'h10 ;
			data[87358] <= 8'h10 ;
			data[87359] <= 8'h10 ;
			data[87360] <= 8'h10 ;
			data[87361] <= 8'h10 ;
			data[87362] <= 8'h10 ;
			data[87363] <= 8'h10 ;
			data[87364] <= 8'h10 ;
			data[87365] <= 8'h10 ;
			data[87366] <= 8'h10 ;
			data[87367] <= 8'h10 ;
			data[87368] <= 8'h10 ;
			data[87369] <= 8'h10 ;
			data[87370] <= 8'h10 ;
			data[87371] <= 8'h10 ;
			data[87372] <= 8'h10 ;
			data[87373] <= 8'h10 ;
			data[87374] <= 8'h10 ;
			data[87375] <= 8'h10 ;
			data[87376] <= 8'h10 ;
			data[87377] <= 8'h10 ;
			data[87378] <= 8'h10 ;
			data[87379] <= 8'h10 ;
			data[87380] <= 8'h10 ;
			data[87381] <= 8'h10 ;
			data[87382] <= 8'h10 ;
			data[87383] <= 8'h10 ;
			data[87384] <= 8'h10 ;
			data[87385] <= 8'h10 ;
			data[87386] <= 8'h10 ;
			data[87387] <= 8'h10 ;
			data[87388] <= 8'h10 ;
			data[87389] <= 8'h10 ;
			data[87390] <= 8'h10 ;
			data[87391] <= 8'h10 ;
			data[87392] <= 8'h10 ;
			data[87393] <= 8'h10 ;
			data[87394] <= 8'h10 ;
			data[87395] <= 8'h10 ;
			data[87396] <= 8'h10 ;
			data[87397] <= 8'h10 ;
			data[87398] <= 8'h10 ;
			data[87399] <= 8'h10 ;
			data[87400] <= 8'h10 ;
			data[87401] <= 8'h10 ;
			data[87402] <= 8'h10 ;
			data[87403] <= 8'h10 ;
			data[87404] <= 8'h10 ;
			data[87405] <= 8'h10 ;
			data[87406] <= 8'h10 ;
			data[87407] <= 8'h10 ;
			data[87408] <= 8'h10 ;
			data[87409] <= 8'h10 ;
			data[87410] <= 8'h10 ;
			data[87411] <= 8'h10 ;
			data[87412] <= 8'h10 ;
			data[87413] <= 8'h10 ;
			data[87414] <= 8'h10 ;
			data[87415] <= 8'h10 ;
			data[87416] <= 8'h10 ;
			data[87417] <= 8'h10 ;
			data[87418] <= 8'h10 ;
			data[87419] <= 8'h10 ;
			data[87420] <= 8'h10 ;
			data[87421] <= 8'h10 ;
			data[87422] <= 8'h10 ;
			data[87423] <= 8'h10 ;
			data[87424] <= 8'h10 ;
			data[87425] <= 8'h10 ;
			data[87426] <= 8'h10 ;
			data[87427] <= 8'h10 ;
			data[87428] <= 8'h10 ;
			data[87429] <= 8'h10 ;
			data[87430] <= 8'h10 ;
			data[87431] <= 8'h10 ;
			data[87432] <= 8'h10 ;
			data[87433] <= 8'h10 ;
			data[87434] <= 8'h10 ;
			data[87435] <= 8'h10 ;
			data[87436] <= 8'h10 ;
			data[87437] <= 8'h10 ;
			data[87438] <= 8'h10 ;
			data[87439] <= 8'h10 ;
			data[87440] <= 8'h10 ;
			data[87441] <= 8'h10 ;
			data[87442] <= 8'h10 ;
			data[87443] <= 8'h10 ;
			data[87444] <= 8'h10 ;
			data[87445] <= 8'h10 ;
			data[87446] <= 8'h10 ;
			data[87447] <= 8'h10 ;
			data[87448] <= 8'h10 ;
			data[87449] <= 8'h10 ;
			data[87450] <= 8'h10 ;
			data[87451] <= 8'h10 ;
			data[87452] <= 8'h10 ;
			data[87453] <= 8'h10 ;
			data[87454] <= 8'h10 ;
			data[87455] <= 8'h10 ;
			data[87456] <= 8'h10 ;
			data[87457] <= 8'h10 ;
			data[87458] <= 8'h10 ;
			data[87459] <= 8'h10 ;
			data[87460] <= 8'h10 ;
			data[87461] <= 8'h10 ;
			data[87462] <= 8'h10 ;
			data[87463] <= 8'h10 ;
			data[87464] <= 8'h10 ;
			data[87465] <= 8'h10 ;
			data[87466] <= 8'h10 ;
			data[87467] <= 8'h10 ;
			data[87468] <= 8'h10 ;
			data[87469] <= 8'h10 ;
			data[87470] <= 8'h10 ;
			data[87471] <= 8'h10 ;
			data[87472] <= 8'h10 ;
			data[87473] <= 8'h10 ;
			data[87474] <= 8'h10 ;
			data[87475] <= 8'h10 ;
			data[87476] <= 8'h10 ;
			data[87477] <= 8'h10 ;
			data[87478] <= 8'h10 ;
			data[87479] <= 8'h10 ;
			data[87480] <= 8'h10 ;
			data[87481] <= 8'h10 ;
			data[87482] <= 8'h10 ;
			data[87483] <= 8'h10 ;
			data[87484] <= 8'h10 ;
			data[87485] <= 8'h10 ;
			data[87486] <= 8'h10 ;
			data[87487] <= 8'h10 ;
			data[87488] <= 8'h10 ;
			data[87489] <= 8'h10 ;
			data[87490] <= 8'h10 ;
			data[87491] <= 8'h10 ;
			data[87492] <= 8'h10 ;
			data[87493] <= 8'h10 ;
			data[87494] <= 8'h10 ;
			data[87495] <= 8'h10 ;
			data[87496] <= 8'h10 ;
			data[87497] <= 8'h10 ;
			data[87498] <= 8'h10 ;
			data[87499] <= 8'h10 ;
			data[87500] <= 8'h10 ;
			data[87501] <= 8'h10 ;
			data[87502] <= 8'h10 ;
			data[87503] <= 8'h10 ;
			data[87504] <= 8'h10 ;
			data[87505] <= 8'h10 ;
			data[87506] <= 8'h10 ;
			data[87507] <= 8'h10 ;
			data[87508] <= 8'h10 ;
			data[87509] <= 8'h10 ;
			data[87510] <= 8'h10 ;
			data[87511] <= 8'h10 ;
			data[87512] <= 8'h10 ;
			data[87513] <= 8'h10 ;
			data[87514] <= 8'h10 ;
			data[87515] <= 8'h10 ;
			data[87516] <= 8'h10 ;
			data[87517] <= 8'h10 ;
			data[87518] <= 8'h10 ;
			data[87519] <= 8'h10 ;
			data[87520] <= 8'h10 ;
			data[87521] <= 8'h10 ;
			data[87522] <= 8'h10 ;
			data[87523] <= 8'h10 ;
			data[87524] <= 8'h10 ;
			data[87525] <= 8'h10 ;
			data[87526] <= 8'h10 ;
			data[87527] <= 8'h10 ;
			data[87528] <= 8'h10 ;
			data[87529] <= 8'h10 ;
			data[87530] <= 8'h10 ;
			data[87531] <= 8'h10 ;
			data[87532] <= 8'h10 ;
			data[87533] <= 8'h10 ;
			data[87534] <= 8'h10 ;
			data[87535] <= 8'h10 ;
			data[87536] <= 8'h10 ;
			data[87537] <= 8'h10 ;
			data[87538] <= 8'h10 ;
			data[87539] <= 8'h10 ;
			data[87540] <= 8'h10 ;
			data[87541] <= 8'h10 ;
			data[87542] <= 8'h10 ;
			data[87543] <= 8'h10 ;
			data[87544] <= 8'h10 ;
			data[87545] <= 8'h10 ;
			data[87546] <= 8'h10 ;
			data[87547] <= 8'h10 ;
			data[87548] <= 8'h10 ;
			data[87549] <= 8'h10 ;
			data[87550] <= 8'h10 ;
			data[87551] <= 8'h10 ;
			data[87552] <= 8'h10 ;
			data[87553] <= 8'h10 ;
			data[87554] <= 8'h10 ;
			data[87555] <= 8'h10 ;
			data[87556] <= 8'h10 ;
			data[87557] <= 8'h10 ;
			data[87558] <= 8'h10 ;
			data[87559] <= 8'h10 ;
			data[87560] <= 8'h10 ;
			data[87561] <= 8'h10 ;
			data[87562] <= 8'h10 ;
			data[87563] <= 8'h10 ;
			data[87564] <= 8'h10 ;
			data[87565] <= 8'h10 ;
			data[87566] <= 8'h10 ;
			data[87567] <= 8'h10 ;
			data[87568] <= 8'h10 ;
			data[87569] <= 8'h10 ;
			data[87570] <= 8'h10 ;
			data[87571] <= 8'h10 ;
			data[87572] <= 8'h10 ;
			data[87573] <= 8'h10 ;
			data[87574] <= 8'h10 ;
			data[87575] <= 8'h10 ;
			data[87576] <= 8'h10 ;
			data[87577] <= 8'h10 ;
			data[87578] <= 8'h10 ;
			data[87579] <= 8'h10 ;
			data[87580] <= 8'h10 ;
			data[87581] <= 8'h10 ;
			data[87582] <= 8'h10 ;
			data[87583] <= 8'h10 ;
			data[87584] <= 8'h10 ;
			data[87585] <= 8'h10 ;
			data[87586] <= 8'h10 ;
			data[87587] <= 8'h10 ;
			data[87588] <= 8'h10 ;
			data[87589] <= 8'h10 ;
			data[87590] <= 8'h10 ;
			data[87591] <= 8'h10 ;
			data[87592] <= 8'h10 ;
			data[87593] <= 8'h10 ;
			data[87594] <= 8'h10 ;
			data[87595] <= 8'h10 ;
			data[87596] <= 8'h10 ;
			data[87597] <= 8'h10 ;
			data[87598] <= 8'h10 ;
			data[87599] <= 8'h10 ;
			data[87600] <= 8'h10 ;
			data[87601] <= 8'h10 ;
			data[87602] <= 8'h10 ;
			data[87603] <= 8'h10 ;
			data[87604] <= 8'h10 ;
			data[87605] <= 8'h10 ;
			data[87606] <= 8'h10 ;
			data[87607] <= 8'h10 ;
			data[87608] <= 8'h10 ;
			data[87609] <= 8'h10 ;
			data[87610] <= 8'h10 ;
			data[87611] <= 8'h10 ;
			data[87612] <= 8'h10 ;
			data[87613] <= 8'h10 ;
			data[87614] <= 8'h10 ;
			data[87615] <= 8'h10 ;
			data[87616] <= 8'h10 ;
			data[87617] <= 8'h10 ;
			data[87618] <= 8'h10 ;
			data[87619] <= 8'h10 ;
			data[87620] <= 8'h10 ;
			data[87621] <= 8'h10 ;
			data[87622] <= 8'h10 ;
			data[87623] <= 8'h10 ;
			data[87624] <= 8'h10 ;
			data[87625] <= 8'h10 ;
			data[87626] <= 8'h10 ;
			data[87627] <= 8'h10 ;
			data[87628] <= 8'h10 ;
			data[87629] <= 8'h10 ;
			data[87630] <= 8'h10 ;
			data[87631] <= 8'h10 ;
			data[87632] <= 8'h10 ;
			data[87633] <= 8'h10 ;
			data[87634] <= 8'h10 ;
			data[87635] <= 8'h10 ;
			data[87636] <= 8'h10 ;
			data[87637] <= 8'h10 ;
			data[87638] <= 8'h10 ;
			data[87639] <= 8'h10 ;
			data[87640] <= 8'h10 ;
			data[87641] <= 8'h10 ;
			data[87642] <= 8'h10 ;
			data[87643] <= 8'h10 ;
			data[87644] <= 8'h10 ;
			data[87645] <= 8'h10 ;
			data[87646] <= 8'h10 ;
			data[87647] <= 8'h10 ;
			data[87648] <= 8'h10 ;
			data[87649] <= 8'h10 ;
			data[87650] <= 8'h10 ;
			data[87651] <= 8'h10 ;
			data[87652] <= 8'h10 ;
			data[87653] <= 8'h10 ;
			data[87654] <= 8'h10 ;
			data[87655] <= 8'h10 ;
			data[87656] <= 8'h10 ;
			data[87657] <= 8'h10 ;
			data[87658] <= 8'h10 ;
			data[87659] <= 8'h10 ;
			data[87660] <= 8'h10 ;
			data[87661] <= 8'h10 ;
			data[87662] <= 8'h10 ;
			data[87663] <= 8'h10 ;
			data[87664] <= 8'h10 ;
			data[87665] <= 8'h10 ;
			data[87666] <= 8'h10 ;
			data[87667] <= 8'h10 ;
			data[87668] <= 8'h10 ;
			data[87669] <= 8'h10 ;
			data[87670] <= 8'h10 ;
			data[87671] <= 8'h10 ;
			data[87672] <= 8'h10 ;
			data[87673] <= 8'h10 ;
			data[87674] <= 8'h10 ;
			data[87675] <= 8'h10 ;
			data[87676] <= 8'h10 ;
			data[87677] <= 8'h10 ;
			data[87678] <= 8'h10 ;
			data[87679] <= 8'h10 ;
			data[87680] <= 8'h10 ;
			data[87681] <= 8'h10 ;
			data[87682] <= 8'h10 ;
			data[87683] <= 8'h10 ;
			data[87684] <= 8'h10 ;
			data[87685] <= 8'h10 ;
			data[87686] <= 8'h10 ;
			data[87687] <= 8'h10 ;
			data[87688] <= 8'h10 ;
			data[87689] <= 8'h10 ;
			data[87690] <= 8'h10 ;
			data[87691] <= 8'h10 ;
			data[87692] <= 8'h10 ;
			data[87693] <= 8'h10 ;
			data[87694] <= 8'h10 ;
			data[87695] <= 8'h10 ;
			data[87696] <= 8'h10 ;
			data[87697] <= 8'h10 ;
			data[87698] <= 8'h10 ;
			data[87699] <= 8'h10 ;
			data[87700] <= 8'h10 ;
			data[87701] <= 8'h10 ;
			data[87702] <= 8'h10 ;
			data[87703] <= 8'h10 ;
			data[87704] <= 8'h10 ;
			data[87705] <= 8'h10 ;
			data[87706] <= 8'h10 ;
			data[87707] <= 8'h10 ;
			data[87708] <= 8'h10 ;
			data[87709] <= 8'h10 ;
			data[87710] <= 8'h10 ;
			data[87711] <= 8'h10 ;
			data[87712] <= 8'h10 ;
			data[87713] <= 8'h10 ;
			data[87714] <= 8'h10 ;
			data[87715] <= 8'h10 ;
			data[87716] <= 8'h10 ;
			data[87717] <= 8'h10 ;
			data[87718] <= 8'h10 ;
			data[87719] <= 8'h10 ;
			data[87720] <= 8'h10 ;
			data[87721] <= 8'h10 ;
			data[87722] <= 8'h10 ;
			data[87723] <= 8'h10 ;
			data[87724] <= 8'h10 ;
			data[87725] <= 8'h10 ;
			data[87726] <= 8'h10 ;
			data[87727] <= 8'h10 ;
			data[87728] <= 8'h10 ;
			data[87729] <= 8'h10 ;
			data[87730] <= 8'h10 ;
			data[87731] <= 8'h10 ;
			data[87732] <= 8'h10 ;
			data[87733] <= 8'h10 ;
			data[87734] <= 8'h10 ;
			data[87735] <= 8'h10 ;
			data[87736] <= 8'h10 ;
			data[87737] <= 8'h10 ;
			data[87738] <= 8'h10 ;
			data[87739] <= 8'h10 ;
			data[87740] <= 8'h10 ;
			data[87741] <= 8'h10 ;
			data[87742] <= 8'h10 ;
			data[87743] <= 8'h10 ;
			data[87744] <= 8'h10 ;
			data[87745] <= 8'h10 ;
			data[87746] <= 8'h10 ;
			data[87747] <= 8'h10 ;
			data[87748] <= 8'h10 ;
			data[87749] <= 8'h10 ;
			data[87750] <= 8'h10 ;
			data[87751] <= 8'h10 ;
			data[87752] <= 8'h10 ;
			data[87753] <= 8'h10 ;
			data[87754] <= 8'h10 ;
			data[87755] <= 8'h10 ;
			data[87756] <= 8'h10 ;
			data[87757] <= 8'h10 ;
			data[87758] <= 8'h10 ;
			data[87759] <= 8'h10 ;
			data[87760] <= 8'h10 ;
			data[87761] <= 8'h10 ;
			data[87762] <= 8'h10 ;
			data[87763] <= 8'h10 ;
			data[87764] <= 8'h10 ;
			data[87765] <= 8'h10 ;
			data[87766] <= 8'h10 ;
			data[87767] <= 8'h10 ;
			data[87768] <= 8'h10 ;
			data[87769] <= 8'h10 ;
			data[87770] <= 8'h10 ;
			data[87771] <= 8'h10 ;
			data[87772] <= 8'h10 ;
			data[87773] <= 8'h10 ;
			data[87774] <= 8'h10 ;
			data[87775] <= 8'h10 ;
			data[87776] <= 8'h10 ;
			data[87777] <= 8'h10 ;
			data[87778] <= 8'h10 ;
			data[87779] <= 8'h10 ;
			data[87780] <= 8'h10 ;
			data[87781] <= 8'h10 ;
			data[87782] <= 8'h10 ;
			data[87783] <= 8'h10 ;
			data[87784] <= 8'h10 ;
			data[87785] <= 8'h10 ;
			data[87786] <= 8'h10 ;
			data[87787] <= 8'h10 ;
			data[87788] <= 8'h10 ;
			data[87789] <= 8'h10 ;
			data[87790] <= 8'h10 ;
			data[87791] <= 8'h10 ;
			data[87792] <= 8'h10 ;
			data[87793] <= 8'h10 ;
			data[87794] <= 8'h10 ;
			data[87795] <= 8'h10 ;
			data[87796] <= 8'h10 ;
			data[87797] <= 8'h10 ;
			data[87798] <= 8'h10 ;
			data[87799] <= 8'h10 ;
			data[87800] <= 8'h10 ;
			data[87801] <= 8'h10 ;
			data[87802] <= 8'h10 ;
			data[87803] <= 8'h10 ;
			data[87804] <= 8'h10 ;
			data[87805] <= 8'h10 ;
			data[87806] <= 8'h10 ;
			data[87807] <= 8'h10 ;
			data[87808] <= 8'h10 ;
			data[87809] <= 8'h10 ;
			data[87810] <= 8'h10 ;
			data[87811] <= 8'h10 ;
			data[87812] <= 8'h10 ;
			data[87813] <= 8'h10 ;
			data[87814] <= 8'h10 ;
			data[87815] <= 8'h10 ;
			data[87816] <= 8'h10 ;
			data[87817] <= 8'h10 ;
			data[87818] <= 8'h10 ;
			data[87819] <= 8'h10 ;
			data[87820] <= 8'h10 ;
			data[87821] <= 8'h10 ;
			data[87822] <= 8'h10 ;
			data[87823] <= 8'h10 ;
			data[87824] <= 8'h10 ;
			data[87825] <= 8'h10 ;
			data[87826] <= 8'h10 ;
			data[87827] <= 8'h10 ;
			data[87828] <= 8'h10 ;
			data[87829] <= 8'h10 ;
			data[87830] <= 8'h10 ;
			data[87831] <= 8'h10 ;
			data[87832] <= 8'h10 ;
			data[87833] <= 8'h10 ;
			data[87834] <= 8'h10 ;
			data[87835] <= 8'h10 ;
			data[87836] <= 8'h10 ;
			data[87837] <= 8'h10 ;
			data[87838] <= 8'h10 ;
			data[87839] <= 8'h10 ;
			data[87840] <= 8'h10 ;
			data[87841] <= 8'h10 ;
			data[87842] <= 8'h10 ;
			data[87843] <= 8'h10 ;
			data[87844] <= 8'h10 ;
			data[87845] <= 8'h10 ;
			data[87846] <= 8'h10 ;
			data[87847] <= 8'h10 ;
			data[87848] <= 8'h10 ;
			data[87849] <= 8'h10 ;
			data[87850] <= 8'h10 ;
			data[87851] <= 8'h10 ;
			data[87852] <= 8'h10 ;
			data[87853] <= 8'h10 ;
			data[87854] <= 8'h10 ;
			data[87855] <= 8'h10 ;
			data[87856] <= 8'h10 ;
			data[87857] <= 8'h10 ;
			data[87858] <= 8'h10 ;
			data[87859] <= 8'h10 ;
			data[87860] <= 8'h10 ;
			data[87861] <= 8'h10 ;
			data[87862] <= 8'h10 ;
			data[87863] <= 8'h10 ;
			data[87864] <= 8'h10 ;
			data[87865] <= 8'h10 ;
			data[87866] <= 8'h10 ;
			data[87867] <= 8'h10 ;
			data[87868] <= 8'h10 ;
			data[87869] <= 8'h10 ;
			data[87870] <= 8'h10 ;
			data[87871] <= 8'h10 ;
			data[87872] <= 8'h10 ;
			data[87873] <= 8'h10 ;
			data[87874] <= 8'h10 ;
			data[87875] <= 8'h10 ;
			data[87876] <= 8'h10 ;
			data[87877] <= 8'h10 ;
			data[87878] <= 8'h10 ;
			data[87879] <= 8'h10 ;
			data[87880] <= 8'h10 ;
			data[87881] <= 8'h10 ;
			data[87882] <= 8'h10 ;
			data[87883] <= 8'h10 ;
			data[87884] <= 8'h10 ;
			data[87885] <= 8'h10 ;
			data[87886] <= 8'h10 ;
			data[87887] <= 8'h10 ;
			data[87888] <= 8'h10 ;
			data[87889] <= 8'h10 ;
			data[87890] <= 8'h10 ;
			data[87891] <= 8'h10 ;
			data[87892] <= 8'h10 ;
			data[87893] <= 8'h10 ;
			data[87894] <= 8'h10 ;
			data[87895] <= 8'h10 ;
			data[87896] <= 8'h10 ;
			data[87897] <= 8'h10 ;
			data[87898] <= 8'h10 ;
			data[87899] <= 8'h10 ;
			data[87900] <= 8'h10 ;
			data[87901] <= 8'h10 ;
			data[87902] <= 8'h10 ;
			data[87903] <= 8'h10 ;
			data[87904] <= 8'h10 ;
			data[87905] <= 8'h10 ;
			data[87906] <= 8'h10 ;
			data[87907] <= 8'h10 ;
			data[87908] <= 8'h10 ;
			data[87909] <= 8'h10 ;
			data[87910] <= 8'h10 ;
			data[87911] <= 8'h10 ;
			data[87912] <= 8'h10 ;
			data[87913] <= 8'h10 ;
			data[87914] <= 8'h10 ;
			data[87915] <= 8'h10 ;
			data[87916] <= 8'h10 ;
			data[87917] <= 8'h10 ;
			data[87918] <= 8'h10 ;
			data[87919] <= 8'h10 ;
			data[87920] <= 8'h10 ;
			data[87921] <= 8'h10 ;
			data[87922] <= 8'h10 ;
			data[87923] <= 8'h10 ;
			data[87924] <= 8'h10 ;
			data[87925] <= 8'h10 ;
			data[87926] <= 8'h10 ;
			data[87927] <= 8'h10 ;
			data[87928] <= 8'h10 ;
			data[87929] <= 8'h10 ;
			data[87930] <= 8'h10 ;
			data[87931] <= 8'h10 ;
			data[87932] <= 8'h10 ;
			data[87933] <= 8'h10 ;
			data[87934] <= 8'h10 ;
			data[87935] <= 8'h10 ;
			data[87936] <= 8'h10 ;
			data[87937] <= 8'h10 ;
			data[87938] <= 8'h10 ;
			data[87939] <= 8'h10 ;
			data[87940] <= 8'h10 ;
			data[87941] <= 8'h10 ;
			data[87942] <= 8'h10 ;
			data[87943] <= 8'h10 ;
			data[87944] <= 8'h10 ;
			data[87945] <= 8'h10 ;
			data[87946] <= 8'h10 ;
			data[87947] <= 8'h10 ;
			data[87948] <= 8'h10 ;
			data[87949] <= 8'h10 ;
			data[87950] <= 8'h10 ;
			data[87951] <= 8'h10 ;
			data[87952] <= 8'h10 ;
			data[87953] <= 8'h10 ;
			data[87954] <= 8'h10 ;
			data[87955] <= 8'h10 ;
			data[87956] <= 8'h10 ;
			data[87957] <= 8'h10 ;
			data[87958] <= 8'h10 ;
			data[87959] <= 8'h10 ;
			data[87960] <= 8'h10 ;
			data[87961] <= 8'h10 ;
			data[87962] <= 8'h10 ;
			data[87963] <= 8'h10 ;
			data[87964] <= 8'h10 ;
			data[87965] <= 8'h10 ;
			data[87966] <= 8'h10 ;
			data[87967] <= 8'h10 ;
			data[87968] <= 8'h10 ;
			data[87969] <= 8'h10 ;
			data[87970] <= 8'h10 ;
			data[87971] <= 8'h10 ;
			data[87972] <= 8'h10 ;
			data[87973] <= 8'h10 ;
			data[87974] <= 8'h10 ;
			data[87975] <= 8'h10 ;
			data[87976] <= 8'h10 ;
			data[87977] <= 8'h10 ;
			data[87978] <= 8'h10 ;
			data[87979] <= 8'h10 ;
			data[87980] <= 8'h10 ;
			data[87981] <= 8'h10 ;
			data[87982] <= 8'h10 ;
			data[87983] <= 8'h10 ;
			data[87984] <= 8'h10 ;
			data[87985] <= 8'h10 ;
			data[87986] <= 8'h10 ;
			data[87987] <= 8'h10 ;
			data[87988] <= 8'h10 ;
			data[87989] <= 8'h10 ;
			data[87990] <= 8'h10 ;
			data[87991] <= 8'h10 ;
			data[87992] <= 8'h10 ;
			data[87993] <= 8'h10 ;
			data[87994] <= 8'h10 ;
			data[87995] <= 8'h10 ;
			data[87996] <= 8'h10 ;
			data[87997] <= 8'h10 ;
			data[87998] <= 8'h10 ;
			data[87999] <= 8'h10 ;
			data[88000] <= 8'h10 ;
			data[88001] <= 8'h10 ;
			data[88002] <= 8'h10 ;
			data[88003] <= 8'h10 ;
			data[88004] <= 8'h10 ;
			data[88005] <= 8'h10 ;
			data[88006] <= 8'h10 ;
			data[88007] <= 8'h10 ;
			data[88008] <= 8'h10 ;
			data[88009] <= 8'h10 ;
			data[88010] <= 8'h10 ;
			data[88011] <= 8'h10 ;
			data[88012] <= 8'h10 ;
			data[88013] <= 8'h10 ;
			data[88014] <= 8'h10 ;
			data[88015] <= 8'h10 ;
			data[88016] <= 8'h10 ;
			data[88017] <= 8'h10 ;
			data[88018] <= 8'h10 ;
			data[88019] <= 8'h10 ;
			data[88020] <= 8'h10 ;
			data[88021] <= 8'h10 ;
			data[88022] <= 8'h10 ;
			data[88023] <= 8'h10 ;
			data[88024] <= 8'h10 ;
			data[88025] <= 8'h10 ;
			data[88026] <= 8'h10 ;
			data[88027] <= 8'h10 ;
			data[88028] <= 8'h10 ;
			data[88029] <= 8'h10 ;
			data[88030] <= 8'h10 ;
			data[88031] <= 8'h10 ;
			data[88032] <= 8'h10 ;
			data[88033] <= 8'h10 ;
			data[88034] <= 8'h10 ;
			data[88035] <= 8'h10 ;
			data[88036] <= 8'h10 ;
			data[88037] <= 8'h10 ;
			data[88038] <= 8'h10 ;
			data[88039] <= 8'h10 ;
			data[88040] <= 8'h10 ;
			data[88041] <= 8'h10 ;
			data[88042] <= 8'h10 ;
			data[88043] <= 8'h10 ;
			data[88044] <= 8'h10 ;
			data[88045] <= 8'h10 ;
			data[88046] <= 8'h10 ;
			data[88047] <= 8'h10 ;
			data[88048] <= 8'h10 ;
			data[88049] <= 8'h10 ;
			data[88050] <= 8'h10 ;
			data[88051] <= 8'h10 ;
			data[88052] <= 8'h10 ;
			data[88053] <= 8'h10 ;
			data[88054] <= 8'h10 ;
			data[88055] <= 8'h10 ;
			data[88056] <= 8'h10 ;
			data[88057] <= 8'h10 ;
			data[88058] <= 8'h10 ;
			data[88059] <= 8'h10 ;
			data[88060] <= 8'h10 ;
			data[88061] <= 8'h10 ;
			data[88062] <= 8'h10 ;
			data[88063] <= 8'h10 ;
			data[88064] <= 8'h10 ;
			data[88065] <= 8'h10 ;
			data[88066] <= 8'h10 ;
			data[88067] <= 8'h10 ;
			data[88068] <= 8'h10 ;
			data[88069] <= 8'h10 ;
			data[88070] <= 8'h10 ;
			data[88071] <= 8'h10 ;
			data[88072] <= 8'h10 ;
			data[88073] <= 8'h10 ;
			data[88074] <= 8'h10 ;
			data[88075] <= 8'h10 ;
			data[88076] <= 8'h10 ;
			data[88077] <= 8'h10 ;
			data[88078] <= 8'h10 ;
			data[88079] <= 8'h10 ;
			data[88080] <= 8'h10 ;
			data[88081] <= 8'h10 ;
			data[88082] <= 8'h10 ;
			data[88083] <= 8'h10 ;
			data[88084] <= 8'h10 ;
			data[88085] <= 8'h10 ;
			data[88086] <= 8'h10 ;
			data[88087] <= 8'h10 ;
			data[88088] <= 8'h10 ;
			data[88089] <= 8'h10 ;
			data[88090] <= 8'h10 ;
			data[88091] <= 8'h10 ;
			data[88092] <= 8'h10 ;
			data[88093] <= 8'h10 ;
			data[88094] <= 8'h10 ;
			data[88095] <= 8'h10 ;
			data[88096] <= 8'h10 ;
			data[88097] <= 8'h10 ;
			data[88098] <= 8'h10 ;
			data[88099] <= 8'h10 ;
			data[88100] <= 8'h10 ;
			data[88101] <= 8'h10 ;
			data[88102] <= 8'h10 ;
			data[88103] <= 8'h10 ;
			data[88104] <= 8'h10 ;
			data[88105] <= 8'h10 ;
			data[88106] <= 8'h10 ;
			data[88107] <= 8'h10 ;
			data[88108] <= 8'h10 ;
			data[88109] <= 8'h10 ;
			data[88110] <= 8'h10 ;
			data[88111] <= 8'h10 ;
			data[88112] <= 8'h10 ;
			data[88113] <= 8'h10 ;
			data[88114] <= 8'h10 ;
			data[88115] <= 8'h10 ;
			data[88116] <= 8'h10 ;
			data[88117] <= 8'h10 ;
			data[88118] <= 8'h10 ;
			data[88119] <= 8'h10 ;
			data[88120] <= 8'h10 ;
			data[88121] <= 8'h10 ;
			data[88122] <= 8'h10 ;
			data[88123] <= 8'h10 ;
			data[88124] <= 8'h10 ;
			data[88125] <= 8'h10 ;
			data[88126] <= 8'h10 ;
			data[88127] <= 8'h10 ;
			data[88128] <= 8'h10 ;
			data[88129] <= 8'h10 ;
			data[88130] <= 8'h10 ;
			data[88131] <= 8'h10 ;
			data[88132] <= 8'h10 ;
			data[88133] <= 8'h10 ;
			data[88134] <= 8'h10 ;
			data[88135] <= 8'h10 ;
			data[88136] <= 8'h10 ;
			data[88137] <= 8'h10 ;
			data[88138] <= 8'h10 ;
			data[88139] <= 8'h10 ;
			data[88140] <= 8'h10 ;
			data[88141] <= 8'h10 ;
			data[88142] <= 8'h10 ;
			data[88143] <= 8'h10 ;
			data[88144] <= 8'h10 ;
			data[88145] <= 8'h10 ;
			data[88146] <= 8'h10 ;
			data[88147] <= 8'h10 ;
			data[88148] <= 8'h10 ;
			data[88149] <= 8'h10 ;
			data[88150] <= 8'h10 ;
			data[88151] <= 8'h10 ;
			data[88152] <= 8'h10 ;
			data[88153] <= 8'h10 ;
			data[88154] <= 8'h10 ;
			data[88155] <= 8'h10 ;
			data[88156] <= 8'h10 ;
			data[88157] <= 8'h10 ;
			data[88158] <= 8'h10 ;
			data[88159] <= 8'h10 ;
			data[88160] <= 8'h10 ;
			data[88161] <= 8'h10 ;
			data[88162] <= 8'h10 ;
			data[88163] <= 8'h10 ;
			data[88164] <= 8'h10 ;
			data[88165] <= 8'h10 ;
			data[88166] <= 8'h10 ;
			data[88167] <= 8'h10 ;
			data[88168] <= 8'h10 ;
			data[88169] <= 8'h10 ;
			data[88170] <= 8'h10 ;
			data[88171] <= 8'h10 ;
			data[88172] <= 8'h10 ;
			data[88173] <= 8'h10 ;
			data[88174] <= 8'h10 ;
			data[88175] <= 8'h10 ;
			data[88176] <= 8'h10 ;
			data[88177] <= 8'h10 ;
			data[88178] <= 8'h10 ;
			data[88179] <= 8'h10 ;
			data[88180] <= 8'h10 ;
			data[88181] <= 8'h10 ;
			data[88182] <= 8'h10 ;
			data[88183] <= 8'h10 ;
			data[88184] <= 8'h10 ;
			data[88185] <= 8'h10 ;
			data[88186] <= 8'h10 ;
			data[88187] <= 8'h10 ;
			data[88188] <= 8'h10 ;
			data[88189] <= 8'h10 ;
			data[88190] <= 8'h10 ;
			data[88191] <= 8'h10 ;
			data[88192] <= 8'h10 ;
			data[88193] <= 8'h10 ;
			data[88194] <= 8'h10 ;
			data[88195] <= 8'h10 ;
			data[88196] <= 8'h10 ;
			data[88197] <= 8'h10 ;
			data[88198] <= 8'h10 ;
			data[88199] <= 8'h10 ;
			data[88200] <= 8'h10 ;
			data[88201] <= 8'h10 ;
			data[88202] <= 8'h10 ;
			data[88203] <= 8'h10 ;
			data[88204] <= 8'h10 ;
			data[88205] <= 8'h10 ;
			data[88206] <= 8'h10 ;
			data[88207] <= 8'h10 ;
			data[88208] <= 8'h10 ;
			data[88209] <= 8'h10 ;
			data[88210] <= 8'h10 ;
			data[88211] <= 8'h10 ;
			data[88212] <= 8'h10 ;
			data[88213] <= 8'h10 ;
			data[88214] <= 8'h10 ;
			data[88215] <= 8'h10 ;
			data[88216] <= 8'h10 ;
			data[88217] <= 8'h10 ;
			data[88218] <= 8'h10 ;
			data[88219] <= 8'h10 ;
			data[88220] <= 8'h10 ;
			data[88221] <= 8'h10 ;
			data[88222] <= 8'h10 ;
			data[88223] <= 8'h10 ;
			data[88224] <= 8'h10 ;
			data[88225] <= 8'h10 ;
			data[88226] <= 8'h10 ;
			data[88227] <= 8'h10 ;
			data[88228] <= 8'h10 ;
			data[88229] <= 8'h10 ;
			data[88230] <= 8'h10 ;
			data[88231] <= 8'h10 ;
			data[88232] <= 8'h10 ;
			data[88233] <= 8'h10 ;
			data[88234] <= 8'h10 ;
			data[88235] <= 8'h10 ;
			data[88236] <= 8'h10 ;
			data[88237] <= 8'h10 ;
			data[88238] <= 8'h10 ;
			data[88239] <= 8'h10 ;
			data[88240] <= 8'h10 ;
			data[88241] <= 8'h10 ;
			data[88242] <= 8'h10 ;
			data[88243] <= 8'h10 ;
			data[88244] <= 8'h10 ;
			data[88245] <= 8'h10 ;
			data[88246] <= 8'h10 ;
			data[88247] <= 8'h10 ;
			data[88248] <= 8'h10 ;
			data[88249] <= 8'h10 ;
			data[88250] <= 8'h10 ;
			data[88251] <= 8'h10 ;
			data[88252] <= 8'h10 ;
			data[88253] <= 8'h10 ;
			data[88254] <= 8'h10 ;
			data[88255] <= 8'h10 ;
			data[88256] <= 8'h10 ;
			data[88257] <= 8'h10 ;
			data[88258] <= 8'h10 ;
			data[88259] <= 8'h10 ;
			data[88260] <= 8'h10 ;
			data[88261] <= 8'h10 ;
			data[88262] <= 8'h10 ;
			data[88263] <= 8'h10 ;
			data[88264] <= 8'h10 ;
			data[88265] <= 8'h10 ;
			data[88266] <= 8'h10 ;
			data[88267] <= 8'h10 ;
			data[88268] <= 8'h10 ;
			data[88269] <= 8'h10 ;
			data[88270] <= 8'h10 ;
			data[88271] <= 8'h10 ;
			data[88272] <= 8'h10 ;
			data[88273] <= 8'h10 ;
			data[88274] <= 8'h10 ;
			data[88275] <= 8'h10 ;
			data[88276] <= 8'h10 ;
			data[88277] <= 8'h10 ;
			data[88278] <= 8'h10 ;
			data[88279] <= 8'h10 ;
			data[88280] <= 8'h10 ;
			data[88281] <= 8'h10 ;
			data[88282] <= 8'h10 ;
			data[88283] <= 8'h10 ;
			data[88284] <= 8'h10 ;
			data[88285] <= 8'h10 ;
			data[88286] <= 8'h10 ;
			data[88287] <= 8'h10 ;
			data[88288] <= 8'h10 ;
			data[88289] <= 8'h10 ;
			data[88290] <= 8'h10 ;
			data[88291] <= 8'h10 ;
			data[88292] <= 8'h10 ;
			data[88293] <= 8'h10 ;
			data[88294] <= 8'h10 ;
			data[88295] <= 8'h10 ;
			data[88296] <= 8'h10 ;
			data[88297] <= 8'h10 ;
			data[88298] <= 8'h10 ;
			data[88299] <= 8'h10 ;
			data[88300] <= 8'h10 ;
			data[88301] <= 8'h10 ;
			data[88302] <= 8'h10 ;
			data[88303] <= 8'h10 ;
			data[88304] <= 8'h10 ;
			data[88305] <= 8'h10 ;
			data[88306] <= 8'h10 ;
			data[88307] <= 8'h10 ;
			data[88308] <= 8'h10 ;
			data[88309] <= 8'h10 ;
			data[88310] <= 8'h10 ;
			data[88311] <= 8'h10 ;
			data[88312] <= 8'h10 ;
			data[88313] <= 8'h10 ;
			data[88314] <= 8'h10 ;
			data[88315] <= 8'h10 ;
			data[88316] <= 8'h10 ;
			data[88317] <= 8'h10 ;
			data[88318] <= 8'h10 ;
			data[88319] <= 8'h10 ;
			data[88320] <= 8'h10 ;
			data[88321] <= 8'h10 ;
			data[88322] <= 8'h10 ;
			data[88323] <= 8'h10 ;
			data[88324] <= 8'h10 ;
			data[88325] <= 8'h10 ;
			data[88326] <= 8'h10 ;
			data[88327] <= 8'h10 ;
			data[88328] <= 8'h10 ;
			data[88329] <= 8'h10 ;
			data[88330] <= 8'h10 ;
			data[88331] <= 8'h10 ;
			data[88332] <= 8'h10 ;
			data[88333] <= 8'h10 ;
			data[88334] <= 8'h10 ;
			data[88335] <= 8'h10 ;
			data[88336] <= 8'h10 ;
			data[88337] <= 8'h10 ;
			data[88338] <= 8'h10 ;
			data[88339] <= 8'h10 ;
			data[88340] <= 8'h10 ;
			data[88341] <= 8'h10 ;
			data[88342] <= 8'h10 ;
			data[88343] <= 8'h10 ;
			data[88344] <= 8'h10 ;
			data[88345] <= 8'h10 ;
			data[88346] <= 8'h10 ;
			data[88347] <= 8'h10 ;
			data[88348] <= 8'h10 ;
			data[88349] <= 8'h10 ;
			data[88350] <= 8'h10 ;
			data[88351] <= 8'h10 ;
			data[88352] <= 8'h10 ;
			data[88353] <= 8'h10 ;
			data[88354] <= 8'h10 ;
			data[88355] <= 8'h10 ;
			data[88356] <= 8'h10 ;
			data[88357] <= 8'h10 ;
			data[88358] <= 8'h10 ;
			data[88359] <= 8'h10 ;
			data[88360] <= 8'h10 ;
			data[88361] <= 8'h10 ;
			data[88362] <= 8'h10 ;
			data[88363] <= 8'h10 ;
			data[88364] <= 8'h10 ;
			data[88365] <= 8'h10 ;
			data[88366] <= 8'h10 ;
			data[88367] <= 8'h10 ;
			data[88368] <= 8'h10 ;
			data[88369] <= 8'h10 ;
			data[88370] <= 8'h10 ;
			data[88371] <= 8'h10 ;
			data[88372] <= 8'h10 ;
			data[88373] <= 8'h10 ;
			data[88374] <= 8'h10 ;
			data[88375] <= 8'h10 ;
			data[88376] <= 8'h10 ;
			data[88377] <= 8'h10 ;
			data[88378] <= 8'h10 ;
			data[88379] <= 8'h10 ;
			data[88380] <= 8'h10 ;
			data[88381] <= 8'h10 ;
			data[88382] <= 8'h10 ;
			data[88383] <= 8'h10 ;
			data[88384] <= 8'h10 ;
			data[88385] <= 8'h10 ;
			data[88386] <= 8'h10 ;
			data[88387] <= 8'h10 ;
			data[88388] <= 8'h10 ;
			data[88389] <= 8'h10 ;
			data[88390] <= 8'h10 ;
			data[88391] <= 8'h10 ;
			data[88392] <= 8'h10 ;
			data[88393] <= 8'h10 ;
			data[88394] <= 8'h10 ;
			data[88395] <= 8'h10 ;
			data[88396] <= 8'h10 ;
			data[88397] <= 8'h10 ;
			data[88398] <= 8'h10 ;
			data[88399] <= 8'h10 ;
			data[88400] <= 8'h10 ;
			data[88401] <= 8'h10 ;
			data[88402] <= 8'h10 ;
			data[88403] <= 8'h10 ;
			data[88404] <= 8'h10 ;
			data[88405] <= 8'h10 ;
			data[88406] <= 8'h10 ;
			data[88407] <= 8'h10 ;
			data[88408] <= 8'h10 ;
			data[88409] <= 8'h10 ;
			data[88410] <= 8'h10 ;
			data[88411] <= 8'h10 ;
			data[88412] <= 8'h10 ;
			data[88413] <= 8'h10 ;
			data[88414] <= 8'h10 ;
			data[88415] <= 8'h10 ;
			data[88416] <= 8'h10 ;
			data[88417] <= 8'h10 ;
			data[88418] <= 8'h10 ;
			data[88419] <= 8'h10 ;
			data[88420] <= 8'h10 ;
			data[88421] <= 8'h10 ;
			data[88422] <= 8'h10 ;
			data[88423] <= 8'h10 ;
			data[88424] <= 8'h10 ;
			data[88425] <= 8'h10 ;
			data[88426] <= 8'h10 ;
			data[88427] <= 8'h10 ;
			data[88428] <= 8'h10 ;
			data[88429] <= 8'h10 ;
			data[88430] <= 8'h10 ;
			data[88431] <= 8'h10 ;
			data[88432] <= 8'h10 ;
			data[88433] <= 8'h10 ;
			data[88434] <= 8'h10 ;
			data[88435] <= 8'h10 ;
			data[88436] <= 8'h10 ;
			data[88437] <= 8'h10 ;
			data[88438] <= 8'h10 ;
			data[88439] <= 8'h10 ;
			data[88440] <= 8'h10 ;
			data[88441] <= 8'h10 ;
			data[88442] <= 8'h10 ;
			data[88443] <= 8'h10 ;
			data[88444] <= 8'h10 ;
			data[88445] <= 8'h10 ;
			data[88446] <= 8'h10 ;
			data[88447] <= 8'h10 ;
			data[88448] <= 8'h10 ;
			data[88449] <= 8'h10 ;
			data[88450] <= 8'h10 ;
			data[88451] <= 8'h10 ;
			data[88452] <= 8'h10 ;
			data[88453] <= 8'h10 ;
			data[88454] <= 8'h10 ;
			data[88455] <= 8'h10 ;
			data[88456] <= 8'h10 ;
			data[88457] <= 8'h10 ;
			data[88458] <= 8'h10 ;
			data[88459] <= 8'h10 ;
			data[88460] <= 8'h10 ;
			data[88461] <= 8'h10 ;
			data[88462] <= 8'h10 ;
			data[88463] <= 8'h10 ;
			data[88464] <= 8'h10 ;
			data[88465] <= 8'h10 ;
			data[88466] <= 8'h10 ;
			data[88467] <= 8'h10 ;
			data[88468] <= 8'h10 ;
			data[88469] <= 8'h10 ;
			data[88470] <= 8'h10 ;
			data[88471] <= 8'h10 ;
			data[88472] <= 8'h10 ;
			data[88473] <= 8'h10 ;
			data[88474] <= 8'h10 ;
			data[88475] <= 8'h10 ;
			data[88476] <= 8'h10 ;
			data[88477] <= 8'h10 ;
			data[88478] <= 8'h10 ;
			data[88479] <= 8'h10 ;
			data[88480] <= 8'h10 ;
			data[88481] <= 8'h10 ;
			data[88482] <= 8'h10 ;
			data[88483] <= 8'h10 ;
			data[88484] <= 8'h10 ;
			data[88485] <= 8'h10 ;
			data[88486] <= 8'h10 ;
			data[88487] <= 8'h10 ;
			data[88488] <= 8'h10 ;
			data[88489] <= 8'h10 ;
			data[88490] <= 8'h10 ;
			data[88491] <= 8'h10 ;
			data[88492] <= 8'h10 ;
			data[88493] <= 8'h10 ;
			data[88494] <= 8'h10 ;
			data[88495] <= 8'h10 ;
			data[88496] <= 8'h10 ;
			data[88497] <= 8'h10 ;
			data[88498] <= 8'h10 ;
			data[88499] <= 8'h10 ;
			data[88500] <= 8'h10 ;
			data[88501] <= 8'h10 ;
			data[88502] <= 8'h10 ;
			data[88503] <= 8'h10 ;
			data[88504] <= 8'h10 ;
			data[88505] <= 8'h10 ;
			data[88506] <= 8'h10 ;
			data[88507] <= 8'h10 ;
			data[88508] <= 8'h10 ;
			data[88509] <= 8'h10 ;
			data[88510] <= 8'h10 ;
			data[88511] <= 8'h10 ;
			data[88512] <= 8'h10 ;
			data[88513] <= 8'h10 ;
			data[88514] <= 8'h10 ;
			data[88515] <= 8'h10 ;
			data[88516] <= 8'h10 ;
			data[88517] <= 8'h10 ;
			data[88518] <= 8'h10 ;
			data[88519] <= 8'h10 ;
			data[88520] <= 8'h10 ;
			data[88521] <= 8'h10 ;
			data[88522] <= 8'h10 ;
			data[88523] <= 8'h10 ;
			data[88524] <= 8'h10 ;
			data[88525] <= 8'h10 ;
			data[88526] <= 8'h10 ;
			data[88527] <= 8'h10 ;
			data[88528] <= 8'h10 ;
			data[88529] <= 8'h10 ;
			data[88530] <= 8'h10 ;
			data[88531] <= 8'h10 ;
			data[88532] <= 8'h10 ;
			data[88533] <= 8'h10 ;
			data[88534] <= 8'h10 ;
			data[88535] <= 8'h10 ;
			data[88536] <= 8'h10 ;
			data[88537] <= 8'h10 ;
			data[88538] <= 8'h10 ;
			data[88539] <= 8'h10 ;
			data[88540] <= 8'h10 ;
			data[88541] <= 8'h10 ;
			data[88542] <= 8'h10 ;
			data[88543] <= 8'h10 ;
			data[88544] <= 8'h10 ;
			data[88545] <= 8'h10 ;
			data[88546] <= 8'h10 ;
			data[88547] <= 8'h10 ;
			data[88548] <= 8'h10 ;
			data[88549] <= 8'h10 ;
			data[88550] <= 8'h10 ;
			data[88551] <= 8'h10 ;
			data[88552] <= 8'h10 ;
			data[88553] <= 8'h10 ;
			data[88554] <= 8'h10 ;
			data[88555] <= 8'h10 ;
			data[88556] <= 8'h10 ;
			data[88557] <= 8'h10 ;
			data[88558] <= 8'h10 ;
			data[88559] <= 8'h10 ;
			data[88560] <= 8'h10 ;
			data[88561] <= 8'h10 ;
			data[88562] <= 8'h10 ;
			data[88563] <= 8'h10 ;
			data[88564] <= 8'h10 ;
			data[88565] <= 8'h10 ;
			data[88566] <= 8'h10 ;
			data[88567] <= 8'h10 ;
			data[88568] <= 8'h10 ;
			data[88569] <= 8'h10 ;
			data[88570] <= 8'h10 ;
			data[88571] <= 8'h10 ;
			data[88572] <= 8'h10 ;
			data[88573] <= 8'h10 ;
			data[88574] <= 8'h10 ;
			data[88575] <= 8'h10 ;
			data[88576] <= 8'h10 ;
			data[88577] <= 8'h10 ;
			data[88578] <= 8'h10 ;
			data[88579] <= 8'h10 ;
			data[88580] <= 8'h10 ;
			data[88581] <= 8'h10 ;
			data[88582] <= 8'h10 ;
			data[88583] <= 8'h10 ;
			data[88584] <= 8'h10 ;
			data[88585] <= 8'h10 ;
			data[88586] <= 8'h10 ;
			data[88587] <= 8'h10 ;
			data[88588] <= 8'h10 ;
			data[88589] <= 8'h10 ;
			data[88590] <= 8'h10 ;
			data[88591] <= 8'h10 ;
			data[88592] <= 8'h10 ;
			data[88593] <= 8'h10 ;
			data[88594] <= 8'h10 ;
			data[88595] <= 8'h10 ;
			data[88596] <= 8'h10 ;
			data[88597] <= 8'h10 ;
			data[88598] <= 8'h10 ;
			data[88599] <= 8'h10 ;
			data[88600] <= 8'h10 ;
			data[88601] <= 8'h10 ;
			data[88602] <= 8'h10 ;
			data[88603] <= 8'h10 ;
			data[88604] <= 8'h10 ;
			data[88605] <= 8'h10 ;
			data[88606] <= 8'h10 ;
			data[88607] <= 8'h10 ;
			data[88608] <= 8'h10 ;
			data[88609] <= 8'h10 ;
			data[88610] <= 8'h10 ;
			data[88611] <= 8'h10 ;
			data[88612] <= 8'h10 ;
			data[88613] <= 8'h10 ;
			data[88614] <= 8'h10 ;
			data[88615] <= 8'h10 ;
			data[88616] <= 8'h10 ;
			data[88617] <= 8'h10 ;
			data[88618] <= 8'h10 ;
			data[88619] <= 8'h10 ;
			data[88620] <= 8'h10 ;
			data[88621] <= 8'h10 ;
			data[88622] <= 8'h10 ;
			data[88623] <= 8'h10 ;
			data[88624] <= 8'h10 ;
			data[88625] <= 8'h10 ;
			data[88626] <= 8'h10 ;
			data[88627] <= 8'h10 ;
			data[88628] <= 8'h10 ;
			data[88629] <= 8'h10 ;
			data[88630] <= 8'h10 ;
			data[88631] <= 8'h10 ;
			data[88632] <= 8'h10 ;
			data[88633] <= 8'h10 ;
			data[88634] <= 8'h10 ;
			data[88635] <= 8'h10 ;
			data[88636] <= 8'h10 ;
			data[88637] <= 8'h10 ;
			data[88638] <= 8'h10 ;
			data[88639] <= 8'h10 ;
			data[88640] <= 8'h10 ;
			data[88641] <= 8'h10 ;
			data[88642] <= 8'h10 ;
			data[88643] <= 8'h10 ;
			data[88644] <= 8'h10 ;
			data[88645] <= 8'h10 ;
			data[88646] <= 8'h10 ;
			data[88647] <= 8'h10 ;
			data[88648] <= 8'h10 ;
			data[88649] <= 8'h10 ;
			data[88650] <= 8'h10 ;
			data[88651] <= 8'h10 ;
			data[88652] <= 8'h10 ;
			data[88653] <= 8'h10 ;
			data[88654] <= 8'h10 ;
			data[88655] <= 8'h10 ;
			data[88656] <= 8'h10 ;
			data[88657] <= 8'h10 ;
			data[88658] <= 8'h10 ;
			data[88659] <= 8'h10 ;
			data[88660] <= 8'h10 ;
			data[88661] <= 8'h10 ;
			data[88662] <= 8'h10 ;
			data[88663] <= 8'h10 ;
			data[88664] <= 8'h10 ;
			data[88665] <= 8'h10 ;
			data[88666] <= 8'h10 ;
			data[88667] <= 8'h10 ;
			data[88668] <= 8'h10 ;
			data[88669] <= 8'h10 ;
			data[88670] <= 8'h10 ;
			data[88671] <= 8'h10 ;
			data[88672] <= 8'h10 ;
			data[88673] <= 8'h10 ;
			data[88674] <= 8'h10 ;
			data[88675] <= 8'h10 ;
			data[88676] <= 8'h10 ;
			data[88677] <= 8'h10 ;
			data[88678] <= 8'h10 ;
			data[88679] <= 8'h10 ;
			data[88680] <= 8'h10 ;
			data[88681] <= 8'h10 ;
			data[88682] <= 8'h10 ;
			data[88683] <= 8'h10 ;
			data[88684] <= 8'h10 ;
			data[88685] <= 8'h10 ;
			data[88686] <= 8'h10 ;
			data[88687] <= 8'h10 ;
			data[88688] <= 8'h10 ;
			data[88689] <= 8'h10 ;
			data[88690] <= 8'h10 ;
			data[88691] <= 8'h10 ;
			data[88692] <= 8'h10 ;
			data[88693] <= 8'h10 ;
			data[88694] <= 8'h10 ;
			data[88695] <= 8'h10 ;
			data[88696] <= 8'h10 ;
			data[88697] <= 8'h10 ;
			data[88698] <= 8'h10 ;
			data[88699] <= 8'h10 ;
			data[88700] <= 8'h10 ;
			data[88701] <= 8'h10 ;
			data[88702] <= 8'h10 ;
			data[88703] <= 8'h10 ;
			data[88704] <= 8'h10 ;
			data[88705] <= 8'h10 ;
			data[88706] <= 8'h10 ;
			data[88707] <= 8'h10 ;
			data[88708] <= 8'h10 ;
			data[88709] <= 8'h10 ;
			data[88710] <= 8'h10 ;
			data[88711] <= 8'h10 ;
			data[88712] <= 8'h10 ;
			data[88713] <= 8'h10 ;
			data[88714] <= 8'h10 ;
			data[88715] <= 8'h10 ;
			data[88716] <= 8'h10 ;
			data[88717] <= 8'h10 ;
			data[88718] <= 8'h10 ;
			data[88719] <= 8'h10 ;
			data[88720] <= 8'h10 ;
			data[88721] <= 8'h10 ;
			data[88722] <= 8'h10 ;
			data[88723] <= 8'h10 ;
			data[88724] <= 8'h10 ;
			data[88725] <= 8'h10 ;
			data[88726] <= 8'h10 ;
			data[88727] <= 8'h10 ;
			data[88728] <= 8'h10 ;
			data[88729] <= 8'h10 ;
			data[88730] <= 8'h10 ;
			data[88731] <= 8'h10 ;
			data[88732] <= 8'h10 ;
			data[88733] <= 8'h10 ;
			data[88734] <= 8'h10 ;
			data[88735] <= 8'h10 ;
			data[88736] <= 8'h10 ;
			data[88737] <= 8'h10 ;
			data[88738] <= 8'h10 ;
			data[88739] <= 8'h10 ;
			data[88740] <= 8'h10 ;
			data[88741] <= 8'h10 ;
			data[88742] <= 8'h10 ;
			data[88743] <= 8'h10 ;
			data[88744] <= 8'h10 ;
			data[88745] <= 8'h10 ;
			data[88746] <= 8'h10 ;
			data[88747] <= 8'h10 ;
			data[88748] <= 8'h10 ;
			data[88749] <= 8'h10 ;
			data[88750] <= 8'h10 ;
			data[88751] <= 8'h10 ;
			data[88752] <= 8'h10 ;
			data[88753] <= 8'h10 ;
			data[88754] <= 8'h10 ;
			data[88755] <= 8'h10 ;
			data[88756] <= 8'h10 ;
			data[88757] <= 8'h10 ;
			data[88758] <= 8'h10 ;
			data[88759] <= 8'h10 ;
			data[88760] <= 8'h10 ;
			data[88761] <= 8'h10 ;
			data[88762] <= 8'h10 ;
			data[88763] <= 8'h10 ;
			data[88764] <= 8'h10 ;
			data[88765] <= 8'h10 ;
			data[88766] <= 8'h10 ;
			data[88767] <= 8'h10 ;
			data[88768] <= 8'h10 ;
			data[88769] <= 8'h10 ;
			data[88770] <= 8'h10 ;
			data[88771] <= 8'h10 ;
			data[88772] <= 8'h10 ;
			data[88773] <= 8'h10 ;
			data[88774] <= 8'h10 ;
			data[88775] <= 8'h10 ;
			data[88776] <= 8'h10 ;
			data[88777] <= 8'h10 ;
			data[88778] <= 8'h10 ;
			data[88779] <= 8'h10 ;
			data[88780] <= 8'h10 ;
			data[88781] <= 8'h10 ;
			data[88782] <= 8'h10 ;
			data[88783] <= 8'h10 ;
			data[88784] <= 8'h10 ;
			data[88785] <= 8'h10 ;
			data[88786] <= 8'h10 ;
			data[88787] <= 8'h10 ;
			data[88788] <= 8'h10 ;
			data[88789] <= 8'h10 ;
			data[88790] <= 8'h10 ;
			data[88791] <= 8'h10 ;
			data[88792] <= 8'h10 ;
			data[88793] <= 8'h10 ;
			data[88794] <= 8'h10 ;
			data[88795] <= 8'h10 ;
			data[88796] <= 8'h10 ;
			data[88797] <= 8'h10 ;
			data[88798] <= 8'h10 ;
			data[88799] <= 8'h10 ;
			data[88800] <= 8'h10 ;
			data[88801] <= 8'h10 ;
			data[88802] <= 8'h10 ;
			data[88803] <= 8'h10 ;
			data[88804] <= 8'h10 ;
			data[88805] <= 8'h10 ;
			data[88806] <= 8'h10 ;
			data[88807] <= 8'h10 ;
			data[88808] <= 8'h10 ;
			data[88809] <= 8'h10 ;
			data[88810] <= 8'h10 ;
			data[88811] <= 8'h10 ;
			data[88812] <= 8'h10 ;
			data[88813] <= 8'h10 ;
			data[88814] <= 8'h10 ;
			data[88815] <= 8'h10 ;
			data[88816] <= 8'h10 ;
			data[88817] <= 8'h10 ;
			data[88818] <= 8'h10 ;
			data[88819] <= 8'h10 ;
			data[88820] <= 8'h10 ;
			data[88821] <= 8'h10 ;
			data[88822] <= 8'h10 ;
			data[88823] <= 8'h10 ;
			data[88824] <= 8'h10 ;
			data[88825] <= 8'h10 ;
			data[88826] <= 8'h10 ;
			data[88827] <= 8'h10 ;
			data[88828] <= 8'h10 ;
			data[88829] <= 8'h10 ;
			data[88830] <= 8'h10 ;
			data[88831] <= 8'h10 ;
			data[88832] <= 8'h10 ;
			data[88833] <= 8'h10 ;
			data[88834] <= 8'h10 ;
			data[88835] <= 8'h10 ;
			data[88836] <= 8'h10 ;
			data[88837] <= 8'h10 ;
			data[88838] <= 8'h10 ;
			data[88839] <= 8'h10 ;
			data[88840] <= 8'h10 ;
			data[88841] <= 8'h10 ;
			data[88842] <= 8'h10 ;
			data[88843] <= 8'h10 ;
			data[88844] <= 8'h10 ;
			data[88845] <= 8'h10 ;
			data[88846] <= 8'h10 ;
			data[88847] <= 8'h10 ;
			data[88848] <= 8'h10 ;
			data[88849] <= 8'h10 ;
			data[88850] <= 8'h10 ;
			data[88851] <= 8'h10 ;
			data[88852] <= 8'h10 ;
			data[88853] <= 8'h10 ;
			data[88854] <= 8'h10 ;
			data[88855] <= 8'h10 ;
			data[88856] <= 8'h10 ;
			data[88857] <= 8'h10 ;
			data[88858] <= 8'h10 ;
			data[88859] <= 8'h10 ;
			data[88860] <= 8'h10 ;
			data[88861] <= 8'h10 ;
			data[88862] <= 8'h10 ;
			data[88863] <= 8'h10 ;
			data[88864] <= 8'h10 ;
			data[88865] <= 8'h10 ;
			data[88866] <= 8'h10 ;
			data[88867] <= 8'h10 ;
			data[88868] <= 8'h10 ;
			data[88869] <= 8'h10 ;
			data[88870] <= 8'h10 ;
			data[88871] <= 8'h10 ;
			data[88872] <= 8'h10 ;
			data[88873] <= 8'h10 ;
			data[88874] <= 8'h10 ;
			data[88875] <= 8'h10 ;
			data[88876] <= 8'h10 ;
			data[88877] <= 8'h10 ;
			data[88878] <= 8'h10 ;
			data[88879] <= 8'h10 ;
			data[88880] <= 8'h10 ;
			data[88881] <= 8'h10 ;
			data[88882] <= 8'h10 ;
			data[88883] <= 8'h10 ;
			data[88884] <= 8'h10 ;
			data[88885] <= 8'h10 ;
			data[88886] <= 8'h10 ;
			data[88887] <= 8'h10 ;
			data[88888] <= 8'h10 ;
			data[88889] <= 8'h10 ;
			data[88890] <= 8'h10 ;
			data[88891] <= 8'h10 ;
			data[88892] <= 8'h10 ;
			data[88893] <= 8'h10 ;
			data[88894] <= 8'h10 ;
			data[88895] <= 8'h10 ;
			data[88896] <= 8'h10 ;
			data[88897] <= 8'h10 ;
			data[88898] <= 8'h10 ;
			data[88899] <= 8'h10 ;
			data[88900] <= 8'h10 ;
			data[88901] <= 8'h10 ;
			data[88902] <= 8'h10 ;
			data[88903] <= 8'h10 ;
			data[88904] <= 8'h10 ;
			data[88905] <= 8'h10 ;
			data[88906] <= 8'h10 ;
			data[88907] <= 8'h10 ;
			data[88908] <= 8'h10 ;
			data[88909] <= 8'h10 ;
			data[88910] <= 8'h10 ;
			data[88911] <= 8'h10 ;
			data[88912] <= 8'h10 ;
			data[88913] <= 8'h10 ;
			data[88914] <= 8'h10 ;
			data[88915] <= 8'h10 ;
			data[88916] <= 8'h10 ;
			data[88917] <= 8'h10 ;
			data[88918] <= 8'h10 ;
			data[88919] <= 8'h10 ;
			data[88920] <= 8'h10 ;
			data[88921] <= 8'h10 ;
			data[88922] <= 8'h10 ;
			data[88923] <= 8'h10 ;
			data[88924] <= 8'h10 ;
			data[88925] <= 8'h10 ;
			data[88926] <= 8'h10 ;
			data[88927] <= 8'h10 ;
			data[88928] <= 8'h10 ;
			data[88929] <= 8'h10 ;
			data[88930] <= 8'h10 ;
			data[88931] <= 8'h10 ;
			data[88932] <= 8'h10 ;
			data[88933] <= 8'h10 ;
			data[88934] <= 8'h10 ;
			data[88935] <= 8'h10 ;
			data[88936] <= 8'h10 ;
			data[88937] <= 8'h10 ;
			data[88938] <= 8'h10 ;
			data[88939] <= 8'h10 ;
			data[88940] <= 8'h10 ;
			data[88941] <= 8'h10 ;
			data[88942] <= 8'h10 ;
			data[88943] <= 8'h10 ;
			data[88944] <= 8'h10 ;
			data[88945] <= 8'h10 ;
			data[88946] <= 8'h10 ;
			data[88947] <= 8'h10 ;
			data[88948] <= 8'h10 ;
			data[88949] <= 8'h10 ;
			data[88950] <= 8'h10 ;
			data[88951] <= 8'h10 ;
			data[88952] <= 8'h10 ;
			data[88953] <= 8'h10 ;
			data[88954] <= 8'h10 ;
			data[88955] <= 8'h10 ;
			data[88956] <= 8'h10 ;
			data[88957] <= 8'h10 ;
			data[88958] <= 8'h10 ;
			data[88959] <= 8'h10 ;
			data[88960] <= 8'h10 ;
			data[88961] <= 8'h10 ;
			data[88962] <= 8'h10 ;
			data[88963] <= 8'h10 ;
			data[88964] <= 8'h10 ;
			data[88965] <= 8'h10 ;
			data[88966] <= 8'h10 ;
			data[88967] <= 8'h10 ;
			data[88968] <= 8'h10 ;
			data[88969] <= 8'h10 ;
			data[88970] <= 8'h10 ;
			data[88971] <= 8'h10 ;
			data[88972] <= 8'h10 ;
			data[88973] <= 8'h10 ;
			data[88974] <= 8'h10 ;
			data[88975] <= 8'h10 ;
			data[88976] <= 8'h10 ;
			data[88977] <= 8'h10 ;
			data[88978] <= 8'h10 ;
			data[88979] <= 8'h10 ;
			data[88980] <= 8'h10 ;
			data[88981] <= 8'h10 ;
			data[88982] <= 8'h10 ;
			data[88983] <= 8'h10 ;
			data[88984] <= 8'h10 ;
			data[88985] <= 8'h10 ;
			data[88986] <= 8'h10 ;
			data[88987] <= 8'h10 ;
			data[88988] <= 8'h10 ;
			data[88989] <= 8'h10 ;
			data[88990] <= 8'h10 ;
			data[88991] <= 8'h10 ;
			data[88992] <= 8'h10 ;
			data[88993] <= 8'h10 ;
			data[88994] <= 8'h10 ;
			data[88995] <= 8'h10 ;
			data[88996] <= 8'h10 ;
			data[88997] <= 8'h10 ;
			data[88998] <= 8'h10 ;
			data[88999] <= 8'h10 ;
			data[89000] <= 8'h10 ;
			data[89001] <= 8'h10 ;
			data[89002] <= 8'h10 ;
			data[89003] <= 8'h10 ;
			data[89004] <= 8'h10 ;
			data[89005] <= 8'h10 ;
			data[89006] <= 8'h10 ;
			data[89007] <= 8'h10 ;
			data[89008] <= 8'h10 ;
			data[89009] <= 8'h10 ;
			data[89010] <= 8'h10 ;
			data[89011] <= 8'h10 ;
			data[89012] <= 8'h10 ;
			data[89013] <= 8'h10 ;
			data[89014] <= 8'h10 ;
			data[89015] <= 8'h10 ;
			data[89016] <= 8'h10 ;
			data[89017] <= 8'h10 ;
			data[89018] <= 8'h10 ;
			data[89019] <= 8'h10 ;
			data[89020] <= 8'h10 ;
			data[89021] <= 8'h10 ;
			data[89022] <= 8'h10 ;
			data[89023] <= 8'h10 ;
			data[89024] <= 8'h10 ;
			data[89025] <= 8'h10 ;
			data[89026] <= 8'h10 ;
			data[89027] <= 8'h10 ;
			data[89028] <= 8'h10 ;
			data[89029] <= 8'h10 ;
			data[89030] <= 8'h10 ;
			data[89031] <= 8'h10 ;
			data[89032] <= 8'h10 ;
			data[89033] <= 8'h10 ;
			data[89034] <= 8'h10 ;
			data[89035] <= 8'h10 ;
			data[89036] <= 8'h10 ;
			data[89037] <= 8'h10 ;
			data[89038] <= 8'h10 ;
			data[89039] <= 8'h10 ;
			data[89040] <= 8'h10 ;
			data[89041] <= 8'h10 ;
			data[89042] <= 8'h10 ;
			data[89043] <= 8'h10 ;
			data[89044] <= 8'h10 ;
			data[89045] <= 8'h10 ;
			data[89046] <= 8'h10 ;
			data[89047] <= 8'h10 ;
			data[89048] <= 8'h10 ;
			data[89049] <= 8'h10 ;
			data[89050] <= 8'h10 ;
			data[89051] <= 8'h10 ;
			data[89052] <= 8'h10 ;
			data[89053] <= 8'h10 ;
			data[89054] <= 8'h10 ;
			data[89055] <= 8'h10 ;
			data[89056] <= 8'h10 ;
			data[89057] <= 8'h10 ;
			data[89058] <= 8'h10 ;
			data[89059] <= 8'h10 ;
			data[89060] <= 8'h10 ;
			data[89061] <= 8'h10 ;
			data[89062] <= 8'h10 ;
			data[89063] <= 8'h10 ;
			data[89064] <= 8'h10 ;
			data[89065] <= 8'h10 ;
			data[89066] <= 8'h10 ;
			data[89067] <= 8'h10 ;
			data[89068] <= 8'h10 ;
			data[89069] <= 8'h10 ;
			data[89070] <= 8'h10 ;
			data[89071] <= 8'h10 ;
			data[89072] <= 8'h10 ;
			data[89073] <= 8'h10 ;
			data[89074] <= 8'h10 ;
			data[89075] <= 8'h10 ;
			data[89076] <= 8'h10 ;
			data[89077] <= 8'h10 ;
			data[89078] <= 8'h10 ;
			data[89079] <= 8'h10 ;
			data[89080] <= 8'h10 ;
			data[89081] <= 8'h10 ;
			data[89082] <= 8'h10 ;
			data[89083] <= 8'h10 ;
			data[89084] <= 8'h10 ;
			data[89085] <= 8'h10 ;
			data[89086] <= 8'h10 ;
			data[89087] <= 8'h10 ;
			data[89088] <= 8'h10 ;
			data[89089] <= 8'h10 ;
			data[89090] <= 8'h10 ;
			data[89091] <= 8'h10 ;
			data[89092] <= 8'h10 ;
			data[89093] <= 8'h10 ;
			data[89094] <= 8'h10 ;
			data[89095] <= 8'h10 ;
			data[89096] <= 8'h10 ;
			data[89097] <= 8'h10 ;
			data[89098] <= 8'h10 ;
			data[89099] <= 8'h10 ;
			data[89100] <= 8'h10 ;
			data[89101] <= 8'h10 ;
			data[89102] <= 8'h10 ;
			data[89103] <= 8'h10 ;
			data[89104] <= 8'h10 ;
			data[89105] <= 8'h10 ;
			data[89106] <= 8'h10 ;
			data[89107] <= 8'h10 ;
			data[89108] <= 8'h10 ;
			data[89109] <= 8'h10 ;
			data[89110] <= 8'h10 ;
			data[89111] <= 8'h10 ;
			data[89112] <= 8'h10 ;
			data[89113] <= 8'h10 ;
			data[89114] <= 8'h10 ;
			data[89115] <= 8'h10 ;
			data[89116] <= 8'h10 ;
			data[89117] <= 8'h10 ;
			data[89118] <= 8'h10 ;
			data[89119] <= 8'h10 ;
			data[89120] <= 8'h10 ;
			data[89121] <= 8'h10 ;
			data[89122] <= 8'h10 ;
			data[89123] <= 8'h10 ;
			data[89124] <= 8'h10 ;
			data[89125] <= 8'h10 ;
			data[89126] <= 8'h10 ;
			data[89127] <= 8'h10 ;
			data[89128] <= 8'h10 ;
			data[89129] <= 8'h10 ;
			data[89130] <= 8'h10 ;
			data[89131] <= 8'h10 ;
			data[89132] <= 8'h10 ;
			data[89133] <= 8'h10 ;
			data[89134] <= 8'h10 ;
			data[89135] <= 8'h10 ;
			data[89136] <= 8'h10 ;
			data[89137] <= 8'h10 ;
			data[89138] <= 8'h10 ;
			data[89139] <= 8'h10 ;
			data[89140] <= 8'h10 ;
			data[89141] <= 8'h10 ;
			data[89142] <= 8'h10 ;
			data[89143] <= 8'h10 ;
			data[89144] <= 8'h10 ;
			data[89145] <= 8'h10 ;
			data[89146] <= 8'h10 ;
			data[89147] <= 8'h10 ;
			data[89148] <= 8'h10 ;
			data[89149] <= 8'h10 ;
			data[89150] <= 8'h10 ;
			data[89151] <= 8'h10 ;
			data[89152] <= 8'h10 ;
			data[89153] <= 8'h10 ;
			data[89154] <= 8'h10 ;
			data[89155] <= 8'h10 ;
			data[89156] <= 8'h10 ;
			data[89157] <= 8'h10 ;
			data[89158] <= 8'h10 ;
			data[89159] <= 8'h10 ;
			data[89160] <= 8'h10 ;
			data[89161] <= 8'h10 ;
			data[89162] <= 8'h10 ;
			data[89163] <= 8'h10 ;
			data[89164] <= 8'h10 ;
			data[89165] <= 8'h10 ;
			data[89166] <= 8'h10 ;
			data[89167] <= 8'h10 ;
			data[89168] <= 8'h10 ;
			data[89169] <= 8'h10 ;
			data[89170] <= 8'h10 ;
			data[89171] <= 8'h10 ;
			data[89172] <= 8'h10 ;
			data[89173] <= 8'h10 ;
			data[89174] <= 8'h10 ;
			data[89175] <= 8'h10 ;
			data[89176] <= 8'h10 ;
			data[89177] <= 8'h10 ;
			data[89178] <= 8'h10 ;
			data[89179] <= 8'h10 ;
			data[89180] <= 8'h10 ;
			data[89181] <= 8'h10 ;
			data[89182] <= 8'h10 ;
			data[89183] <= 8'h10 ;
			data[89184] <= 8'h10 ;
			data[89185] <= 8'h10 ;
			data[89186] <= 8'h10 ;
			data[89187] <= 8'h10 ;
			data[89188] <= 8'h10 ;
			data[89189] <= 8'h10 ;
			data[89190] <= 8'h10 ;
			data[89191] <= 8'h10 ;
			data[89192] <= 8'h10 ;
			data[89193] <= 8'h10 ;
			data[89194] <= 8'h10 ;
			data[89195] <= 8'h10 ;
			data[89196] <= 8'h10 ;
			data[89197] <= 8'h10 ;
			data[89198] <= 8'h10 ;
			data[89199] <= 8'h10 ;
			data[89200] <= 8'h10 ;
			data[89201] <= 8'h10 ;
			data[89202] <= 8'h10 ;
			data[89203] <= 8'h10 ;
			data[89204] <= 8'h10 ;
			data[89205] <= 8'h10 ;
			data[89206] <= 8'h10 ;
			data[89207] <= 8'h10 ;
			data[89208] <= 8'h10 ;
			data[89209] <= 8'h10 ;
			data[89210] <= 8'h10 ;
			data[89211] <= 8'h10 ;
			data[89212] <= 8'h10 ;
			data[89213] <= 8'h10 ;
			data[89214] <= 8'h10 ;
			data[89215] <= 8'h10 ;
			data[89216] <= 8'h10 ;
			data[89217] <= 8'h10 ;
			data[89218] <= 8'h10 ;
			data[89219] <= 8'h10 ;
			data[89220] <= 8'h10 ;
			data[89221] <= 8'h10 ;
			data[89222] <= 8'h10 ;
			data[89223] <= 8'h10 ;
			data[89224] <= 8'h10 ;
			data[89225] <= 8'h10 ;
			data[89226] <= 8'h10 ;
			data[89227] <= 8'h10 ;
			data[89228] <= 8'h10 ;
			data[89229] <= 8'h10 ;
			data[89230] <= 8'h10 ;
			data[89231] <= 8'h10 ;
			data[89232] <= 8'h10 ;
			data[89233] <= 8'h10 ;
			data[89234] <= 8'h10 ;
			data[89235] <= 8'h10 ;
			data[89236] <= 8'h10 ;
			data[89237] <= 8'h10 ;
			data[89238] <= 8'h10 ;
			data[89239] <= 8'h10 ;
			data[89240] <= 8'h10 ;
			data[89241] <= 8'h10 ;
			data[89242] <= 8'h10 ;
			data[89243] <= 8'h10 ;
			data[89244] <= 8'h10 ;
			data[89245] <= 8'h10 ;
			data[89246] <= 8'h10 ;
			data[89247] <= 8'h10 ;
			data[89248] <= 8'h10 ;
			data[89249] <= 8'h10 ;
			data[89250] <= 8'h10 ;
			data[89251] <= 8'h10 ;
			data[89252] <= 8'h10 ;
			data[89253] <= 8'h10 ;
			data[89254] <= 8'h10 ;
			data[89255] <= 8'h10 ;
			data[89256] <= 8'h10 ;
			data[89257] <= 8'h10 ;
			data[89258] <= 8'h10 ;
			data[89259] <= 8'h10 ;
			data[89260] <= 8'h10 ;
			data[89261] <= 8'h10 ;
			data[89262] <= 8'h10 ;
			data[89263] <= 8'h10 ;
			data[89264] <= 8'h10 ;
			data[89265] <= 8'h10 ;
			data[89266] <= 8'h10 ;
			data[89267] <= 8'h10 ;
			data[89268] <= 8'h10 ;
			data[89269] <= 8'h10 ;
			data[89270] <= 8'h10 ;
			data[89271] <= 8'h10 ;
			data[89272] <= 8'h10 ;
			data[89273] <= 8'h10 ;
			data[89274] <= 8'h10 ;
			data[89275] <= 8'h10 ;
			data[89276] <= 8'h10 ;
			data[89277] <= 8'h10 ;
			data[89278] <= 8'h10 ;
			data[89279] <= 8'h10 ;
			data[89280] <= 8'h10 ;
			data[89281] <= 8'h10 ;
			data[89282] <= 8'h10 ;
			data[89283] <= 8'h10 ;
			data[89284] <= 8'h10 ;
			data[89285] <= 8'h10 ;
			data[89286] <= 8'h10 ;
			data[89287] <= 8'h10 ;
			data[89288] <= 8'h10 ;
			data[89289] <= 8'h10 ;
			data[89290] <= 8'h10 ;
			data[89291] <= 8'h10 ;
			data[89292] <= 8'h10 ;
			data[89293] <= 8'h10 ;
			data[89294] <= 8'h10 ;
			data[89295] <= 8'h10 ;
			data[89296] <= 8'h10 ;
			data[89297] <= 8'h10 ;
			data[89298] <= 8'h10 ;
			data[89299] <= 8'h10 ;
			data[89300] <= 8'h10 ;
			data[89301] <= 8'h10 ;
			data[89302] <= 8'h10 ;
			data[89303] <= 8'h10 ;
			data[89304] <= 8'h10 ;
			data[89305] <= 8'h10 ;
			data[89306] <= 8'h10 ;
			data[89307] <= 8'h10 ;
			data[89308] <= 8'h10 ;
			data[89309] <= 8'h10 ;
			data[89310] <= 8'h10 ;
			data[89311] <= 8'h10 ;
			data[89312] <= 8'h10 ;
			data[89313] <= 8'h10 ;
			data[89314] <= 8'h10 ;
			data[89315] <= 8'h10 ;
			data[89316] <= 8'h10 ;
			data[89317] <= 8'h10 ;
			data[89318] <= 8'h10 ;
			data[89319] <= 8'h10 ;
			data[89320] <= 8'h10 ;
			data[89321] <= 8'h10 ;
			data[89322] <= 8'h10 ;
			data[89323] <= 8'h10 ;
			data[89324] <= 8'h10 ;
			data[89325] <= 8'h10 ;
			data[89326] <= 8'h10 ;
			data[89327] <= 8'h10 ;
			data[89328] <= 8'h10 ;
			data[89329] <= 8'h10 ;
			data[89330] <= 8'h10 ;
			data[89331] <= 8'h10 ;
			data[89332] <= 8'h10 ;
			data[89333] <= 8'h10 ;
			data[89334] <= 8'h10 ;
			data[89335] <= 8'h10 ;
			data[89336] <= 8'h10 ;
			data[89337] <= 8'h10 ;
			data[89338] <= 8'h10 ;
			data[89339] <= 8'h10 ;
			data[89340] <= 8'h10 ;
			data[89341] <= 8'h10 ;
			data[89342] <= 8'h10 ;
			data[89343] <= 8'h10 ;
			data[89344] <= 8'h10 ;
			data[89345] <= 8'h10 ;
			data[89346] <= 8'h10 ;
			data[89347] <= 8'h10 ;
			data[89348] <= 8'h10 ;
			data[89349] <= 8'h10 ;
			data[89350] <= 8'h10 ;
			data[89351] <= 8'h10 ;
			data[89352] <= 8'h10 ;
			data[89353] <= 8'h10 ;
			data[89354] <= 8'h10 ;
			data[89355] <= 8'h10 ;
			data[89356] <= 8'h10 ;
			data[89357] <= 8'h10 ;
			data[89358] <= 8'h10 ;
			data[89359] <= 8'h10 ;
			data[89360] <= 8'h10 ;
			data[89361] <= 8'h10 ;
			data[89362] <= 8'h10 ;
			data[89363] <= 8'h10 ;
			data[89364] <= 8'h10 ;
			data[89365] <= 8'h10 ;
			data[89366] <= 8'h10 ;
			data[89367] <= 8'h10 ;
			data[89368] <= 8'h10 ;
			data[89369] <= 8'h10 ;
			data[89370] <= 8'h10 ;
			data[89371] <= 8'h10 ;
			data[89372] <= 8'h10 ;
			data[89373] <= 8'h10 ;
			data[89374] <= 8'h10 ;
			data[89375] <= 8'h10 ;
			data[89376] <= 8'h10 ;
			data[89377] <= 8'h10 ;
			data[89378] <= 8'h10 ;
			data[89379] <= 8'h10 ;
			data[89380] <= 8'h10 ;
			data[89381] <= 8'h10 ;
			data[89382] <= 8'h10 ;
			data[89383] <= 8'h10 ;
			data[89384] <= 8'h10 ;
			data[89385] <= 8'h10 ;
			data[89386] <= 8'h10 ;
			data[89387] <= 8'h10 ;
			data[89388] <= 8'h10 ;
			data[89389] <= 8'h10 ;
			data[89390] <= 8'h10 ;
			data[89391] <= 8'h10 ;
			data[89392] <= 8'h10 ;
			data[89393] <= 8'h10 ;
			data[89394] <= 8'h10 ;
			data[89395] <= 8'h10 ;
			data[89396] <= 8'h10 ;
			data[89397] <= 8'h10 ;
			data[89398] <= 8'h10 ;
			data[89399] <= 8'h10 ;
			data[89400] <= 8'h10 ;
			data[89401] <= 8'h10 ;
			data[89402] <= 8'h10 ;
			data[89403] <= 8'h10 ;
			data[89404] <= 8'h10 ;
			data[89405] <= 8'h10 ;
			data[89406] <= 8'h10 ;
			data[89407] <= 8'h10 ;
			data[89408] <= 8'h10 ;
			data[89409] <= 8'h10 ;
			data[89410] <= 8'h10 ;
			data[89411] <= 8'h10 ;
			data[89412] <= 8'h10 ;
			data[89413] <= 8'h10 ;
			data[89414] <= 8'h10 ;
			data[89415] <= 8'h10 ;
			data[89416] <= 8'h10 ;
			data[89417] <= 8'h10 ;
			data[89418] <= 8'h10 ;
			data[89419] <= 8'h10 ;
			data[89420] <= 8'h10 ;
			data[89421] <= 8'h10 ;
			data[89422] <= 8'h10 ;
			data[89423] <= 8'h10 ;
			data[89424] <= 8'h10 ;
			data[89425] <= 8'h10 ;
			data[89426] <= 8'h10 ;
			data[89427] <= 8'h10 ;
			data[89428] <= 8'h10 ;
			data[89429] <= 8'h10 ;
			data[89430] <= 8'h10 ;
			data[89431] <= 8'h10 ;
			data[89432] <= 8'h10 ;
			data[89433] <= 8'h10 ;
			data[89434] <= 8'h10 ;
			data[89435] <= 8'h10 ;
			data[89436] <= 8'h10 ;
			data[89437] <= 8'h10 ;
			data[89438] <= 8'h10 ;
			data[89439] <= 8'h10 ;
			data[89440] <= 8'h10 ;
			data[89441] <= 8'h10 ;
			data[89442] <= 8'h10 ;
			data[89443] <= 8'h10 ;
			data[89444] <= 8'h10 ;
			data[89445] <= 8'h10 ;
			data[89446] <= 8'h10 ;
			data[89447] <= 8'h10 ;
			data[89448] <= 8'h10 ;
			data[89449] <= 8'h10 ;
			data[89450] <= 8'h10 ;
			data[89451] <= 8'h10 ;
			data[89452] <= 8'h10 ;
			data[89453] <= 8'h10 ;
			data[89454] <= 8'h10 ;
			data[89455] <= 8'h10 ;
			data[89456] <= 8'h10 ;
			data[89457] <= 8'h10 ;
			data[89458] <= 8'h10 ;
			data[89459] <= 8'h10 ;
			data[89460] <= 8'h10 ;
			data[89461] <= 8'h10 ;
			data[89462] <= 8'h10 ;
			data[89463] <= 8'h10 ;
			data[89464] <= 8'h10 ;
			data[89465] <= 8'h10 ;
			data[89466] <= 8'h10 ;
			data[89467] <= 8'h10 ;
			data[89468] <= 8'h10 ;
			data[89469] <= 8'h10 ;
			data[89470] <= 8'h10 ;
			data[89471] <= 8'h10 ;
			data[89472] <= 8'h10 ;
			data[89473] <= 8'h10 ;
			data[89474] <= 8'h10 ;
			data[89475] <= 8'h10 ;
			data[89476] <= 8'h10 ;
			data[89477] <= 8'h10 ;
			data[89478] <= 8'h10 ;
			data[89479] <= 8'h10 ;
			data[89480] <= 8'h10 ;
			data[89481] <= 8'h10 ;
			data[89482] <= 8'h10 ;
			data[89483] <= 8'h10 ;
			data[89484] <= 8'h10 ;
			data[89485] <= 8'h10 ;
			data[89486] <= 8'h10 ;
			data[89487] <= 8'h10 ;
			data[89488] <= 8'h10 ;
			data[89489] <= 8'h10 ;
			data[89490] <= 8'h10 ;
			data[89491] <= 8'h10 ;
			data[89492] <= 8'h10 ;
			data[89493] <= 8'h10 ;
			data[89494] <= 8'h10 ;
			data[89495] <= 8'h10 ;
			data[89496] <= 8'h10 ;
			data[89497] <= 8'h10 ;
			data[89498] <= 8'h10 ;
			data[89499] <= 8'h10 ;
			data[89500] <= 8'h10 ;
			data[89501] <= 8'h10 ;
			data[89502] <= 8'h10 ;
			data[89503] <= 8'h10 ;
			data[89504] <= 8'h10 ;
			data[89505] <= 8'h10 ;
			data[89506] <= 8'h10 ;
			data[89507] <= 8'h10 ;
			data[89508] <= 8'h10 ;
			data[89509] <= 8'h10 ;
			data[89510] <= 8'h10 ;
			data[89511] <= 8'h10 ;
			data[89512] <= 8'h10 ;
			data[89513] <= 8'h10 ;
			data[89514] <= 8'h10 ;
			data[89515] <= 8'h10 ;
			data[89516] <= 8'h10 ;
			data[89517] <= 8'h10 ;
			data[89518] <= 8'h10 ;
			data[89519] <= 8'h10 ;
			data[89520] <= 8'h10 ;
			data[89521] <= 8'h10 ;
			data[89522] <= 8'h10 ;
			data[89523] <= 8'h10 ;
			data[89524] <= 8'h10 ;
			data[89525] <= 8'h10 ;
			data[89526] <= 8'h10 ;
			data[89527] <= 8'h10 ;
			data[89528] <= 8'h10 ;
			data[89529] <= 8'h10 ;
			data[89530] <= 8'h10 ;
			data[89531] <= 8'h10 ;
			data[89532] <= 8'h10 ;
			data[89533] <= 8'h10 ;
			data[89534] <= 8'h10 ;
			data[89535] <= 8'h10 ;
			data[89536] <= 8'h10 ;
			data[89537] <= 8'h10 ;
			data[89538] <= 8'h10 ;
			data[89539] <= 8'h10 ;
			data[89540] <= 8'h10 ;
			data[89541] <= 8'h10 ;
			data[89542] <= 8'h10 ;
			data[89543] <= 8'h10 ;
			data[89544] <= 8'h10 ;
			data[89545] <= 8'h10 ;
			data[89546] <= 8'h10 ;
			data[89547] <= 8'h10 ;
			data[89548] <= 8'h10 ;
			data[89549] <= 8'h10 ;
			data[89550] <= 8'h10 ;
			data[89551] <= 8'h10 ;
			data[89552] <= 8'h10 ;
			data[89553] <= 8'h10 ;
			data[89554] <= 8'h10 ;
			data[89555] <= 8'h10 ;
			data[89556] <= 8'h10 ;
			data[89557] <= 8'h10 ;
			data[89558] <= 8'h10 ;
			data[89559] <= 8'h10 ;
			data[89560] <= 8'h10 ;
			data[89561] <= 8'h10 ;
			data[89562] <= 8'h10 ;
			data[89563] <= 8'h10 ;
			data[89564] <= 8'h10 ;
			data[89565] <= 8'h10 ;
			data[89566] <= 8'h10 ;
			data[89567] <= 8'h10 ;
			data[89568] <= 8'h10 ;
			data[89569] <= 8'h10 ;
			data[89570] <= 8'h10 ;
			data[89571] <= 8'h10 ;
			data[89572] <= 8'h10 ;
			data[89573] <= 8'h10 ;
			data[89574] <= 8'h10 ;
			data[89575] <= 8'h10 ;
			data[89576] <= 8'h10 ;
			data[89577] <= 8'h10 ;
			data[89578] <= 8'h10 ;
			data[89579] <= 8'h10 ;
			data[89580] <= 8'h10 ;
			data[89581] <= 8'h10 ;
			data[89582] <= 8'h10 ;
			data[89583] <= 8'h10 ;
			data[89584] <= 8'h10 ;
			data[89585] <= 8'h10 ;
			data[89586] <= 8'h10 ;
			data[89587] <= 8'h10 ;
			data[89588] <= 8'h10 ;
			data[89589] <= 8'h10 ;
			data[89590] <= 8'h10 ;
			data[89591] <= 8'h10 ;
			data[89592] <= 8'h10 ;
			data[89593] <= 8'h10 ;
			data[89594] <= 8'h10 ;
			data[89595] <= 8'h10 ;
			data[89596] <= 8'h10 ;
			data[89597] <= 8'h10 ;
			data[89598] <= 8'h10 ;
			data[89599] <= 8'h10 ;
			data[89600] <= 8'h10 ;
			data[89601] <= 8'h10 ;
			data[89602] <= 8'h10 ;
			data[89603] <= 8'h10 ;
			data[89604] <= 8'h10 ;
			data[89605] <= 8'h10 ;
			data[89606] <= 8'h10 ;
			data[89607] <= 8'h10 ;
			data[89608] <= 8'h10 ;
			data[89609] <= 8'h10 ;
			data[89610] <= 8'h10 ;
			data[89611] <= 8'h10 ;
			data[89612] <= 8'h10 ;
			data[89613] <= 8'h10 ;
			data[89614] <= 8'h10 ;
			data[89615] <= 8'h10 ;
			data[89616] <= 8'h10 ;
			data[89617] <= 8'h10 ;
			data[89618] <= 8'h10 ;
			data[89619] <= 8'h10 ;
			data[89620] <= 8'h10 ;
			data[89621] <= 8'h10 ;
			data[89622] <= 8'h10 ;
			data[89623] <= 8'h10 ;
			data[89624] <= 8'h10 ;
			data[89625] <= 8'h10 ;
			data[89626] <= 8'h10 ;
			data[89627] <= 8'h10 ;
			data[89628] <= 8'h10 ;
			data[89629] <= 8'h10 ;
			data[89630] <= 8'h10 ;
			data[89631] <= 8'h10 ;
			data[89632] <= 8'h10 ;
			data[89633] <= 8'h10 ;
			data[89634] <= 8'h10 ;
			data[89635] <= 8'h10 ;
			data[89636] <= 8'h10 ;
			data[89637] <= 8'h10 ;
			data[89638] <= 8'h10 ;
			data[89639] <= 8'h10 ;
			data[89640] <= 8'h10 ;
			data[89641] <= 8'h10 ;
			data[89642] <= 8'h10 ;
			data[89643] <= 8'h10 ;
			data[89644] <= 8'h10 ;
			data[89645] <= 8'h10 ;
			data[89646] <= 8'h10 ;
			data[89647] <= 8'h10 ;
			data[89648] <= 8'h10 ;
			data[89649] <= 8'h10 ;
			data[89650] <= 8'h10 ;
			data[89651] <= 8'h10 ;
			data[89652] <= 8'h10 ;
			data[89653] <= 8'h10 ;
			data[89654] <= 8'h10 ;
			data[89655] <= 8'h10 ;
			data[89656] <= 8'h10 ;
			data[89657] <= 8'h10 ;
			data[89658] <= 8'h10 ;
			data[89659] <= 8'h10 ;
			data[89660] <= 8'h10 ;
			data[89661] <= 8'h10 ;
			data[89662] <= 8'h10 ;
			data[89663] <= 8'h10 ;
			data[89664] <= 8'h10 ;
			data[89665] <= 8'h10 ;
			data[89666] <= 8'h10 ;
			data[89667] <= 8'h10 ;
			data[89668] <= 8'h10 ;
			data[89669] <= 8'h10 ;
			data[89670] <= 8'h10 ;
			data[89671] <= 8'h10 ;
			data[89672] <= 8'h10 ;
			data[89673] <= 8'h10 ;
			data[89674] <= 8'h10 ;
			data[89675] <= 8'h10 ;
			data[89676] <= 8'h10 ;
			data[89677] <= 8'h10 ;
			data[89678] <= 8'h10 ;
			data[89679] <= 8'h10 ;
			data[89680] <= 8'h10 ;
			data[89681] <= 8'h10 ;
			data[89682] <= 8'h10 ;
			data[89683] <= 8'h10 ;
			data[89684] <= 8'h10 ;
			data[89685] <= 8'h10 ;
			data[89686] <= 8'h10 ;
			data[89687] <= 8'h10 ;
			data[89688] <= 8'h10 ;
			data[89689] <= 8'h10 ;
			data[89690] <= 8'h10 ;
			data[89691] <= 8'h10 ;
			data[89692] <= 8'h10 ;
			data[89693] <= 8'h10 ;
			data[89694] <= 8'h10 ;
			data[89695] <= 8'h10 ;
			data[89696] <= 8'h10 ;
			data[89697] <= 8'h10 ;
			data[89698] <= 8'h10 ;
			data[89699] <= 8'h10 ;
			data[89700] <= 8'h10 ;
			data[89701] <= 8'h10 ;
			data[89702] <= 8'h10 ;
			data[89703] <= 8'h10 ;
			data[89704] <= 8'h10 ;
			data[89705] <= 8'h10 ;
			data[89706] <= 8'h10 ;
			data[89707] <= 8'h10 ;
			data[89708] <= 8'h10 ;
			data[89709] <= 8'h10 ;
			data[89710] <= 8'h10 ;
			data[89711] <= 8'h10 ;
			data[89712] <= 8'h10 ;
			data[89713] <= 8'h10 ;
			data[89714] <= 8'h10 ;
			data[89715] <= 8'h10 ;
			data[89716] <= 8'h10 ;
			data[89717] <= 8'h10 ;
			data[89718] <= 8'h10 ;
			data[89719] <= 8'h10 ;
			data[89720] <= 8'h10 ;
			data[89721] <= 8'h10 ;
			data[89722] <= 8'h10 ;
			data[89723] <= 8'h10 ;
			data[89724] <= 8'h10 ;
			data[89725] <= 8'h10 ;
			data[89726] <= 8'h10 ;
			data[89727] <= 8'h10 ;
			data[89728] <= 8'h10 ;
			data[89729] <= 8'h10 ;
			data[89730] <= 8'h10 ;
			data[89731] <= 8'h10 ;
			data[89732] <= 8'h10 ;
			data[89733] <= 8'h10 ;
			data[89734] <= 8'h10 ;
			data[89735] <= 8'h10 ;
			data[89736] <= 8'h10 ;
			data[89737] <= 8'h10 ;
			data[89738] <= 8'h10 ;
			data[89739] <= 8'h10 ;
			data[89740] <= 8'h10 ;
			data[89741] <= 8'h10 ;
			data[89742] <= 8'h10 ;
			data[89743] <= 8'h10 ;
			data[89744] <= 8'h10 ;
			data[89745] <= 8'h10 ;
			data[89746] <= 8'h10 ;
			data[89747] <= 8'h10 ;
			data[89748] <= 8'h10 ;
			data[89749] <= 8'h10 ;
			data[89750] <= 8'h10 ;
			data[89751] <= 8'h10 ;
			data[89752] <= 8'h10 ;
			data[89753] <= 8'h10 ;
			data[89754] <= 8'h10 ;
			data[89755] <= 8'h10 ;
			data[89756] <= 8'h10 ;
			data[89757] <= 8'h10 ;
			data[89758] <= 8'h10 ;
			data[89759] <= 8'h10 ;
			data[89760] <= 8'h10 ;
			data[89761] <= 8'h10 ;
			data[89762] <= 8'h10 ;
			data[89763] <= 8'h10 ;
			data[89764] <= 8'h10 ;
			data[89765] <= 8'h10 ;
			data[89766] <= 8'h10 ;
			data[89767] <= 8'h10 ;
			data[89768] <= 8'h10 ;
			data[89769] <= 8'h10 ;
			data[89770] <= 8'h10 ;
			data[89771] <= 8'h10 ;
			data[89772] <= 8'h10 ;
			data[89773] <= 8'h10 ;
			data[89774] <= 8'h10 ;
			data[89775] <= 8'h10 ;
			data[89776] <= 8'h10 ;
			data[89777] <= 8'h10 ;
			data[89778] <= 8'h10 ;
			data[89779] <= 8'h10 ;
			data[89780] <= 8'h10 ;
			data[89781] <= 8'h10 ;
			data[89782] <= 8'h10 ;
			data[89783] <= 8'h10 ;
			data[89784] <= 8'h10 ;
			data[89785] <= 8'h10 ;
			data[89786] <= 8'h10 ;
			data[89787] <= 8'h10 ;
			data[89788] <= 8'h10 ;
			data[89789] <= 8'h10 ;
			data[89790] <= 8'h10 ;
			data[89791] <= 8'h10 ;
			data[89792] <= 8'h10 ;
			data[89793] <= 8'h10 ;
			data[89794] <= 8'h10 ;
			data[89795] <= 8'h10 ;
			data[89796] <= 8'h10 ;
			data[89797] <= 8'h10 ;
			data[89798] <= 8'h10 ;
			data[89799] <= 8'h10 ;
			data[89800] <= 8'h10 ;
			data[89801] <= 8'h10 ;
			data[89802] <= 8'h10 ;
			data[89803] <= 8'h10 ;
			data[89804] <= 8'h10 ;
			data[89805] <= 8'h10 ;
			data[89806] <= 8'h10 ;
			data[89807] <= 8'h10 ;
			data[89808] <= 8'h10 ;
			data[89809] <= 8'h10 ;
			data[89810] <= 8'h10 ;
			data[89811] <= 8'h10 ;
			data[89812] <= 8'h10 ;
			data[89813] <= 8'h10 ;
			data[89814] <= 8'h10 ;
			data[89815] <= 8'h10 ;
			data[89816] <= 8'h10 ;
			data[89817] <= 8'h10 ;
			data[89818] <= 8'h10 ;
			data[89819] <= 8'h10 ;
			data[89820] <= 8'h10 ;
			data[89821] <= 8'h10 ;
			data[89822] <= 8'h10 ;
			data[89823] <= 8'h10 ;
			data[89824] <= 8'h10 ;
			data[89825] <= 8'h10 ;
			data[89826] <= 8'h10 ;
			data[89827] <= 8'h10 ;
			data[89828] <= 8'h10 ;
			data[89829] <= 8'h10 ;
			data[89830] <= 8'h10 ;
			data[89831] <= 8'h10 ;
			data[89832] <= 8'h10 ;
			data[89833] <= 8'h10 ;
			data[89834] <= 8'h10 ;
			data[89835] <= 8'h10 ;
			data[89836] <= 8'h10 ;
			data[89837] <= 8'h10 ;
			data[89838] <= 8'h10 ;
			data[89839] <= 8'h10 ;
			data[89840] <= 8'h10 ;
			data[89841] <= 8'h10 ;
			data[89842] <= 8'h10 ;
			data[89843] <= 8'h10 ;
			data[89844] <= 8'h10 ;
			data[89845] <= 8'h10 ;
			data[89846] <= 8'h10 ;
			data[89847] <= 8'h10 ;
			data[89848] <= 8'h10 ;
			data[89849] <= 8'h10 ;
			data[89850] <= 8'h10 ;
			data[89851] <= 8'h10 ;
			data[89852] <= 8'h10 ;
			data[89853] <= 8'h10 ;
			data[89854] <= 8'h10 ;
			data[89855] <= 8'h10 ;
			data[89856] <= 8'h10 ;
			data[89857] <= 8'h10 ;
			data[89858] <= 8'h10 ;
			data[89859] <= 8'h10 ;
			data[89860] <= 8'h10 ;
			data[89861] <= 8'h10 ;
			data[89862] <= 8'h10 ;
			data[89863] <= 8'h10 ;
			data[89864] <= 8'h10 ;
			data[89865] <= 8'h10 ;
			data[89866] <= 8'h10 ;
			data[89867] <= 8'h10 ;
			data[89868] <= 8'h10 ;
			data[89869] <= 8'h10 ;
			data[89870] <= 8'h10 ;
			data[89871] <= 8'h10 ;
			data[89872] <= 8'h10 ;
			data[89873] <= 8'h10 ;
			data[89874] <= 8'h10 ;
			data[89875] <= 8'h10 ;
			data[89876] <= 8'h10 ;
			data[89877] <= 8'h10 ;
			data[89878] <= 8'h10 ;
			data[89879] <= 8'h10 ;
			data[89880] <= 8'h10 ;
			data[89881] <= 8'h10 ;
			data[89882] <= 8'h10 ;
			data[89883] <= 8'h10 ;
			data[89884] <= 8'h10 ;
			data[89885] <= 8'h10 ;
			data[89886] <= 8'h10 ;
			data[89887] <= 8'h10 ;
			data[89888] <= 8'h10 ;
			data[89889] <= 8'h10 ;
			data[89890] <= 8'h10 ;
			data[89891] <= 8'h10 ;
			data[89892] <= 8'h10 ;
			data[89893] <= 8'h10 ;
			data[89894] <= 8'h10 ;
			data[89895] <= 8'h10 ;
			data[89896] <= 8'h10 ;
			data[89897] <= 8'h10 ;
			data[89898] <= 8'h10 ;
			data[89899] <= 8'h10 ;
			data[89900] <= 8'h10 ;
			data[89901] <= 8'h10 ;
			data[89902] <= 8'h10 ;
			data[89903] <= 8'h10 ;
			data[89904] <= 8'h10 ;
			data[89905] <= 8'h10 ;
			data[89906] <= 8'h10 ;
			data[89907] <= 8'h10 ;
			data[89908] <= 8'h10 ;
			data[89909] <= 8'h10 ;
			data[89910] <= 8'h10 ;
			data[89911] <= 8'h10 ;
			data[89912] <= 8'h10 ;
			data[89913] <= 8'h10 ;
			data[89914] <= 8'h10 ;
			data[89915] <= 8'h10 ;
			data[89916] <= 8'h10 ;
			data[89917] <= 8'h10 ;
			data[89918] <= 8'h10 ;
			data[89919] <= 8'h10 ;
			data[89920] <= 8'h10 ;
			data[89921] <= 8'h10 ;
			data[89922] <= 8'h10 ;
			data[89923] <= 8'h10 ;
			data[89924] <= 8'h10 ;
			data[89925] <= 8'h10 ;
			data[89926] <= 8'h10 ;
			data[89927] <= 8'h10 ;
			data[89928] <= 8'h10 ;
			data[89929] <= 8'h10 ;
			data[89930] <= 8'h10 ;
			data[89931] <= 8'h10 ;
			data[89932] <= 8'h10 ;
			data[89933] <= 8'h10 ;
			data[89934] <= 8'h10 ;
			data[89935] <= 8'h10 ;
			data[89936] <= 8'h10 ;
			data[89937] <= 8'h10 ;
			data[89938] <= 8'h10 ;
			data[89939] <= 8'h10 ;
			data[89940] <= 8'h10 ;
			data[89941] <= 8'h10 ;
			data[89942] <= 8'h10 ;
			data[89943] <= 8'h10 ;
			data[89944] <= 8'h10 ;
			data[89945] <= 8'h10 ;
			data[89946] <= 8'h10 ;
			data[89947] <= 8'h10 ;
			data[89948] <= 8'h10 ;
			data[89949] <= 8'h10 ;
			data[89950] <= 8'h10 ;
			data[89951] <= 8'h10 ;
			data[89952] <= 8'h10 ;
			data[89953] <= 8'h10 ;
			data[89954] <= 8'h10 ;
			data[89955] <= 8'h10 ;
			data[89956] <= 8'h10 ;
			data[89957] <= 8'h10 ;
			data[89958] <= 8'h10 ;
			data[89959] <= 8'h10 ;
			data[89960] <= 8'h10 ;
			data[89961] <= 8'h10 ;
			data[89962] <= 8'h10 ;
			data[89963] <= 8'h10 ;
			data[89964] <= 8'h10 ;
			data[89965] <= 8'h10 ;
			data[89966] <= 8'h10 ;
			data[89967] <= 8'h10 ;
			data[89968] <= 8'h10 ;
			data[89969] <= 8'h10 ;
			data[89970] <= 8'h10 ;
			data[89971] <= 8'h10 ;
			data[89972] <= 8'h10 ;
			data[89973] <= 8'h10 ;
			data[89974] <= 8'h10 ;
			data[89975] <= 8'h10 ;
			data[89976] <= 8'h10 ;
			data[89977] <= 8'h10 ;
			data[89978] <= 8'h10 ;
			data[89979] <= 8'h10 ;
			data[89980] <= 8'h10 ;
			data[89981] <= 8'h10 ;
			data[89982] <= 8'h10 ;
			data[89983] <= 8'h10 ;
			data[89984] <= 8'h10 ;
			data[89985] <= 8'h10 ;
			data[89986] <= 8'h10 ;
			data[89987] <= 8'h10 ;
			data[89988] <= 8'h10 ;
			data[89989] <= 8'h10 ;
			data[89990] <= 8'h10 ;
			data[89991] <= 8'h10 ;
			data[89992] <= 8'h10 ;
			data[89993] <= 8'h10 ;
			data[89994] <= 8'h10 ;
			data[89995] <= 8'h10 ;
			data[89996] <= 8'h10 ;
			data[89997] <= 8'h10 ;
			data[89998] <= 8'h10 ;
			data[89999] <= 8'h10 ;
			data[90000] <= 8'h10 ;
			data[90001] <= 8'h10 ;
			data[90002] <= 8'h10 ;
			data[90003] <= 8'h10 ;
			data[90004] <= 8'h10 ;
			data[90005] <= 8'h10 ;
			data[90006] <= 8'h10 ;
			data[90007] <= 8'h10 ;
			data[90008] <= 8'h10 ;
			data[90009] <= 8'h10 ;
			data[90010] <= 8'h10 ;
			data[90011] <= 8'h10 ;
			data[90012] <= 8'h10 ;
			data[90013] <= 8'h10 ;
			data[90014] <= 8'h10 ;
			data[90015] <= 8'h10 ;
			data[90016] <= 8'h10 ;
			data[90017] <= 8'h10 ;
			data[90018] <= 8'h10 ;
			data[90019] <= 8'h10 ;
			data[90020] <= 8'h10 ;
			data[90021] <= 8'h10 ;
			data[90022] <= 8'h10 ;
			data[90023] <= 8'h10 ;
			data[90024] <= 8'h10 ;
			data[90025] <= 8'h10 ;
			data[90026] <= 8'h10 ;
			data[90027] <= 8'h10 ;
			data[90028] <= 8'h10 ;
			data[90029] <= 8'h10 ;
			data[90030] <= 8'h10 ;
			data[90031] <= 8'h10 ;
			data[90032] <= 8'h10 ;
			data[90033] <= 8'h10 ;
			data[90034] <= 8'h10 ;
			data[90035] <= 8'h10 ;
			data[90036] <= 8'h10 ;
			data[90037] <= 8'h10 ;
			data[90038] <= 8'h10 ;
			data[90039] <= 8'h10 ;
			data[90040] <= 8'h10 ;
			data[90041] <= 8'h10 ;
			data[90042] <= 8'h10 ;
			data[90043] <= 8'h10 ;
			data[90044] <= 8'h10 ;
			data[90045] <= 8'h10 ;
			data[90046] <= 8'h10 ;
			data[90047] <= 8'h10 ;
			data[90048] <= 8'h10 ;
			data[90049] <= 8'h10 ;
			data[90050] <= 8'h10 ;
			data[90051] <= 8'h10 ;
			data[90052] <= 8'h10 ;
			data[90053] <= 8'h10 ;
			data[90054] <= 8'h10 ;
			data[90055] <= 8'h10 ;
			data[90056] <= 8'h10 ;
			data[90057] <= 8'h10 ;
			data[90058] <= 8'h10 ;
			data[90059] <= 8'h10 ;
			data[90060] <= 8'h10 ;
			data[90061] <= 8'h10 ;
			data[90062] <= 8'h10 ;
			data[90063] <= 8'h10 ;
			data[90064] <= 8'h10 ;
			data[90065] <= 8'h10 ;
			data[90066] <= 8'h10 ;
			data[90067] <= 8'h10 ;
			data[90068] <= 8'h10 ;
			data[90069] <= 8'h10 ;
			data[90070] <= 8'h10 ;
			data[90071] <= 8'h10 ;
			data[90072] <= 8'h10 ;
			data[90073] <= 8'h10 ;
			data[90074] <= 8'h10 ;
			data[90075] <= 8'h10 ;
			data[90076] <= 8'h10 ;
			data[90077] <= 8'h10 ;
			data[90078] <= 8'h10 ;
			data[90079] <= 8'h10 ;
			data[90080] <= 8'h10 ;
			data[90081] <= 8'h10 ;
			data[90082] <= 8'h10 ;
			data[90083] <= 8'h10 ;
			data[90084] <= 8'h10 ;
			data[90085] <= 8'h10 ;
			data[90086] <= 8'h10 ;
			data[90087] <= 8'h10 ;
			data[90088] <= 8'h10 ;
			data[90089] <= 8'h10 ;
			data[90090] <= 8'h10 ;
			data[90091] <= 8'h10 ;
			data[90092] <= 8'h10 ;
			data[90093] <= 8'h10 ;
			data[90094] <= 8'h10 ;
			data[90095] <= 8'h10 ;
			data[90096] <= 8'h10 ;
			data[90097] <= 8'h10 ;
			data[90098] <= 8'h10 ;
			data[90099] <= 8'h10 ;
			data[90100] <= 8'h10 ;
			data[90101] <= 8'h10 ;
			data[90102] <= 8'h10 ;
			data[90103] <= 8'h10 ;
			data[90104] <= 8'h10 ;
			data[90105] <= 8'h10 ;
			data[90106] <= 8'h10 ;
			data[90107] <= 8'h10 ;
			data[90108] <= 8'h10 ;
			data[90109] <= 8'h10 ;
			data[90110] <= 8'h10 ;
			data[90111] <= 8'h10 ;
			data[90112] <= 8'h10 ;
			data[90113] <= 8'h10 ;
			data[90114] <= 8'h10 ;
			data[90115] <= 8'h10 ;
			data[90116] <= 8'h10 ;
			data[90117] <= 8'h10 ;
			data[90118] <= 8'h10 ;
			data[90119] <= 8'h10 ;
			data[90120] <= 8'h10 ;
			data[90121] <= 8'h10 ;
			data[90122] <= 8'h10 ;
			data[90123] <= 8'h10 ;
			data[90124] <= 8'h10 ;
			data[90125] <= 8'h10 ;
			data[90126] <= 8'h10 ;
			data[90127] <= 8'h10 ;
			data[90128] <= 8'h10 ;
			data[90129] <= 8'h10 ;
			data[90130] <= 8'h10 ;
			data[90131] <= 8'h10 ;
			data[90132] <= 8'h10 ;
			data[90133] <= 8'h10 ;
			data[90134] <= 8'h10 ;
			data[90135] <= 8'h10 ;
			data[90136] <= 8'h10 ;
			data[90137] <= 8'h10 ;
			data[90138] <= 8'h10 ;
			data[90139] <= 8'h10 ;
			data[90140] <= 8'h10 ;
			data[90141] <= 8'h10 ;
			data[90142] <= 8'h10 ;
			data[90143] <= 8'h10 ;
			data[90144] <= 8'h10 ;
			data[90145] <= 8'h10 ;
			data[90146] <= 8'h10 ;
			data[90147] <= 8'h10 ;
			data[90148] <= 8'h10 ;
			data[90149] <= 8'h10 ;
			data[90150] <= 8'h10 ;
			data[90151] <= 8'h10 ;
			data[90152] <= 8'h10 ;
			data[90153] <= 8'h10 ;
			data[90154] <= 8'h10 ;
			data[90155] <= 8'h10 ;
			data[90156] <= 8'h10 ;
			data[90157] <= 8'h10 ;
			data[90158] <= 8'h10 ;
			data[90159] <= 8'h10 ;
			data[90160] <= 8'h10 ;
			data[90161] <= 8'h10 ;
			data[90162] <= 8'h10 ;
			data[90163] <= 8'h10 ;
			data[90164] <= 8'h10 ;
			data[90165] <= 8'h10 ;
			data[90166] <= 8'h10 ;
			data[90167] <= 8'h10 ;
			data[90168] <= 8'h10 ;
			data[90169] <= 8'h10 ;
			data[90170] <= 8'h10 ;
			data[90171] <= 8'h10 ;
			data[90172] <= 8'h10 ;
			data[90173] <= 8'h10 ;
			data[90174] <= 8'h10 ;
			data[90175] <= 8'h10 ;
			data[90176] <= 8'h10 ;
			data[90177] <= 8'h10 ;
			data[90178] <= 8'h10 ;
			data[90179] <= 8'h10 ;
			data[90180] <= 8'h10 ;
			data[90181] <= 8'h10 ;
			data[90182] <= 8'h10 ;
			data[90183] <= 8'h10 ;
			data[90184] <= 8'h10 ;
			data[90185] <= 8'h10 ;
			data[90186] <= 8'h10 ;
			data[90187] <= 8'h10 ;
			data[90188] <= 8'h10 ;
			data[90189] <= 8'h10 ;
			data[90190] <= 8'h10 ;
			data[90191] <= 8'h10 ;
			data[90192] <= 8'h10 ;
			data[90193] <= 8'h10 ;
			data[90194] <= 8'h10 ;
			data[90195] <= 8'h10 ;
			data[90196] <= 8'h10 ;
			data[90197] <= 8'h10 ;
			data[90198] <= 8'h10 ;
			data[90199] <= 8'h10 ;
			data[90200] <= 8'h10 ;
			data[90201] <= 8'h10 ;
			data[90202] <= 8'h10 ;
			data[90203] <= 8'h10 ;
			data[90204] <= 8'h10 ;
			data[90205] <= 8'h10 ;
			data[90206] <= 8'h10 ;
			data[90207] <= 8'h10 ;
			data[90208] <= 8'h10 ;
			data[90209] <= 8'h10 ;
			data[90210] <= 8'h10 ;
			data[90211] <= 8'h10 ;
			data[90212] <= 8'h10 ;
			data[90213] <= 8'h10 ;
			data[90214] <= 8'h10 ;
			data[90215] <= 8'h10 ;
			data[90216] <= 8'h10 ;
			data[90217] <= 8'h10 ;
			data[90218] <= 8'h10 ;
			data[90219] <= 8'h10 ;
			data[90220] <= 8'h10 ;
			data[90221] <= 8'h10 ;
			data[90222] <= 8'h10 ;
			data[90223] <= 8'h10 ;
			data[90224] <= 8'h10 ;
			data[90225] <= 8'h10 ;
			data[90226] <= 8'h10 ;
			data[90227] <= 8'h10 ;
			data[90228] <= 8'h10 ;
			data[90229] <= 8'h10 ;
			data[90230] <= 8'h10 ;
			data[90231] <= 8'h10 ;
			data[90232] <= 8'h10 ;
			data[90233] <= 8'h10 ;
			data[90234] <= 8'h10 ;
			data[90235] <= 8'h10 ;
			data[90236] <= 8'h10 ;
			data[90237] <= 8'h10 ;
			data[90238] <= 8'h10 ;
			data[90239] <= 8'h10 ;
			data[90240] <= 8'h10 ;
			data[90241] <= 8'h10 ;
			data[90242] <= 8'h10 ;
			data[90243] <= 8'h10 ;
			data[90244] <= 8'h10 ;
			data[90245] <= 8'h10 ;
			data[90246] <= 8'h10 ;
			data[90247] <= 8'h10 ;
			data[90248] <= 8'h10 ;
			data[90249] <= 8'h10 ;
			data[90250] <= 8'h10 ;
			data[90251] <= 8'h10 ;
			data[90252] <= 8'h10 ;
			data[90253] <= 8'h10 ;
			data[90254] <= 8'h10 ;
			data[90255] <= 8'h10 ;
			data[90256] <= 8'h10 ;
			data[90257] <= 8'h10 ;
			data[90258] <= 8'h10 ;
			data[90259] <= 8'h10 ;
			data[90260] <= 8'h10 ;
			data[90261] <= 8'h10 ;
			data[90262] <= 8'h10 ;
			data[90263] <= 8'h10 ;
			data[90264] <= 8'h10 ;
			data[90265] <= 8'h10 ;
			data[90266] <= 8'h10 ;
			data[90267] <= 8'h10 ;
			data[90268] <= 8'h10 ;
			data[90269] <= 8'h10 ;
			data[90270] <= 8'h10 ;
			data[90271] <= 8'h10 ;
			data[90272] <= 8'h10 ;
			data[90273] <= 8'h10 ;
			data[90274] <= 8'h10 ;
			data[90275] <= 8'h10 ;
			data[90276] <= 8'h10 ;
			data[90277] <= 8'h10 ;
			data[90278] <= 8'h10 ;
			data[90279] <= 8'h10 ;
			data[90280] <= 8'h10 ;
			data[90281] <= 8'h10 ;
			data[90282] <= 8'h10 ;
			data[90283] <= 8'h10 ;
			data[90284] <= 8'h10 ;
			data[90285] <= 8'h10 ;
			data[90286] <= 8'h10 ;
			data[90287] <= 8'h10 ;
			data[90288] <= 8'h10 ;
			data[90289] <= 8'h10 ;
			data[90290] <= 8'h10 ;
			data[90291] <= 8'h10 ;
			data[90292] <= 8'h10 ;
			data[90293] <= 8'h10 ;
			data[90294] <= 8'h10 ;
			data[90295] <= 8'h10 ;
			data[90296] <= 8'h10 ;
			data[90297] <= 8'h10 ;
			data[90298] <= 8'h10 ;
			data[90299] <= 8'h10 ;
			data[90300] <= 8'h10 ;
			data[90301] <= 8'h10 ;
			data[90302] <= 8'h10 ;
			data[90303] <= 8'h10 ;
			data[90304] <= 8'h10 ;
			data[90305] <= 8'h10 ;
			data[90306] <= 8'h10 ;
			data[90307] <= 8'h10 ;
			data[90308] <= 8'h10 ;
			data[90309] <= 8'h10 ;
			data[90310] <= 8'h10 ;
			data[90311] <= 8'h10 ;
			data[90312] <= 8'h10 ;
			data[90313] <= 8'h10 ;
			data[90314] <= 8'h10 ;
			data[90315] <= 8'h10 ;
			data[90316] <= 8'h10 ;
			data[90317] <= 8'h10 ;
			data[90318] <= 8'h10 ;
			data[90319] <= 8'h10 ;
			data[90320] <= 8'h10 ;
			data[90321] <= 8'h10 ;
			data[90322] <= 8'h10 ;
			data[90323] <= 8'h10 ;
			data[90324] <= 8'h10 ;
			data[90325] <= 8'h10 ;
			data[90326] <= 8'h10 ;
			data[90327] <= 8'h10 ;
			data[90328] <= 8'h10 ;
			data[90329] <= 8'h10 ;
			data[90330] <= 8'h10 ;
			data[90331] <= 8'h10 ;
			data[90332] <= 8'h10 ;
			data[90333] <= 8'h10 ;
			data[90334] <= 8'h10 ;
			data[90335] <= 8'h10 ;
			data[90336] <= 8'h10 ;
			data[90337] <= 8'h10 ;
			data[90338] <= 8'h10 ;
			data[90339] <= 8'h10 ;
			data[90340] <= 8'h10 ;
			data[90341] <= 8'h10 ;
			data[90342] <= 8'h10 ;
			data[90343] <= 8'h10 ;
			data[90344] <= 8'h10 ;
			data[90345] <= 8'h10 ;
			data[90346] <= 8'h10 ;
			data[90347] <= 8'h10 ;
			data[90348] <= 8'h10 ;
			data[90349] <= 8'h10 ;
			data[90350] <= 8'h10 ;
			data[90351] <= 8'h10 ;
			data[90352] <= 8'h10 ;
			data[90353] <= 8'h10 ;
			data[90354] <= 8'h10 ;
			data[90355] <= 8'h10 ;
			data[90356] <= 8'h10 ;
			data[90357] <= 8'h10 ;
			data[90358] <= 8'h10 ;
			data[90359] <= 8'h10 ;
			data[90360] <= 8'h10 ;
			data[90361] <= 8'h10 ;
			data[90362] <= 8'h10 ;
			data[90363] <= 8'h10 ;
			data[90364] <= 8'h10 ;
			data[90365] <= 8'h10 ;
			data[90366] <= 8'h10 ;
			data[90367] <= 8'h10 ;
			data[90368] <= 8'h10 ;
			data[90369] <= 8'h10 ;
			data[90370] <= 8'h10 ;
			data[90371] <= 8'h10 ;
			data[90372] <= 8'h10 ;
			data[90373] <= 8'h10 ;
			data[90374] <= 8'h10 ;
			data[90375] <= 8'h10 ;
			data[90376] <= 8'h10 ;
			data[90377] <= 8'h10 ;
			data[90378] <= 8'h10 ;
			data[90379] <= 8'h10 ;
			data[90380] <= 8'h10 ;
			data[90381] <= 8'h10 ;
			data[90382] <= 8'h10 ;
			data[90383] <= 8'h10 ;
			data[90384] <= 8'h10 ;
			data[90385] <= 8'h10 ;
			data[90386] <= 8'h10 ;
			data[90387] <= 8'h10 ;
			data[90388] <= 8'h10 ;
			data[90389] <= 8'h10 ;
			data[90390] <= 8'h10 ;
			data[90391] <= 8'h10 ;
			data[90392] <= 8'h10 ;
			data[90393] <= 8'h10 ;
			data[90394] <= 8'h10 ;
			data[90395] <= 8'h10 ;
			data[90396] <= 8'h10 ;
			data[90397] <= 8'h10 ;
			data[90398] <= 8'h10 ;
			data[90399] <= 8'h10 ;
			data[90400] <= 8'h10 ;
			data[90401] <= 8'h10 ;
			data[90402] <= 8'h10 ;
			data[90403] <= 8'h10 ;
			data[90404] <= 8'h10 ;
			data[90405] <= 8'h10 ;
			data[90406] <= 8'h10 ;
			data[90407] <= 8'h10 ;
			data[90408] <= 8'h10 ;
			data[90409] <= 8'h10 ;
			data[90410] <= 8'h10 ;
			data[90411] <= 8'h10 ;
			data[90412] <= 8'h10 ;
			data[90413] <= 8'h10 ;
			data[90414] <= 8'h10 ;
			data[90415] <= 8'h10 ;
			data[90416] <= 8'h10 ;
			data[90417] <= 8'h10 ;
			data[90418] <= 8'h10 ;
			data[90419] <= 8'h10 ;
			data[90420] <= 8'h10 ;
			data[90421] <= 8'h10 ;
			data[90422] <= 8'h10 ;
			data[90423] <= 8'h10 ;
			data[90424] <= 8'h10 ;
			data[90425] <= 8'h10 ;
			data[90426] <= 8'h10 ;
			data[90427] <= 8'h10 ;
			data[90428] <= 8'h10 ;
			data[90429] <= 8'h10 ;
			data[90430] <= 8'h10 ;
			data[90431] <= 8'h10 ;
			data[90432] <= 8'h10 ;
			data[90433] <= 8'h10 ;
			data[90434] <= 8'h10 ;
			data[90435] <= 8'h10 ;
			data[90436] <= 8'h10 ;
			data[90437] <= 8'h10 ;
			data[90438] <= 8'h10 ;
			data[90439] <= 8'h10 ;
			data[90440] <= 8'h10 ;
			data[90441] <= 8'h10 ;
			data[90442] <= 8'h10 ;
			data[90443] <= 8'h10 ;
			data[90444] <= 8'h10 ;
			data[90445] <= 8'h10 ;
			data[90446] <= 8'h10 ;
			data[90447] <= 8'h10 ;
			data[90448] <= 8'h10 ;
			data[90449] <= 8'h10 ;
			data[90450] <= 8'h10 ;
			data[90451] <= 8'h10 ;
			data[90452] <= 8'h10 ;
			data[90453] <= 8'h10 ;
			data[90454] <= 8'h10 ;
			data[90455] <= 8'h10 ;
			data[90456] <= 8'h10 ;
			data[90457] <= 8'h10 ;
			data[90458] <= 8'h10 ;
			data[90459] <= 8'h10 ;
			data[90460] <= 8'h10 ;
			data[90461] <= 8'h10 ;
			data[90462] <= 8'h10 ;
			data[90463] <= 8'h10 ;
			data[90464] <= 8'h10 ;
			data[90465] <= 8'h10 ;
			data[90466] <= 8'h10 ;
			data[90467] <= 8'h10 ;
			data[90468] <= 8'h10 ;
			data[90469] <= 8'h10 ;
			data[90470] <= 8'h10 ;
			data[90471] <= 8'h10 ;
			data[90472] <= 8'h10 ;
			data[90473] <= 8'h10 ;
			data[90474] <= 8'h10 ;
			data[90475] <= 8'h10 ;
			data[90476] <= 8'h10 ;
			data[90477] <= 8'h10 ;
			data[90478] <= 8'h10 ;
			data[90479] <= 8'h10 ;
			data[90480] <= 8'h10 ;
			data[90481] <= 8'h10 ;
			data[90482] <= 8'h10 ;
			data[90483] <= 8'h10 ;
			data[90484] <= 8'h10 ;
			data[90485] <= 8'h10 ;
			data[90486] <= 8'h10 ;
			data[90487] <= 8'h10 ;
			data[90488] <= 8'h10 ;
			data[90489] <= 8'h10 ;
			data[90490] <= 8'h10 ;
			data[90491] <= 8'h10 ;
			data[90492] <= 8'h10 ;
			data[90493] <= 8'h10 ;
			data[90494] <= 8'h10 ;
			data[90495] <= 8'h10 ;
			data[90496] <= 8'h10 ;
			data[90497] <= 8'h10 ;
			data[90498] <= 8'h10 ;
			data[90499] <= 8'h10 ;
			data[90500] <= 8'h10 ;
			data[90501] <= 8'h10 ;
			data[90502] <= 8'h10 ;
			data[90503] <= 8'h10 ;
			data[90504] <= 8'h10 ;
			data[90505] <= 8'h10 ;
			data[90506] <= 8'h10 ;
			data[90507] <= 8'h10 ;
			data[90508] <= 8'h10 ;
			data[90509] <= 8'h10 ;
			data[90510] <= 8'h10 ;
			data[90511] <= 8'h10 ;
			data[90512] <= 8'h10 ;
			data[90513] <= 8'h10 ;
			data[90514] <= 8'h10 ;
			data[90515] <= 8'h10 ;
			data[90516] <= 8'h10 ;
			data[90517] <= 8'h10 ;
			data[90518] <= 8'h10 ;
			data[90519] <= 8'h10 ;
			data[90520] <= 8'h10 ;
			data[90521] <= 8'h10 ;
			data[90522] <= 8'h10 ;
			data[90523] <= 8'h10 ;
			data[90524] <= 8'h10 ;
			data[90525] <= 8'h10 ;
			data[90526] <= 8'h10 ;
			data[90527] <= 8'h10 ;
			data[90528] <= 8'h10 ;
			data[90529] <= 8'h10 ;
			data[90530] <= 8'h10 ;
			data[90531] <= 8'h10 ;
			data[90532] <= 8'h10 ;
			data[90533] <= 8'h10 ;
			data[90534] <= 8'h10 ;
			data[90535] <= 8'h10 ;
			data[90536] <= 8'h10 ;
			data[90537] <= 8'h10 ;
			data[90538] <= 8'h10 ;
			data[90539] <= 8'h10 ;
			data[90540] <= 8'h10 ;
			data[90541] <= 8'h10 ;
			data[90542] <= 8'h10 ;
			data[90543] <= 8'h10 ;
			data[90544] <= 8'h10 ;
			data[90545] <= 8'h10 ;
			data[90546] <= 8'h10 ;
			data[90547] <= 8'h10 ;
			data[90548] <= 8'h10 ;
			data[90549] <= 8'h10 ;
			data[90550] <= 8'h10 ;
			data[90551] <= 8'h10 ;
			data[90552] <= 8'h10 ;
			data[90553] <= 8'h10 ;
			data[90554] <= 8'h10 ;
			data[90555] <= 8'h10 ;
			data[90556] <= 8'h10 ;
			data[90557] <= 8'h10 ;
			data[90558] <= 8'h10 ;
			data[90559] <= 8'h10 ;
			data[90560] <= 8'h10 ;
			data[90561] <= 8'h10 ;
			data[90562] <= 8'h10 ;
			data[90563] <= 8'h10 ;
			data[90564] <= 8'h10 ;
			data[90565] <= 8'h10 ;
			data[90566] <= 8'h10 ;
			data[90567] <= 8'h10 ;
			data[90568] <= 8'h10 ;
			data[90569] <= 8'h10 ;
			data[90570] <= 8'h10 ;
			data[90571] <= 8'h10 ;
			data[90572] <= 8'h10 ;
			data[90573] <= 8'h10 ;
			data[90574] <= 8'h10 ;
			data[90575] <= 8'h10 ;
			data[90576] <= 8'h10 ;
			data[90577] <= 8'h10 ;
			data[90578] <= 8'h10 ;
			data[90579] <= 8'h10 ;
			data[90580] <= 8'h10 ;
			data[90581] <= 8'h10 ;
			data[90582] <= 8'h10 ;
			data[90583] <= 8'h10 ;
			data[90584] <= 8'h10 ;
			data[90585] <= 8'h10 ;
			data[90586] <= 8'h10 ;
			data[90587] <= 8'h10 ;
			data[90588] <= 8'h10 ;
			data[90589] <= 8'h10 ;
			data[90590] <= 8'h10 ;
			data[90591] <= 8'h10 ;
			data[90592] <= 8'h10 ;
			data[90593] <= 8'h10 ;
			data[90594] <= 8'h10 ;
			data[90595] <= 8'h10 ;
			data[90596] <= 8'h10 ;
			data[90597] <= 8'h10 ;
			data[90598] <= 8'h10 ;
			data[90599] <= 8'h10 ;
			data[90600] <= 8'h10 ;
			data[90601] <= 8'h10 ;
			data[90602] <= 8'h10 ;
			data[90603] <= 8'h10 ;
			data[90604] <= 8'h10 ;
			data[90605] <= 8'h10 ;
			data[90606] <= 8'h10 ;
			data[90607] <= 8'h10 ;
			data[90608] <= 8'h10 ;
			data[90609] <= 8'h10 ;
			data[90610] <= 8'h10 ;
			data[90611] <= 8'h10 ;
			data[90612] <= 8'h10 ;
			data[90613] <= 8'h10 ;
			data[90614] <= 8'h10 ;
			data[90615] <= 8'h10 ;
			data[90616] <= 8'h10 ;
			data[90617] <= 8'h10 ;
			data[90618] <= 8'h10 ;
			data[90619] <= 8'h10 ;
			data[90620] <= 8'h10 ;
			data[90621] <= 8'h10 ;
			data[90622] <= 8'h10 ;
			data[90623] <= 8'h10 ;
			data[90624] <= 8'h10 ;
			data[90625] <= 8'h10 ;
			data[90626] <= 8'h10 ;
			data[90627] <= 8'h10 ;
			data[90628] <= 8'h10 ;
			data[90629] <= 8'h10 ;
			data[90630] <= 8'h10 ;
			data[90631] <= 8'h10 ;
			data[90632] <= 8'h10 ;
			data[90633] <= 8'h10 ;
			data[90634] <= 8'h10 ;
			data[90635] <= 8'h10 ;
			data[90636] <= 8'h10 ;
			data[90637] <= 8'h10 ;
			data[90638] <= 8'h10 ;
			data[90639] <= 8'h10 ;
			data[90640] <= 8'h10 ;
			data[90641] <= 8'h10 ;
			data[90642] <= 8'h10 ;
			data[90643] <= 8'h10 ;
			data[90644] <= 8'h10 ;
			data[90645] <= 8'h10 ;
			data[90646] <= 8'h10 ;
			data[90647] <= 8'h10 ;
			data[90648] <= 8'h10 ;
			data[90649] <= 8'h10 ;
			data[90650] <= 8'h10 ;
			data[90651] <= 8'h10 ;
			data[90652] <= 8'h10 ;
			data[90653] <= 8'h10 ;
			data[90654] <= 8'h10 ;
			data[90655] <= 8'h10 ;
			data[90656] <= 8'h10 ;
			data[90657] <= 8'h10 ;
			data[90658] <= 8'h10 ;
			data[90659] <= 8'h10 ;
			data[90660] <= 8'h10 ;
			data[90661] <= 8'h10 ;
			data[90662] <= 8'h10 ;
			data[90663] <= 8'h10 ;
			data[90664] <= 8'h10 ;
			data[90665] <= 8'h10 ;
			data[90666] <= 8'h10 ;
			data[90667] <= 8'h10 ;
			data[90668] <= 8'h10 ;
			data[90669] <= 8'h10 ;
			data[90670] <= 8'h10 ;
			data[90671] <= 8'h10 ;
			data[90672] <= 8'h10 ;
			data[90673] <= 8'h10 ;
			data[90674] <= 8'h10 ;
			data[90675] <= 8'h10 ;
			data[90676] <= 8'h10 ;
			data[90677] <= 8'h10 ;
			data[90678] <= 8'h10 ;
			data[90679] <= 8'h10 ;
			data[90680] <= 8'h10 ;
			data[90681] <= 8'h10 ;
			data[90682] <= 8'h10 ;
			data[90683] <= 8'h10 ;
			data[90684] <= 8'h10 ;
			data[90685] <= 8'h10 ;
			data[90686] <= 8'h10 ;
			data[90687] <= 8'h10 ;
			data[90688] <= 8'h10 ;
			data[90689] <= 8'h10 ;
			data[90690] <= 8'h10 ;
			data[90691] <= 8'h10 ;
			data[90692] <= 8'h10 ;
			data[90693] <= 8'h10 ;
			data[90694] <= 8'h10 ;
			data[90695] <= 8'h10 ;
			data[90696] <= 8'h10 ;
			data[90697] <= 8'h10 ;
			data[90698] <= 8'h10 ;
			data[90699] <= 8'h10 ;
			data[90700] <= 8'h10 ;
			data[90701] <= 8'h10 ;
			data[90702] <= 8'h10 ;
			data[90703] <= 8'h10 ;
			data[90704] <= 8'h10 ;
			data[90705] <= 8'h10 ;
			data[90706] <= 8'h10 ;
			data[90707] <= 8'h10 ;
			data[90708] <= 8'h10 ;
			data[90709] <= 8'h10 ;
			data[90710] <= 8'h10 ;
			data[90711] <= 8'h10 ;
			data[90712] <= 8'h10 ;
			data[90713] <= 8'h10 ;
			data[90714] <= 8'h10 ;
			data[90715] <= 8'h10 ;
			data[90716] <= 8'h10 ;
			data[90717] <= 8'h10 ;
			data[90718] <= 8'h10 ;
			data[90719] <= 8'h10 ;
			data[90720] <= 8'h10 ;
			data[90721] <= 8'h10 ;
			data[90722] <= 8'h10 ;
			data[90723] <= 8'h10 ;
			data[90724] <= 8'h10 ;
			data[90725] <= 8'h10 ;
			data[90726] <= 8'h10 ;
			data[90727] <= 8'h10 ;
			data[90728] <= 8'h10 ;
			data[90729] <= 8'h10 ;
			data[90730] <= 8'h10 ;
			data[90731] <= 8'h10 ;
			data[90732] <= 8'h10 ;
			data[90733] <= 8'h10 ;
			data[90734] <= 8'h10 ;
			data[90735] <= 8'h10 ;
			data[90736] <= 8'h10 ;
			data[90737] <= 8'h10 ;
			data[90738] <= 8'h10 ;
			data[90739] <= 8'h10 ;
			data[90740] <= 8'h10 ;
			data[90741] <= 8'h10 ;
			data[90742] <= 8'h10 ;
			data[90743] <= 8'h10 ;
			data[90744] <= 8'h10 ;
			data[90745] <= 8'h10 ;
			data[90746] <= 8'h10 ;
			data[90747] <= 8'h10 ;
			data[90748] <= 8'h10 ;
			data[90749] <= 8'h10 ;
			data[90750] <= 8'h10 ;
			data[90751] <= 8'h10 ;
			data[90752] <= 8'h10 ;
			data[90753] <= 8'h10 ;
			data[90754] <= 8'h10 ;
			data[90755] <= 8'h10 ;
			data[90756] <= 8'h10 ;
			data[90757] <= 8'h10 ;
			data[90758] <= 8'h10 ;
			data[90759] <= 8'h10 ;
			data[90760] <= 8'h10 ;
			data[90761] <= 8'h10 ;
			data[90762] <= 8'h10 ;
			data[90763] <= 8'h10 ;
			data[90764] <= 8'h10 ;
			data[90765] <= 8'h10 ;
			data[90766] <= 8'h10 ;
			data[90767] <= 8'h10 ;
			data[90768] <= 8'h10 ;
			data[90769] <= 8'h10 ;
			data[90770] <= 8'h10 ;
			data[90771] <= 8'h10 ;
			data[90772] <= 8'h10 ;
			data[90773] <= 8'h10 ;
			data[90774] <= 8'h10 ;
			data[90775] <= 8'h10 ;
			data[90776] <= 8'h10 ;
			data[90777] <= 8'h10 ;
			data[90778] <= 8'h10 ;
			data[90779] <= 8'h10 ;
			data[90780] <= 8'h10 ;
			data[90781] <= 8'h10 ;
			data[90782] <= 8'h10 ;
			data[90783] <= 8'h10 ;
			data[90784] <= 8'h10 ;
			data[90785] <= 8'h10 ;
			data[90786] <= 8'h10 ;
			data[90787] <= 8'h10 ;
			data[90788] <= 8'h10 ;
			data[90789] <= 8'h10 ;
			data[90790] <= 8'h10 ;
			data[90791] <= 8'h10 ;
			data[90792] <= 8'h10 ;
			data[90793] <= 8'h10 ;
			data[90794] <= 8'h10 ;
			data[90795] <= 8'h10 ;
			data[90796] <= 8'h10 ;
			data[90797] <= 8'h10 ;
			data[90798] <= 8'h10 ;
			data[90799] <= 8'h10 ;
			data[90800] <= 8'h10 ;
			data[90801] <= 8'h10 ;
			data[90802] <= 8'h10 ;
			data[90803] <= 8'h10 ;
			data[90804] <= 8'h10 ;
			data[90805] <= 8'h10 ;
			data[90806] <= 8'h10 ;
			data[90807] <= 8'h10 ;
			data[90808] <= 8'h10 ;
			data[90809] <= 8'h10 ;
			data[90810] <= 8'h10 ;
			data[90811] <= 8'h10 ;
			data[90812] <= 8'h10 ;
			data[90813] <= 8'h10 ;
			data[90814] <= 8'h10 ;
			data[90815] <= 8'h10 ;
			data[90816] <= 8'h10 ;
			data[90817] <= 8'h10 ;
			data[90818] <= 8'h10 ;
			data[90819] <= 8'h10 ;
			data[90820] <= 8'h10 ;
			data[90821] <= 8'h10 ;
			data[90822] <= 8'h10 ;
			data[90823] <= 8'h10 ;
			data[90824] <= 8'h10 ;
			data[90825] <= 8'h10 ;
			data[90826] <= 8'h10 ;
			data[90827] <= 8'h10 ;
			data[90828] <= 8'h10 ;
			data[90829] <= 8'h10 ;
			data[90830] <= 8'h10 ;
			data[90831] <= 8'h10 ;
			data[90832] <= 8'h10 ;
			data[90833] <= 8'h10 ;
			data[90834] <= 8'h10 ;
			data[90835] <= 8'h10 ;
			data[90836] <= 8'h10 ;
			data[90837] <= 8'h10 ;
			data[90838] <= 8'h10 ;
			data[90839] <= 8'h10 ;
			data[90840] <= 8'h10 ;
			data[90841] <= 8'h10 ;
			data[90842] <= 8'h10 ;
			data[90843] <= 8'h10 ;
			data[90844] <= 8'h10 ;
			data[90845] <= 8'h10 ;
			data[90846] <= 8'h10 ;
			data[90847] <= 8'h10 ;
			data[90848] <= 8'h10 ;
			data[90849] <= 8'h10 ;
			data[90850] <= 8'h10 ;
			data[90851] <= 8'h10 ;
			data[90852] <= 8'h10 ;
			data[90853] <= 8'h10 ;
			data[90854] <= 8'h10 ;
			data[90855] <= 8'h10 ;
			data[90856] <= 8'h10 ;
			data[90857] <= 8'h10 ;
			data[90858] <= 8'h10 ;
			data[90859] <= 8'h10 ;
			data[90860] <= 8'h10 ;
			data[90861] <= 8'h10 ;
			data[90862] <= 8'h10 ;
			data[90863] <= 8'h10 ;
			data[90864] <= 8'h10 ;
			data[90865] <= 8'h10 ;
			data[90866] <= 8'h10 ;
			data[90867] <= 8'h10 ;
			data[90868] <= 8'h10 ;
			data[90869] <= 8'h10 ;
			data[90870] <= 8'h10 ;
			data[90871] <= 8'h10 ;
			data[90872] <= 8'h10 ;
			data[90873] <= 8'h10 ;
			data[90874] <= 8'h10 ;
			data[90875] <= 8'h10 ;
			data[90876] <= 8'h10 ;
			data[90877] <= 8'h10 ;
			data[90878] <= 8'h10 ;
			data[90879] <= 8'h10 ;
			data[90880] <= 8'h10 ;
			data[90881] <= 8'h10 ;
			data[90882] <= 8'h10 ;
			data[90883] <= 8'h10 ;
			data[90884] <= 8'h10 ;
			data[90885] <= 8'h10 ;
			data[90886] <= 8'h10 ;
			data[90887] <= 8'h10 ;
			data[90888] <= 8'h10 ;
			data[90889] <= 8'h10 ;
			data[90890] <= 8'h10 ;
			data[90891] <= 8'h10 ;
			data[90892] <= 8'h10 ;
			data[90893] <= 8'h10 ;
			data[90894] <= 8'h10 ;
			data[90895] <= 8'h10 ;
			data[90896] <= 8'h10 ;
			data[90897] <= 8'h10 ;
			data[90898] <= 8'h10 ;
			data[90899] <= 8'h10 ;
			data[90900] <= 8'h10 ;
			data[90901] <= 8'h10 ;
			data[90902] <= 8'h10 ;
			data[90903] <= 8'h10 ;
			data[90904] <= 8'h10 ;
			data[90905] <= 8'h10 ;
			data[90906] <= 8'h10 ;
			data[90907] <= 8'h10 ;
			data[90908] <= 8'h10 ;
			data[90909] <= 8'h10 ;
			data[90910] <= 8'h10 ;
			data[90911] <= 8'h10 ;
			data[90912] <= 8'h10 ;
			data[90913] <= 8'h10 ;
			data[90914] <= 8'h10 ;
			data[90915] <= 8'h10 ;
			data[90916] <= 8'h10 ;
			data[90917] <= 8'h10 ;
			data[90918] <= 8'h10 ;
			data[90919] <= 8'h10 ;
			data[90920] <= 8'h10 ;
			data[90921] <= 8'h10 ;
			data[90922] <= 8'h10 ;
			data[90923] <= 8'h10 ;
			data[90924] <= 8'h10 ;
			data[90925] <= 8'h10 ;
			data[90926] <= 8'h10 ;
			data[90927] <= 8'h10 ;
			data[90928] <= 8'h10 ;
			data[90929] <= 8'h10 ;
			data[90930] <= 8'h10 ;
			data[90931] <= 8'h10 ;
			data[90932] <= 8'h10 ;
			data[90933] <= 8'h10 ;
			data[90934] <= 8'h10 ;
			data[90935] <= 8'h10 ;
			data[90936] <= 8'h10 ;
			data[90937] <= 8'h10 ;
			data[90938] <= 8'h10 ;
			data[90939] <= 8'h10 ;
			data[90940] <= 8'h10 ;
			data[90941] <= 8'h10 ;
			data[90942] <= 8'h10 ;
			data[90943] <= 8'h10 ;
			data[90944] <= 8'h10 ;
			data[90945] <= 8'h10 ;
			data[90946] <= 8'h10 ;
			data[90947] <= 8'h10 ;
			data[90948] <= 8'h10 ;
			data[90949] <= 8'h10 ;
			data[90950] <= 8'h10 ;
			data[90951] <= 8'h10 ;
			data[90952] <= 8'h10 ;
			data[90953] <= 8'h10 ;
			data[90954] <= 8'h10 ;
			data[90955] <= 8'h10 ;
			data[90956] <= 8'h10 ;
			data[90957] <= 8'h10 ;
			data[90958] <= 8'h10 ;
			data[90959] <= 8'h10 ;
			data[90960] <= 8'h10 ;
			data[90961] <= 8'h10 ;
			data[90962] <= 8'h10 ;
			data[90963] <= 8'h10 ;
			data[90964] <= 8'h10 ;
			data[90965] <= 8'h10 ;
			data[90966] <= 8'h10 ;
			data[90967] <= 8'h10 ;
			data[90968] <= 8'h10 ;
			data[90969] <= 8'h10 ;
			data[90970] <= 8'h10 ;
			data[90971] <= 8'h10 ;
			data[90972] <= 8'h10 ;
			data[90973] <= 8'h10 ;
			data[90974] <= 8'h10 ;
			data[90975] <= 8'h10 ;
			data[90976] <= 8'h10 ;
			data[90977] <= 8'h10 ;
			data[90978] <= 8'h10 ;
			data[90979] <= 8'h10 ;
			data[90980] <= 8'h10 ;
			data[90981] <= 8'h10 ;
			data[90982] <= 8'h10 ;
			data[90983] <= 8'h10 ;
			data[90984] <= 8'h10 ;
			data[90985] <= 8'h10 ;
			data[90986] <= 8'h10 ;
			data[90987] <= 8'h10 ;
			data[90988] <= 8'h10 ;
			data[90989] <= 8'h10 ;
			data[90990] <= 8'h10 ;
			data[90991] <= 8'h10 ;
			data[90992] <= 8'h10 ;
			data[90993] <= 8'h10 ;
			data[90994] <= 8'h10 ;
			data[90995] <= 8'h10 ;
			data[90996] <= 8'h10 ;
			data[90997] <= 8'h10 ;
			data[90998] <= 8'h10 ;
			data[90999] <= 8'h10 ;
			data[91000] <= 8'h10 ;
			data[91001] <= 8'h10 ;
			data[91002] <= 8'h10 ;
			data[91003] <= 8'h10 ;
			data[91004] <= 8'h10 ;
			data[91005] <= 8'h10 ;
			data[91006] <= 8'h10 ;
			data[91007] <= 8'h10 ;
			data[91008] <= 8'h10 ;
			data[91009] <= 8'h10 ;
			data[91010] <= 8'h10 ;
			data[91011] <= 8'h10 ;
			data[91012] <= 8'h10 ;
			data[91013] <= 8'h10 ;
			data[91014] <= 8'h10 ;
			data[91015] <= 8'h10 ;
			data[91016] <= 8'h10 ;
			data[91017] <= 8'h10 ;
			data[91018] <= 8'h10 ;
			data[91019] <= 8'h10 ;
			data[91020] <= 8'h10 ;
			data[91021] <= 8'h10 ;
			data[91022] <= 8'h10 ;
			data[91023] <= 8'h10 ;
			data[91024] <= 8'h10 ;
			data[91025] <= 8'h10 ;
			data[91026] <= 8'h10 ;
			data[91027] <= 8'h10 ;
			data[91028] <= 8'h10 ;
			data[91029] <= 8'h10 ;
			data[91030] <= 8'h10 ;
			data[91031] <= 8'h10 ;
			data[91032] <= 8'h10 ;
			data[91033] <= 8'h10 ;
			data[91034] <= 8'h10 ;
			data[91035] <= 8'h10 ;
			data[91036] <= 8'h10 ;
			data[91037] <= 8'h10 ;
			data[91038] <= 8'h10 ;
			data[91039] <= 8'h10 ;
			data[91040] <= 8'h10 ;
			data[91041] <= 8'h10 ;
			data[91042] <= 8'h10 ;
			data[91043] <= 8'h10 ;
			data[91044] <= 8'h10 ;
			data[91045] <= 8'h10 ;
			data[91046] <= 8'h10 ;
			data[91047] <= 8'h10 ;
			data[91048] <= 8'h10 ;
			data[91049] <= 8'h10 ;
			data[91050] <= 8'h10 ;
			data[91051] <= 8'h10 ;
			data[91052] <= 8'h10 ;
			data[91053] <= 8'h10 ;
			data[91054] <= 8'h10 ;
			data[91055] <= 8'h10 ;
			data[91056] <= 8'h10 ;
			data[91057] <= 8'h10 ;
			data[91058] <= 8'h10 ;
			data[91059] <= 8'h10 ;
			data[91060] <= 8'h10 ;
			data[91061] <= 8'h10 ;
			data[91062] <= 8'h10 ;
			data[91063] <= 8'h10 ;
			data[91064] <= 8'h10 ;
			data[91065] <= 8'h10 ;
			data[91066] <= 8'h10 ;
			data[91067] <= 8'h10 ;
			data[91068] <= 8'h10 ;
			data[91069] <= 8'h10 ;
			data[91070] <= 8'h10 ;
			data[91071] <= 8'h10 ;
			data[91072] <= 8'h10 ;
			data[91073] <= 8'h10 ;
			data[91074] <= 8'h10 ;
			data[91075] <= 8'h10 ;
			data[91076] <= 8'h10 ;
			data[91077] <= 8'h10 ;
			data[91078] <= 8'h10 ;
			data[91079] <= 8'h10 ;
			data[91080] <= 8'h10 ;
			data[91081] <= 8'h10 ;
			data[91082] <= 8'h10 ;
			data[91083] <= 8'h10 ;
			data[91084] <= 8'h10 ;
			data[91085] <= 8'h10 ;
			data[91086] <= 8'h10 ;
			data[91087] <= 8'h10 ;
			data[91088] <= 8'h10 ;
			data[91089] <= 8'h10 ;
			data[91090] <= 8'h10 ;
			data[91091] <= 8'h10 ;
			data[91092] <= 8'h10 ;
			data[91093] <= 8'h10 ;
			data[91094] <= 8'h10 ;
			data[91095] <= 8'h10 ;
			data[91096] <= 8'h10 ;
			data[91097] <= 8'h10 ;
			data[91098] <= 8'h10 ;
			data[91099] <= 8'h10 ;
			data[91100] <= 8'h10 ;
			data[91101] <= 8'h10 ;
			data[91102] <= 8'h10 ;
			data[91103] <= 8'h10 ;
			data[91104] <= 8'h10 ;
			data[91105] <= 8'h10 ;
			data[91106] <= 8'h10 ;
			data[91107] <= 8'h10 ;
			data[91108] <= 8'h10 ;
			data[91109] <= 8'h10 ;
			data[91110] <= 8'h10 ;
			data[91111] <= 8'h10 ;
			data[91112] <= 8'h10 ;
			data[91113] <= 8'h10 ;
			data[91114] <= 8'h10 ;
			data[91115] <= 8'h10 ;
			data[91116] <= 8'h10 ;
			data[91117] <= 8'h10 ;
			data[91118] <= 8'h10 ;
			data[91119] <= 8'h10 ;
			data[91120] <= 8'h10 ;
			data[91121] <= 8'h10 ;
			data[91122] <= 8'h10 ;
			data[91123] <= 8'h10 ;
			data[91124] <= 8'h10 ;
			data[91125] <= 8'h10 ;
			data[91126] <= 8'h10 ;
			data[91127] <= 8'h10 ;
			data[91128] <= 8'h10 ;
			data[91129] <= 8'h10 ;
			data[91130] <= 8'h10 ;
			data[91131] <= 8'h10 ;
			data[91132] <= 8'h10 ;
			data[91133] <= 8'h10 ;
			data[91134] <= 8'h10 ;
			data[91135] <= 8'h10 ;
			data[91136] <= 8'h10 ;
			data[91137] <= 8'h10 ;
			data[91138] <= 8'h10 ;
			data[91139] <= 8'h10 ;
			data[91140] <= 8'h10 ;
			data[91141] <= 8'h10 ;
			data[91142] <= 8'h10 ;
			data[91143] <= 8'h10 ;
			data[91144] <= 8'h10 ;
			data[91145] <= 8'h10 ;
			data[91146] <= 8'h10 ;
			data[91147] <= 8'h10 ;
			data[91148] <= 8'h10 ;
			data[91149] <= 8'h10 ;
			data[91150] <= 8'h10 ;
			data[91151] <= 8'h10 ;
			data[91152] <= 8'h10 ;
			data[91153] <= 8'h10 ;
			data[91154] <= 8'h10 ;
			data[91155] <= 8'h10 ;
			data[91156] <= 8'h10 ;
			data[91157] <= 8'h10 ;
			data[91158] <= 8'h10 ;
			data[91159] <= 8'h10 ;
			data[91160] <= 8'h10 ;
			data[91161] <= 8'h10 ;
			data[91162] <= 8'h10 ;
			data[91163] <= 8'h10 ;
			data[91164] <= 8'h10 ;
			data[91165] <= 8'h10 ;
			data[91166] <= 8'h10 ;
			data[91167] <= 8'h10 ;
			data[91168] <= 8'h10 ;
			data[91169] <= 8'h10 ;
			data[91170] <= 8'h10 ;
			data[91171] <= 8'h10 ;
			data[91172] <= 8'h10 ;
			data[91173] <= 8'h10 ;
			data[91174] <= 8'h10 ;
			data[91175] <= 8'h10 ;
			data[91176] <= 8'h10 ;
			data[91177] <= 8'h10 ;
			data[91178] <= 8'h10 ;
			data[91179] <= 8'h10 ;
			data[91180] <= 8'h10 ;
			data[91181] <= 8'h10 ;
			data[91182] <= 8'h10 ;
			data[91183] <= 8'h10 ;
			data[91184] <= 8'h10 ;
			data[91185] <= 8'h10 ;
			data[91186] <= 8'h10 ;
			data[91187] <= 8'h10 ;
			data[91188] <= 8'h10 ;
			data[91189] <= 8'h10 ;
			data[91190] <= 8'h10 ;
			data[91191] <= 8'h10 ;
			data[91192] <= 8'h10 ;
			data[91193] <= 8'h10 ;
			data[91194] <= 8'h10 ;
			data[91195] <= 8'h10 ;
			data[91196] <= 8'h10 ;
			data[91197] <= 8'h10 ;
			data[91198] <= 8'h10 ;
			data[91199] <= 8'h10 ;
			data[91200] <= 8'h10 ;
			data[91201] <= 8'h10 ;
			data[91202] <= 8'h10 ;
			data[91203] <= 8'h10 ;
			data[91204] <= 8'h10 ;
			data[91205] <= 8'h10 ;
			data[91206] <= 8'h10 ;
			data[91207] <= 8'h10 ;
			data[91208] <= 8'h10 ;
			data[91209] <= 8'h10 ;
			data[91210] <= 8'h10 ;
			data[91211] <= 8'h10 ;
			data[91212] <= 8'h10 ;
			data[91213] <= 8'h10 ;
			data[91214] <= 8'h10 ;
			data[91215] <= 8'h10 ;
			data[91216] <= 8'h10 ;
			data[91217] <= 8'h10 ;
			data[91218] <= 8'h10 ;
			data[91219] <= 8'h10 ;
			data[91220] <= 8'h10 ;
			data[91221] <= 8'h10 ;
			data[91222] <= 8'h10 ;
			data[91223] <= 8'h10 ;
			data[91224] <= 8'h10 ;
			data[91225] <= 8'h10 ;
			data[91226] <= 8'h10 ;
			data[91227] <= 8'h10 ;
			data[91228] <= 8'h10 ;
			data[91229] <= 8'h10 ;
			data[91230] <= 8'h10 ;
			data[91231] <= 8'h10 ;
			data[91232] <= 8'h10 ;
			data[91233] <= 8'h10 ;
			data[91234] <= 8'h10 ;
			data[91235] <= 8'h10 ;
			data[91236] <= 8'h10 ;
			data[91237] <= 8'h10 ;
			data[91238] <= 8'h10 ;
			data[91239] <= 8'h10 ;
			data[91240] <= 8'h10 ;
			data[91241] <= 8'h10 ;
			data[91242] <= 8'h10 ;
			data[91243] <= 8'h10 ;
			data[91244] <= 8'h10 ;
			data[91245] <= 8'h10 ;
			data[91246] <= 8'h10 ;
			data[91247] <= 8'h10 ;
			data[91248] <= 8'h10 ;
			data[91249] <= 8'h10 ;
			data[91250] <= 8'h10 ;
			data[91251] <= 8'h10 ;
			data[91252] <= 8'h10 ;
			data[91253] <= 8'h10 ;
			data[91254] <= 8'h10 ;
			data[91255] <= 8'h10 ;
			data[91256] <= 8'h10 ;
			data[91257] <= 8'h10 ;
			data[91258] <= 8'h10 ;
			data[91259] <= 8'h10 ;
			data[91260] <= 8'h10 ;
			data[91261] <= 8'h10 ;
			data[91262] <= 8'h10 ;
			data[91263] <= 8'h10 ;
			data[91264] <= 8'h10 ;
			data[91265] <= 8'h10 ;
			data[91266] <= 8'h10 ;
			data[91267] <= 8'h10 ;
			data[91268] <= 8'h10 ;
			data[91269] <= 8'h10 ;
			data[91270] <= 8'h10 ;
			data[91271] <= 8'h10 ;
			data[91272] <= 8'h10 ;
			data[91273] <= 8'h10 ;
			data[91274] <= 8'h10 ;
			data[91275] <= 8'h10 ;
			data[91276] <= 8'h10 ;
			data[91277] <= 8'h10 ;
			data[91278] <= 8'h10 ;
			data[91279] <= 8'h10 ;
			data[91280] <= 8'h10 ;
			data[91281] <= 8'h10 ;
			data[91282] <= 8'h10 ;
			data[91283] <= 8'h10 ;
			data[91284] <= 8'h10 ;
			data[91285] <= 8'h10 ;
			data[91286] <= 8'h10 ;
			data[91287] <= 8'h10 ;
			data[91288] <= 8'h10 ;
			data[91289] <= 8'h10 ;
			data[91290] <= 8'h10 ;
			data[91291] <= 8'h10 ;
			data[91292] <= 8'h10 ;
			data[91293] <= 8'h10 ;
			data[91294] <= 8'h10 ;
			data[91295] <= 8'h10 ;
			data[91296] <= 8'h10 ;
			data[91297] <= 8'h10 ;
			data[91298] <= 8'h10 ;
			data[91299] <= 8'h10 ;
			data[91300] <= 8'h10 ;
			data[91301] <= 8'h10 ;
			data[91302] <= 8'h10 ;
			data[91303] <= 8'h10 ;
			data[91304] <= 8'h10 ;
			data[91305] <= 8'h10 ;
			data[91306] <= 8'h10 ;
			data[91307] <= 8'h10 ;
			data[91308] <= 8'h10 ;
			data[91309] <= 8'h10 ;
			data[91310] <= 8'h10 ;
			data[91311] <= 8'h10 ;
			data[91312] <= 8'h10 ;
			data[91313] <= 8'h10 ;
			data[91314] <= 8'h10 ;
			data[91315] <= 8'h10 ;
			data[91316] <= 8'h10 ;
			data[91317] <= 8'h10 ;
			data[91318] <= 8'h10 ;
			data[91319] <= 8'h10 ;
			data[91320] <= 8'h10 ;
			data[91321] <= 8'h10 ;
			data[91322] <= 8'h10 ;
			data[91323] <= 8'h10 ;
			data[91324] <= 8'h10 ;
			data[91325] <= 8'h10 ;
			data[91326] <= 8'h10 ;
			data[91327] <= 8'h10 ;
			data[91328] <= 8'h10 ;
			data[91329] <= 8'h10 ;
			data[91330] <= 8'h10 ;
			data[91331] <= 8'h10 ;
			data[91332] <= 8'h10 ;
			data[91333] <= 8'h10 ;
			data[91334] <= 8'h10 ;
			data[91335] <= 8'h10 ;
			data[91336] <= 8'h10 ;
			data[91337] <= 8'h10 ;
			data[91338] <= 8'h10 ;
			data[91339] <= 8'h10 ;
			data[91340] <= 8'h10 ;
			data[91341] <= 8'h10 ;
			data[91342] <= 8'h10 ;
			data[91343] <= 8'h10 ;
			data[91344] <= 8'h10 ;
			data[91345] <= 8'h10 ;
			data[91346] <= 8'h10 ;
			data[91347] <= 8'h10 ;
			data[91348] <= 8'h10 ;
			data[91349] <= 8'h10 ;
			data[91350] <= 8'h10 ;
			data[91351] <= 8'h10 ;
			data[91352] <= 8'h10 ;
			data[91353] <= 8'h10 ;
			data[91354] <= 8'h10 ;
			data[91355] <= 8'h10 ;
			data[91356] <= 8'h10 ;
			data[91357] <= 8'h10 ;
			data[91358] <= 8'h10 ;
			data[91359] <= 8'h10 ;
			data[91360] <= 8'h10 ;
			data[91361] <= 8'h10 ;
			data[91362] <= 8'h10 ;
			data[91363] <= 8'h10 ;
			data[91364] <= 8'h10 ;
			data[91365] <= 8'h10 ;
			data[91366] <= 8'h10 ;
			data[91367] <= 8'h10 ;
			data[91368] <= 8'h10 ;
			data[91369] <= 8'h10 ;
			data[91370] <= 8'h10 ;
			data[91371] <= 8'h10 ;
			data[91372] <= 8'h10 ;
			data[91373] <= 8'h10 ;
			data[91374] <= 8'h10 ;
			data[91375] <= 8'h10 ;
			data[91376] <= 8'h10 ;
			data[91377] <= 8'h10 ;
			data[91378] <= 8'h10 ;
			data[91379] <= 8'h10 ;
			data[91380] <= 8'h10 ;
			data[91381] <= 8'h10 ;
			data[91382] <= 8'h10 ;
			data[91383] <= 8'h10 ;
			data[91384] <= 8'h10 ;
			data[91385] <= 8'h10 ;
			data[91386] <= 8'h10 ;
			data[91387] <= 8'h10 ;
			data[91388] <= 8'h10 ;
			data[91389] <= 8'h10 ;
			data[91390] <= 8'h10 ;
			data[91391] <= 8'h10 ;
			data[91392] <= 8'h10 ;
			data[91393] <= 8'h10 ;
			data[91394] <= 8'h10 ;
			data[91395] <= 8'h10 ;
			data[91396] <= 8'h10 ;
			data[91397] <= 8'h10 ;
			data[91398] <= 8'h10 ;
			data[91399] <= 8'h10 ;
			data[91400] <= 8'h10 ;
			data[91401] <= 8'h10 ;
			data[91402] <= 8'h10 ;
			data[91403] <= 8'h10 ;
			data[91404] <= 8'h10 ;
			data[91405] <= 8'h10 ;
			data[91406] <= 8'h10 ;
			data[91407] <= 8'h10 ;
			data[91408] <= 8'h10 ;
			data[91409] <= 8'h10 ;
			data[91410] <= 8'h10 ;
			data[91411] <= 8'h10 ;
			data[91412] <= 8'h10 ;
			data[91413] <= 8'h10 ;
			data[91414] <= 8'h10 ;
			data[91415] <= 8'h10 ;
			data[91416] <= 8'h10 ;
			data[91417] <= 8'h10 ;
			data[91418] <= 8'h10 ;
			data[91419] <= 8'h10 ;
			data[91420] <= 8'h10 ;
			data[91421] <= 8'h10 ;
			data[91422] <= 8'h10 ;
			data[91423] <= 8'h10 ;
			data[91424] <= 8'h10 ;
			data[91425] <= 8'h10 ;
			data[91426] <= 8'h10 ;
			data[91427] <= 8'h10 ;
			data[91428] <= 8'h10 ;
			data[91429] <= 8'h10 ;
			data[91430] <= 8'h10 ;
			data[91431] <= 8'h10 ;
			data[91432] <= 8'h10 ;
			data[91433] <= 8'h10 ;
			data[91434] <= 8'h10 ;
			data[91435] <= 8'h10 ;
			data[91436] <= 8'h10 ;
			data[91437] <= 8'h10 ;
			data[91438] <= 8'h10 ;
			data[91439] <= 8'h10 ;
			data[91440] <= 8'h10 ;
			data[91441] <= 8'h10 ;
			data[91442] <= 8'h10 ;
			data[91443] <= 8'h10 ;
			data[91444] <= 8'h10 ;
			data[91445] <= 8'h10 ;
			data[91446] <= 8'h10 ;
			data[91447] <= 8'h10 ;
			data[91448] <= 8'h10 ;
			data[91449] <= 8'h10 ;
			data[91450] <= 8'h10 ;
			data[91451] <= 8'h10 ;
			data[91452] <= 8'h10 ;
			data[91453] <= 8'h10 ;
			data[91454] <= 8'h10 ;
			data[91455] <= 8'h10 ;
			data[91456] <= 8'h10 ;
			data[91457] <= 8'h10 ;
			data[91458] <= 8'h10 ;
			data[91459] <= 8'h10 ;
			data[91460] <= 8'h10 ;
			data[91461] <= 8'h10 ;
			data[91462] <= 8'h10 ;
			data[91463] <= 8'h10 ;
			data[91464] <= 8'h10 ;
			data[91465] <= 8'h10 ;
			data[91466] <= 8'h10 ;
			data[91467] <= 8'h10 ;
			data[91468] <= 8'h10 ;
			data[91469] <= 8'h10 ;
			data[91470] <= 8'h10 ;
			data[91471] <= 8'h10 ;
			data[91472] <= 8'h10 ;
			data[91473] <= 8'h10 ;
			data[91474] <= 8'h10 ;
			data[91475] <= 8'h10 ;
			data[91476] <= 8'h10 ;
			data[91477] <= 8'h10 ;
			data[91478] <= 8'h10 ;
			data[91479] <= 8'h10 ;
			data[91480] <= 8'h10 ;
			data[91481] <= 8'h10 ;
			data[91482] <= 8'h10 ;
			data[91483] <= 8'h10 ;
			data[91484] <= 8'h10 ;
			data[91485] <= 8'h10 ;
			data[91486] <= 8'h10 ;
			data[91487] <= 8'h10 ;
			data[91488] <= 8'h10 ;
			data[91489] <= 8'h10 ;
			data[91490] <= 8'h10 ;
			data[91491] <= 8'h10 ;
			data[91492] <= 8'h10 ;
			data[91493] <= 8'h10 ;
			data[91494] <= 8'h10 ;
			data[91495] <= 8'h10 ;
			data[91496] <= 8'h10 ;
			data[91497] <= 8'h10 ;
			data[91498] <= 8'h10 ;
			data[91499] <= 8'h10 ;
			data[91500] <= 8'h10 ;
			data[91501] <= 8'h10 ;
			data[91502] <= 8'h10 ;
			data[91503] <= 8'h10 ;
			data[91504] <= 8'h10 ;
			data[91505] <= 8'h10 ;
			data[91506] <= 8'h10 ;
			data[91507] <= 8'h10 ;
			data[91508] <= 8'h10 ;
			data[91509] <= 8'h10 ;
			data[91510] <= 8'h10 ;
			data[91511] <= 8'h10 ;
			data[91512] <= 8'h10 ;
			data[91513] <= 8'h10 ;
			data[91514] <= 8'h10 ;
			data[91515] <= 8'h10 ;
			data[91516] <= 8'h10 ;
			data[91517] <= 8'h10 ;
			data[91518] <= 8'h10 ;
			data[91519] <= 8'h10 ;
			data[91520] <= 8'h10 ;
			data[91521] <= 8'h10 ;
			data[91522] <= 8'h10 ;
			data[91523] <= 8'h10 ;
			data[91524] <= 8'h10 ;
			data[91525] <= 8'h10 ;
			data[91526] <= 8'h10 ;
			data[91527] <= 8'h10 ;
			data[91528] <= 8'h10 ;
			data[91529] <= 8'h10 ;
			data[91530] <= 8'h10 ;
			data[91531] <= 8'h10 ;
			data[91532] <= 8'h10 ;
			data[91533] <= 8'h10 ;
			data[91534] <= 8'h10 ;
			data[91535] <= 8'h10 ;
			data[91536] <= 8'h10 ;
			data[91537] <= 8'h10 ;
			data[91538] <= 8'h10 ;
			data[91539] <= 8'h10 ;
			data[91540] <= 8'h10 ;
			data[91541] <= 8'h10 ;
			data[91542] <= 8'h10 ;
			data[91543] <= 8'h10 ;
			data[91544] <= 8'h10 ;
			data[91545] <= 8'h10 ;
			data[91546] <= 8'h10 ;
			data[91547] <= 8'h10 ;
			data[91548] <= 8'h10 ;
			data[91549] <= 8'h10 ;
			data[91550] <= 8'h10 ;
			data[91551] <= 8'h10 ;
			data[91552] <= 8'h10 ;
			data[91553] <= 8'h10 ;
			data[91554] <= 8'h10 ;
			data[91555] <= 8'h10 ;
			data[91556] <= 8'h10 ;
			data[91557] <= 8'h10 ;
			data[91558] <= 8'h10 ;
			data[91559] <= 8'h10 ;
			data[91560] <= 8'h10 ;
			data[91561] <= 8'h10 ;
			data[91562] <= 8'h10 ;
			data[91563] <= 8'h10 ;
			data[91564] <= 8'h10 ;
			data[91565] <= 8'h10 ;
			data[91566] <= 8'h10 ;
			data[91567] <= 8'h10 ;
			data[91568] <= 8'h10 ;
			data[91569] <= 8'h10 ;
			data[91570] <= 8'h10 ;
			data[91571] <= 8'h10 ;
			data[91572] <= 8'h10 ;
			data[91573] <= 8'h10 ;
			data[91574] <= 8'h10 ;
			data[91575] <= 8'h10 ;
			data[91576] <= 8'h10 ;
			data[91577] <= 8'h10 ;
			data[91578] <= 8'h10 ;
			data[91579] <= 8'h10 ;
			data[91580] <= 8'h10 ;
			data[91581] <= 8'h10 ;
			data[91582] <= 8'h10 ;
			data[91583] <= 8'h10 ;
			data[91584] <= 8'h10 ;
			data[91585] <= 8'h10 ;
			data[91586] <= 8'h10 ;
			data[91587] <= 8'h10 ;
			data[91588] <= 8'h10 ;
			data[91589] <= 8'h10 ;
			data[91590] <= 8'h10 ;
			data[91591] <= 8'h10 ;
			data[91592] <= 8'h10 ;
			data[91593] <= 8'h10 ;
			data[91594] <= 8'h10 ;
			data[91595] <= 8'h10 ;
			data[91596] <= 8'h10 ;
			data[91597] <= 8'h10 ;
			data[91598] <= 8'h10 ;
			data[91599] <= 8'h10 ;
			data[91600] <= 8'h10 ;
			data[91601] <= 8'h10 ;
			data[91602] <= 8'h10 ;
			data[91603] <= 8'h10 ;
			data[91604] <= 8'h10 ;
			data[91605] <= 8'h10 ;
			data[91606] <= 8'h10 ;
			data[91607] <= 8'h10 ;
			data[91608] <= 8'h10 ;
			data[91609] <= 8'h10 ;
			data[91610] <= 8'h10 ;
			data[91611] <= 8'h10 ;
			data[91612] <= 8'h10 ;
			data[91613] <= 8'h10 ;
			data[91614] <= 8'h10 ;
			data[91615] <= 8'h10 ;
			data[91616] <= 8'h10 ;
			data[91617] <= 8'h10 ;
			data[91618] <= 8'h10 ;
			data[91619] <= 8'h10 ;
			data[91620] <= 8'h10 ;
			data[91621] <= 8'h10 ;
			data[91622] <= 8'h10 ;
			data[91623] <= 8'h10 ;
			data[91624] <= 8'h10 ;
			data[91625] <= 8'h10 ;
			data[91626] <= 8'h10 ;
			data[91627] <= 8'h10 ;
			data[91628] <= 8'h10 ;
			data[91629] <= 8'h10 ;
			data[91630] <= 8'h10 ;
			data[91631] <= 8'h10 ;
			data[91632] <= 8'h10 ;
			data[91633] <= 8'h10 ;
			data[91634] <= 8'h10 ;
			data[91635] <= 8'h10 ;
			data[91636] <= 8'h10 ;
			data[91637] <= 8'h10 ;
			data[91638] <= 8'h10 ;
			data[91639] <= 8'h10 ;
			data[91640] <= 8'h10 ;
			data[91641] <= 8'h10 ;
			data[91642] <= 8'h10 ;
			data[91643] <= 8'h10 ;
			data[91644] <= 8'h10 ;
			data[91645] <= 8'h10 ;
			data[91646] <= 8'h10 ;
			data[91647] <= 8'h10 ;
			data[91648] <= 8'h10 ;
			data[91649] <= 8'h10 ;
			data[91650] <= 8'h10 ;
			data[91651] <= 8'h10 ;
			data[91652] <= 8'h10 ;
			data[91653] <= 8'h10 ;
			data[91654] <= 8'h10 ;
			data[91655] <= 8'h10 ;
			data[91656] <= 8'h10 ;
			data[91657] <= 8'h10 ;
			data[91658] <= 8'h10 ;
			data[91659] <= 8'h10 ;
			data[91660] <= 8'h10 ;
			data[91661] <= 8'h10 ;
			data[91662] <= 8'h10 ;
			data[91663] <= 8'h10 ;
			data[91664] <= 8'h10 ;
			data[91665] <= 8'h10 ;
			data[91666] <= 8'h10 ;
			data[91667] <= 8'h10 ;
			data[91668] <= 8'h10 ;
			data[91669] <= 8'h10 ;
			data[91670] <= 8'h10 ;
			data[91671] <= 8'h10 ;
			data[91672] <= 8'h10 ;
			data[91673] <= 8'h10 ;
			data[91674] <= 8'h10 ;
			data[91675] <= 8'h10 ;
			data[91676] <= 8'h10 ;
			data[91677] <= 8'h10 ;
			data[91678] <= 8'h10 ;
			data[91679] <= 8'h10 ;
			data[91680] <= 8'h10 ;
			data[91681] <= 8'h10 ;
			data[91682] <= 8'h10 ;
			data[91683] <= 8'h10 ;
			data[91684] <= 8'h10 ;
			data[91685] <= 8'h10 ;
			data[91686] <= 8'h10 ;
			data[91687] <= 8'h10 ;
			data[91688] <= 8'h10 ;
			data[91689] <= 8'h10 ;
			data[91690] <= 8'h10 ;
			data[91691] <= 8'h10 ;
			data[91692] <= 8'h10 ;
			data[91693] <= 8'h10 ;
			data[91694] <= 8'h10 ;
			data[91695] <= 8'h10 ;
			data[91696] <= 8'h10 ;
			data[91697] <= 8'h10 ;
			data[91698] <= 8'h10 ;
			data[91699] <= 8'h10 ;
			data[91700] <= 8'h10 ;
			data[91701] <= 8'h10 ;
			data[91702] <= 8'h10 ;
			data[91703] <= 8'h10 ;
			data[91704] <= 8'h10 ;
			data[91705] <= 8'h10 ;
			data[91706] <= 8'h10 ;
			data[91707] <= 8'h10 ;
			data[91708] <= 8'h10 ;
			data[91709] <= 8'h10 ;
			data[91710] <= 8'h10 ;
			data[91711] <= 8'h10 ;
			data[91712] <= 8'h10 ;
			data[91713] <= 8'h10 ;
			data[91714] <= 8'h10 ;
			data[91715] <= 8'h10 ;
			data[91716] <= 8'h10 ;
			data[91717] <= 8'h10 ;
			data[91718] <= 8'h10 ;
			data[91719] <= 8'h10 ;
			data[91720] <= 8'h10 ;
			data[91721] <= 8'h10 ;
			data[91722] <= 8'h10 ;
			data[91723] <= 8'h10 ;
			data[91724] <= 8'h10 ;
			data[91725] <= 8'h10 ;
			data[91726] <= 8'h10 ;
			data[91727] <= 8'h10 ;
			data[91728] <= 8'h10 ;
			data[91729] <= 8'h10 ;
			data[91730] <= 8'h10 ;
			data[91731] <= 8'h10 ;
			data[91732] <= 8'h10 ;
			data[91733] <= 8'h10 ;
			data[91734] <= 8'h10 ;
			data[91735] <= 8'h10 ;
			data[91736] <= 8'h10 ;
			data[91737] <= 8'h10 ;
			data[91738] <= 8'h10 ;
			data[91739] <= 8'h10 ;
			data[91740] <= 8'h10 ;
			data[91741] <= 8'h10 ;
			data[91742] <= 8'h10 ;
			data[91743] <= 8'h10 ;
			data[91744] <= 8'h10 ;
			data[91745] <= 8'h10 ;
			data[91746] <= 8'h10 ;
			data[91747] <= 8'h10 ;
			data[91748] <= 8'h10 ;
			data[91749] <= 8'h10 ;
			data[91750] <= 8'h10 ;
			data[91751] <= 8'h10 ;
			data[91752] <= 8'h10 ;
			data[91753] <= 8'h10 ;
			data[91754] <= 8'h10 ;
			data[91755] <= 8'h10 ;
			data[91756] <= 8'h10 ;
			data[91757] <= 8'h10 ;
			data[91758] <= 8'h10 ;
			data[91759] <= 8'h10 ;
			data[91760] <= 8'h10 ;
			data[91761] <= 8'h10 ;
			data[91762] <= 8'h10 ;
			data[91763] <= 8'h10 ;
			data[91764] <= 8'h10 ;
			data[91765] <= 8'h10 ;
			data[91766] <= 8'h10 ;
			data[91767] <= 8'h10 ;
			data[91768] <= 8'h10 ;
			data[91769] <= 8'h10 ;
			data[91770] <= 8'h10 ;
			data[91771] <= 8'h10 ;
			data[91772] <= 8'h10 ;
			data[91773] <= 8'h10 ;
			data[91774] <= 8'h10 ;
			data[91775] <= 8'h10 ;
			data[91776] <= 8'h10 ;
			data[91777] <= 8'h10 ;
			data[91778] <= 8'h10 ;
			data[91779] <= 8'h10 ;
			data[91780] <= 8'h10 ;
			data[91781] <= 8'h10 ;
			data[91782] <= 8'h10 ;
			data[91783] <= 8'h10 ;
			data[91784] <= 8'h10 ;
			data[91785] <= 8'h10 ;
			data[91786] <= 8'h10 ;
			data[91787] <= 8'h10 ;
			data[91788] <= 8'h10 ;
			data[91789] <= 8'h10 ;
			data[91790] <= 8'h10 ;
			data[91791] <= 8'h10 ;
			data[91792] <= 8'h10 ;
			data[91793] <= 8'h10 ;
			data[91794] <= 8'h10 ;
			data[91795] <= 8'h10 ;
			data[91796] <= 8'h10 ;
			data[91797] <= 8'h10 ;
			data[91798] <= 8'h10 ;
			data[91799] <= 8'h10 ;
			data[91800] <= 8'h10 ;
			data[91801] <= 8'h10 ;
			data[91802] <= 8'h10 ;
			data[91803] <= 8'h10 ;
			data[91804] <= 8'h10 ;
			data[91805] <= 8'h10 ;
			data[91806] <= 8'h10 ;
			data[91807] <= 8'h10 ;
			data[91808] <= 8'h10 ;
			data[91809] <= 8'h10 ;
			data[91810] <= 8'h10 ;
			data[91811] <= 8'h10 ;
			data[91812] <= 8'h10 ;
			data[91813] <= 8'h10 ;
			data[91814] <= 8'h10 ;
			data[91815] <= 8'h10 ;
			data[91816] <= 8'h10 ;
			data[91817] <= 8'h10 ;
			data[91818] <= 8'h10 ;
			data[91819] <= 8'h10 ;
			data[91820] <= 8'h10 ;
			data[91821] <= 8'h10 ;
			data[91822] <= 8'h10 ;
			data[91823] <= 8'h10 ;
			data[91824] <= 8'h10 ;
			data[91825] <= 8'h10 ;
			data[91826] <= 8'h10 ;
			data[91827] <= 8'h10 ;
			data[91828] <= 8'h10 ;
			data[91829] <= 8'h10 ;
			data[91830] <= 8'h10 ;
			data[91831] <= 8'h10 ;
			data[91832] <= 8'h10 ;
			data[91833] <= 8'h10 ;
			data[91834] <= 8'h10 ;
			data[91835] <= 8'h10 ;
			data[91836] <= 8'h10 ;
			data[91837] <= 8'h10 ;
			data[91838] <= 8'h10 ;
			data[91839] <= 8'h10 ;
			data[91840] <= 8'h10 ;
			data[91841] <= 8'h10 ;
			data[91842] <= 8'h10 ;
			data[91843] <= 8'h10 ;
			data[91844] <= 8'h10 ;
			data[91845] <= 8'h10 ;
			data[91846] <= 8'h10 ;
			data[91847] <= 8'h10 ;
			data[91848] <= 8'h10 ;
			data[91849] <= 8'h10 ;
			data[91850] <= 8'h10 ;
			data[91851] <= 8'h10 ;
			data[91852] <= 8'h10 ;
			data[91853] <= 8'h10 ;
			data[91854] <= 8'h10 ;
			data[91855] <= 8'h10 ;
			data[91856] <= 8'h10 ;
			data[91857] <= 8'h10 ;
			data[91858] <= 8'h10 ;
			data[91859] <= 8'h10 ;
			data[91860] <= 8'h10 ;
			data[91861] <= 8'h10 ;
			data[91862] <= 8'h10 ;
			data[91863] <= 8'h10 ;
			data[91864] <= 8'h10 ;
			data[91865] <= 8'h10 ;
			data[91866] <= 8'h10 ;
			data[91867] <= 8'h10 ;
			data[91868] <= 8'h10 ;
			data[91869] <= 8'h10 ;
			data[91870] <= 8'h10 ;
			data[91871] <= 8'h10 ;
			data[91872] <= 8'h10 ;
			data[91873] <= 8'h10 ;
			data[91874] <= 8'h10 ;
			data[91875] <= 8'h10 ;
			data[91876] <= 8'h10 ;
			data[91877] <= 8'h10 ;
			data[91878] <= 8'h10 ;
			data[91879] <= 8'h10 ;
			data[91880] <= 8'h10 ;
			data[91881] <= 8'h10 ;
			data[91882] <= 8'h10 ;
			data[91883] <= 8'h10 ;
			data[91884] <= 8'h10 ;
			data[91885] <= 8'h10 ;
			data[91886] <= 8'h10 ;
			data[91887] <= 8'h10 ;
			data[91888] <= 8'h10 ;
			data[91889] <= 8'h10 ;
			data[91890] <= 8'h10 ;
			data[91891] <= 8'h10 ;
			data[91892] <= 8'h10 ;
			data[91893] <= 8'h10 ;
			data[91894] <= 8'h10 ;
			data[91895] <= 8'h10 ;
			data[91896] <= 8'h10 ;
			data[91897] <= 8'h10 ;
			data[91898] <= 8'h10 ;
			data[91899] <= 8'h10 ;
			data[91900] <= 8'h10 ;
			data[91901] <= 8'h10 ;
			data[91902] <= 8'h10 ;
			data[91903] <= 8'h10 ;
			data[91904] <= 8'h10 ;
			data[91905] <= 8'h10 ;
			data[91906] <= 8'h10 ;
			data[91907] <= 8'h10 ;
			data[91908] <= 8'h10 ;
			data[91909] <= 8'h10 ;
			data[91910] <= 8'h10 ;
			data[91911] <= 8'h10 ;
			data[91912] <= 8'h10 ;
			data[91913] <= 8'h10 ;
			data[91914] <= 8'h10 ;
			data[91915] <= 8'h10 ;
			data[91916] <= 8'h10 ;
			data[91917] <= 8'h10 ;
			data[91918] <= 8'h10 ;
			data[91919] <= 8'h10 ;
			data[91920] <= 8'h10 ;
			data[91921] <= 8'h10 ;
			data[91922] <= 8'h10 ;
			data[91923] <= 8'h10 ;
			data[91924] <= 8'h10 ;
			data[91925] <= 8'h10 ;
			data[91926] <= 8'h10 ;
			data[91927] <= 8'h10 ;
			data[91928] <= 8'h10 ;
			data[91929] <= 8'h10 ;
			data[91930] <= 8'h10 ;
			data[91931] <= 8'h10 ;
			data[91932] <= 8'h10 ;
			data[91933] <= 8'h10 ;
			data[91934] <= 8'h10 ;
			data[91935] <= 8'h10 ;
			data[91936] <= 8'h10 ;
			data[91937] <= 8'h10 ;
			data[91938] <= 8'h10 ;
			data[91939] <= 8'h10 ;
			data[91940] <= 8'h10 ;
			data[91941] <= 8'h10 ;
			data[91942] <= 8'h10 ;
			data[91943] <= 8'h10 ;
			data[91944] <= 8'h10 ;
			data[91945] <= 8'h10 ;
			data[91946] <= 8'h10 ;
			data[91947] <= 8'h10 ;
			data[91948] <= 8'h10 ;
			data[91949] <= 8'h10 ;
			data[91950] <= 8'h10 ;
			data[91951] <= 8'h10 ;
			data[91952] <= 8'h10 ;
			data[91953] <= 8'h10 ;
			data[91954] <= 8'h10 ;
			data[91955] <= 8'h10 ;
			data[91956] <= 8'h10 ;
			data[91957] <= 8'h10 ;
			data[91958] <= 8'h10 ;
			data[91959] <= 8'h10 ;
			data[91960] <= 8'h10 ;
			data[91961] <= 8'h10 ;
			data[91962] <= 8'h10 ;
			data[91963] <= 8'h10 ;
			data[91964] <= 8'h10 ;
			data[91965] <= 8'h10 ;
			data[91966] <= 8'h10 ;
			data[91967] <= 8'h10 ;
			data[91968] <= 8'h10 ;
			data[91969] <= 8'h10 ;
			data[91970] <= 8'h10 ;
			data[91971] <= 8'h10 ;
			data[91972] <= 8'h10 ;
			data[91973] <= 8'h10 ;
			data[91974] <= 8'h10 ;
			data[91975] <= 8'h10 ;
			data[91976] <= 8'h10 ;
			data[91977] <= 8'h10 ;
			data[91978] <= 8'h10 ;
			data[91979] <= 8'h10 ;
			data[91980] <= 8'h10 ;
			data[91981] <= 8'h10 ;
			data[91982] <= 8'h10 ;
			data[91983] <= 8'h10 ;
			data[91984] <= 8'h10 ;
			data[91985] <= 8'h10 ;
			data[91986] <= 8'h10 ;
			data[91987] <= 8'h10 ;
			data[91988] <= 8'h10 ;
			data[91989] <= 8'h10 ;
			data[91990] <= 8'h10 ;
			data[91991] <= 8'h10 ;
			data[91992] <= 8'h10 ;
			data[91993] <= 8'h10 ;
			data[91994] <= 8'h10 ;
			data[91995] <= 8'h10 ;
			data[91996] <= 8'h10 ;
			data[91997] <= 8'h10 ;
			data[91998] <= 8'h10 ;
			data[91999] <= 8'h10 ;
			data[92000] <= 8'h10 ;
			data[92001] <= 8'h10 ;
			data[92002] <= 8'h10 ;
			data[92003] <= 8'h10 ;
			data[92004] <= 8'h10 ;
			data[92005] <= 8'h10 ;
			data[92006] <= 8'h10 ;
			data[92007] <= 8'h10 ;
			data[92008] <= 8'h10 ;
			data[92009] <= 8'h10 ;
			data[92010] <= 8'h10 ;
			data[92011] <= 8'h10 ;
			data[92012] <= 8'h10 ;
			data[92013] <= 8'h10 ;
			data[92014] <= 8'h10 ;
			data[92015] <= 8'h10 ;
			data[92016] <= 8'h10 ;
			data[92017] <= 8'h10 ;
			data[92018] <= 8'h10 ;
			data[92019] <= 8'h10 ;
			data[92020] <= 8'h10 ;
			data[92021] <= 8'h10 ;
			data[92022] <= 8'h10 ;
			data[92023] <= 8'h10 ;
			data[92024] <= 8'h10 ;
			data[92025] <= 8'h10 ;
			data[92026] <= 8'h10 ;
			data[92027] <= 8'h10 ;
			data[92028] <= 8'h10 ;
			data[92029] <= 8'h10 ;
			data[92030] <= 8'h10 ;
			data[92031] <= 8'h10 ;
			data[92032] <= 8'h10 ;
			data[92033] <= 8'h10 ;
			data[92034] <= 8'h10 ;
			data[92035] <= 8'h10 ;
			data[92036] <= 8'h10 ;
			data[92037] <= 8'h10 ;
			data[92038] <= 8'h10 ;
			data[92039] <= 8'h10 ;
			data[92040] <= 8'h10 ;
			data[92041] <= 8'h10 ;
			data[92042] <= 8'h10 ;
			data[92043] <= 8'h10 ;
			data[92044] <= 8'h10 ;
			data[92045] <= 8'h10 ;
			data[92046] <= 8'h10 ;
			data[92047] <= 8'h10 ;
			data[92048] <= 8'h10 ;
			data[92049] <= 8'h10 ;
			data[92050] <= 8'h10 ;
			data[92051] <= 8'h10 ;
			data[92052] <= 8'h10 ;
			data[92053] <= 8'h10 ;
			data[92054] <= 8'h10 ;
			data[92055] <= 8'h10 ;
			data[92056] <= 8'h10 ;
			data[92057] <= 8'h10 ;
			data[92058] <= 8'h10 ;
			data[92059] <= 8'h10 ;
			data[92060] <= 8'h10 ;
			data[92061] <= 8'h10 ;
			data[92062] <= 8'h10 ;
			data[92063] <= 8'h10 ;
			data[92064] <= 8'h10 ;
			data[92065] <= 8'h10 ;
			data[92066] <= 8'h10 ;
			data[92067] <= 8'h10 ;
			data[92068] <= 8'h10 ;
			data[92069] <= 8'h10 ;
			data[92070] <= 8'h10 ;
			data[92071] <= 8'h10 ;
			data[92072] <= 8'h10 ;
			data[92073] <= 8'h10 ;
			data[92074] <= 8'h10 ;
			data[92075] <= 8'h10 ;
			data[92076] <= 8'h10 ;
			data[92077] <= 8'h10 ;
			data[92078] <= 8'h10 ;
			data[92079] <= 8'h10 ;
			data[92080] <= 8'h10 ;
			data[92081] <= 8'h10 ;
			data[92082] <= 8'h10 ;
			data[92083] <= 8'h10 ;
			data[92084] <= 8'h10 ;
			data[92085] <= 8'h10 ;
			data[92086] <= 8'h10 ;
			data[92087] <= 8'h10 ;
			data[92088] <= 8'h10 ;
			data[92089] <= 8'h10 ;
			data[92090] <= 8'h10 ;
			data[92091] <= 8'h10 ;
			data[92092] <= 8'h10 ;
			data[92093] <= 8'h10 ;
			data[92094] <= 8'h10 ;
			data[92095] <= 8'h10 ;
			data[92096] <= 8'h10 ;
			data[92097] <= 8'h10 ;
			data[92098] <= 8'h10 ;
			data[92099] <= 8'h10 ;
			data[92100] <= 8'h10 ;
			data[92101] <= 8'h10 ;
			data[92102] <= 8'h10 ;
			data[92103] <= 8'h10 ;
			data[92104] <= 8'h10 ;
			data[92105] <= 8'h10 ;
			data[92106] <= 8'h10 ;
			data[92107] <= 8'h10 ;
			data[92108] <= 8'h10 ;
			data[92109] <= 8'h10 ;
			data[92110] <= 8'h10 ;
			data[92111] <= 8'h10 ;
			data[92112] <= 8'h10 ;
			data[92113] <= 8'h10 ;
			data[92114] <= 8'h10 ;
			data[92115] <= 8'h10 ;
			data[92116] <= 8'h10 ;
			data[92117] <= 8'h10 ;
			data[92118] <= 8'h10 ;
			data[92119] <= 8'h10 ;
			data[92120] <= 8'h10 ;
			data[92121] <= 8'h10 ;
			data[92122] <= 8'h10 ;
			data[92123] <= 8'h10 ;
			data[92124] <= 8'h10 ;
			data[92125] <= 8'h10 ;
			data[92126] <= 8'h10 ;
			data[92127] <= 8'h10 ;
			data[92128] <= 8'h10 ;
			data[92129] <= 8'h10 ;
			data[92130] <= 8'h10 ;
			data[92131] <= 8'h10 ;
			data[92132] <= 8'h10 ;
			data[92133] <= 8'h10 ;
			data[92134] <= 8'h10 ;
			data[92135] <= 8'h10 ;
			data[92136] <= 8'h10 ;
			data[92137] <= 8'h10 ;
			data[92138] <= 8'h10 ;
			data[92139] <= 8'h10 ;
			data[92140] <= 8'h10 ;
			data[92141] <= 8'h10 ;
			data[92142] <= 8'h10 ;
			data[92143] <= 8'h10 ;
			data[92144] <= 8'h10 ;
			data[92145] <= 8'h10 ;
			data[92146] <= 8'h10 ;
			data[92147] <= 8'h10 ;
			data[92148] <= 8'h10 ;
			data[92149] <= 8'h10 ;
			data[92150] <= 8'h10 ;
			data[92151] <= 8'h10 ;
			data[92152] <= 8'h10 ;
			data[92153] <= 8'h10 ;
			data[92154] <= 8'h10 ;
			data[92155] <= 8'h10 ;
			data[92156] <= 8'h10 ;
			data[92157] <= 8'h10 ;
			data[92158] <= 8'h10 ;
			data[92159] <= 8'h10 ;
			data[92160] <= 8'h10 ;
			data[92161] <= 8'h10 ;
			data[92162] <= 8'h10 ;
			data[92163] <= 8'h10 ;
			data[92164] <= 8'h10 ;
			data[92165] <= 8'h10 ;
			data[92166] <= 8'h10 ;
			data[92167] <= 8'h10 ;
			data[92168] <= 8'h10 ;
			data[92169] <= 8'h10 ;
			data[92170] <= 8'h10 ;
			data[92171] <= 8'h10 ;
			data[92172] <= 8'h10 ;
			data[92173] <= 8'h10 ;
			data[92174] <= 8'h10 ;
			data[92175] <= 8'h10 ;
			data[92176] <= 8'h10 ;
			data[92177] <= 8'h10 ;
			data[92178] <= 8'h10 ;
			data[92179] <= 8'h10 ;
			data[92180] <= 8'h10 ;
			data[92181] <= 8'h10 ;
			data[92182] <= 8'h10 ;
			data[92183] <= 8'h10 ;
			data[92184] <= 8'h10 ;
			data[92185] <= 8'h10 ;
			data[92186] <= 8'h10 ;
			data[92187] <= 8'h10 ;
			data[92188] <= 8'h10 ;
			data[92189] <= 8'h10 ;
			data[92190] <= 8'h10 ;
			data[92191] <= 8'h10 ;
			data[92192] <= 8'h10 ;
			data[92193] <= 8'h10 ;
			data[92194] <= 8'h10 ;
			data[92195] <= 8'h10 ;
			data[92196] <= 8'h10 ;
			data[92197] <= 8'h10 ;
			data[92198] <= 8'h10 ;
			data[92199] <= 8'h10 ;
			data[92200] <= 8'h10 ;
			data[92201] <= 8'h10 ;
			data[92202] <= 8'h10 ;
			data[92203] <= 8'h10 ;
			data[92204] <= 8'h10 ;
			data[92205] <= 8'h10 ;
			data[92206] <= 8'h10 ;
			data[92207] <= 8'h10 ;
			data[92208] <= 8'h10 ;
			data[92209] <= 8'h10 ;
			data[92210] <= 8'h10 ;
			data[92211] <= 8'h10 ;
			data[92212] <= 8'h10 ;
			data[92213] <= 8'h10 ;
			data[92214] <= 8'h10 ;
			data[92215] <= 8'h10 ;
			data[92216] <= 8'h10 ;
			data[92217] <= 8'h10 ;
			data[92218] <= 8'h10 ;
			data[92219] <= 8'h10 ;
			data[92220] <= 8'h10 ;
			data[92221] <= 8'h10 ;
			data[92222] <= 8'h10 ;
			data[92223] <= 8'h10 ;
			data[92224] <= 8'h10 ;
			data[92225] <= 8'h10 ;
			data[92226] <= 8'h10 ;
			data[92227] <= 8'h10 ;
			data[92228] <= 8'h10 ;
			data[92229] <= 8'h10 ;
			data[92230] <= 8'h10 ;
			data[92231] <= 8'h10 ;
			data[92232] <= 8'h10 ;
			data[92233] <= 8'h10 ;
			data[92234] <= 8'h10 ;
			data[92235] <= 8'h10 ;
			data[92236] <= 8'h10 ;
			data[92237] <= 8'h10 ;
			data[92238] <= 8'h10 ;
			data[92239] <= 8'h10 ;
			data[92240] <= 8'h10 ;
			data[92241] <= 8'h10 ;
			data[92242] <= 8'h10 ;
			data[92243] <= 8'h10 ;
			data[92244] <= 8'h10 ;
			data[92245] <= 8'h10 ;
			data[92246] <= 8'h10 ;
			data[92247] <= 8'h10 ;
			data[92248] <= 8'h10 ;
			data[92249] <= 8'h10 ;
			data[92250] <= 8'h10 ;
			data[92251] <= 8'h10 ;
			data[92252] <= 8'h10 ;
			data[92253] <= 8'h10 ;
			data[92254] <= 8'h10 ;
			data[92255] <= 8'h10 ;
			data[92256] <= 8'h10 ;
			data[92257] <= 8'h10 ;
			data[92258] <= 8'h10 ;
			data[92259] <= 8'h10 ;
			data[92260] <= 8'h10 ;
			data[92261] <= 8'h10 ;
			data[92262] <= 8'h10 ;
			data[92263] <= 8'h10 ;
			data[92264] <= 8'h10 ;
			data[92265] <= 8'h10 ;
			data[92266] <= 8'h10 ;
			data[92267] <= 8'h10 ;
			data[92268] <= 8'h10 ;
			data[92269] <= 8'h10 ;
			data[92270] <= 8'h10 ;
			data[92271] <= 8'h10 ;
			data[92272] <= 8'h10 ;
			data[92273] <= 8'h10 ;
			data[92274] <= 8'h10 ;
			data[92275] <= 8'h10 ;
			data[92276] <= 8'h10 ;
			data[92277] <= 8'h10 ;
			data[92278] <= 8'h10 ;
			data[92279] <= 8'h10 ;
			data[92280] <= 8'h10 ;
			data[92281] <= 8'h10 ;
			data[92282] <= 8'h10 ;
			data[92283] <= 8'h10 ;
			data[92284] <= 8'h10 ;
			data[92285] <= 8'h10 ;
			data[92286] <= 8'h10 ;
			data[92287] <= 8'h10 ;
			data[92288] <= 8'h10 ;
			data[92289] <= 8'h10 ;
			data[92290] <= 8'h10 ;
			data[92291] <= 8'h10 ;
			data[92292] <= 8'h10 ;
			data[92293] <= 8'h10 ;
			data[92294] <= 8'h10 ;
			data[92295] <= 8'h10 ;
			data[92296] <= 8'h10 ;
			data[92297] <= 8'h10 ;
			data[92298] <= 8'h10 ;
			data[92299] <= 8'h10 ;
			data[92300] <= 8'h10 ;
			data[92301] <= 8'h10 ;
			data[92302] <= 8'h10 ;
			data[92303] <= 8'h10 ;
			data[92304] <= 8'h10 ;
			data[92305] <= 8'h10 ;
			data[92306] <= 8'h10 ;
			data[92307] <= 8'h10 ;
			data[92308] <= 8'h10 ;
			data[92309] <= 8'h10 ;
			data[92310] <= 8'h10 ;
			data[92311] <= 8'h10 ;
			data[92312] <= 8'h10 ;
			data[92313] <= 8'h10 ;
			data[92314] <= 8'h10 ;
			data[92315] <= 8'h10 ;
			data[92316] <= 8'h10 ;
			data[92317] <= 8'h10 ;
			data[92318] <= 8'h10 ;
			data[92319] <= 8'h10 ;
			data[92320] <= 8'h10 ;
			data[92321] <= 8'h10 ;
			data[92322] <= 8'h10 ;
			data[92323] <= 8'h10 ;
			data[92324] <= 8'h10 ;
			data[92325] <= 8'h10 ;
			data[92326] <= 8'h10 ;
			data[92327] <= 8'h10 ;
			data[92328] <= 8'h10 ;
			data[92329] <= 8'h10 ;
			data[92330] <= 8'h10 ;
			data[92331] <= 8'h10 ;
			data[92332] <= 8'h10 ;
			data[92333] <= 8'h10 ;
			data[92334] <= 8'h10 ;
			data[92335] <= 8'h10 ;
			data[92336] <= 8'h10 ;
			data[92337] <= 8'h10 ;
			data[92338] <= 8'h10 ;
			data[92339] <= 8'h10 ;
			data[92340] <= 8'h10 ;
			data[92341] <= 8'h10 ;
			data[92342] <= 8'h10 ;
			data[92343] <= 8'h10 ;
			data[92344] <= 8'h10 ;
			data[92345] <= 8'h10 ;
			data[92346] <= 8'h10 ;
			data[92347] <= 8'h10 ;
			data[92348] <= 8'h10 ;
			data[92349] <= 8'h10 ;
			data[92350] <= 8'h10 ;
			data[92351] <= 8'h10 ;
			data[92352] <= 8'h10 ;
			data[92353] <= 8'h10 ;
			data[92354] <= 8'h10 ;
			data[92355] <= 8'h10 ;
			data[92356] <= 8'h10 ;
			data[92357] <= 8'h10 ;
			data[92358] <= 8'h10 ;
			data[92359] <= 8'h10 ;
			data[92360] <= 8'h10 ;
			data[92361] <= 8'h10 ;
			data[92362] <= 8'h10 ;
			data[92363] <= 8'h10 ;
			data[92364] <= 8'h10 ;
			data[92365] <= 8'h10 ;
			data[92366] <= 8'h10 ;
			data[92367] <= 8'h10 ;
			data[92368] <= 8'h10 ;
			data[92369] <= 8'h10 ;
			data[92370] <= 8'h10 ;
			data[92371] <= 8'h10 ;
			data[92372] <= 8'h10 ;
			data[92373] <= 8'h10 ;
			data[92374] <= 8'h10 ;
			data[92375] <= 8'h10 ;
			data[92376] <= 8'h10 ;
			data[92377] <= 8'h10 ;
			data[92378] <= 8'h10 ;
			data[92379] <= 8'h10 ;
			data[92380] <= 8'h10 ;
			data[92381] <= 8'h10 ;
			data[92382] <= 8'h10 ;
			data[92383] <= 8'h10 ;
			data[92384] <= 8'h10 ;
			data[92385] <= 8'h10 ;
			data[92386] <= 8'h10 ;
			data[92387] <= 8'h10 ;
			data[92388] <= 8'h10 ;
			data[92389] <= 8'h10 ;
			data[92390] <= 8'h10 ;
			data[92391] <= 8'h10 ;
			data[92392] <= 8'h10 ;
			data[92393] <= 8'h10 ;
			data[92394] <= 8'h10 ;
			data[92395] <= 8'h10 ;
			data[92396] <= 8'h10 ;
			data[92397] <= 8'h10 ;
			data[92398] <= 8'h10 ;
			data[92399] <= 8'h10 ;
			data[92400] <= 8'h10 ;
			data[92401] <= 8'h10 ;
			data[92402] <= 8'h10 ;
			data[92403] <= 8'h10 ;
			data[92404] <= 8'h10 ;
			data[92405] <= 8'h10 ;
			data[92406] <= 8'h10 ;
			data[92407] <= 8'h10 ;
			data[92408] <= 8'h10 ;
			data[92409] <= 8'h10 ;
			data[92410] <= 8'h10 ;
			data[92411] <= 8'h10 ;
			data[92412] <= 8'h10 ;
			data[92413] <= 8'h10 ;
			data[92414] <= 8'h10 ;
			data[92415] <= 8'h10 ;
			data[92416] <= 8'h10 ;
			data[92417] <= 8'h10 ;
			data[92418] <= 8'h10 ;
			data[92419] <= 8'h10 ;
			data[92420] <= 8'h10 ;
			data[92421] <= 8'h10 ;
			data[92422] <= 8'h10 ;
			data[92423] <= 8'h10 ;
			data[92424] <= 8'h10 ;
			data[92425] <= 8'h10 ;
			data[92426] <= 8'h10 ;
			data[92427] <= 8'h10 ;
			data[92428] <= 8'h10 ;
			data[92429] <= 8'h10 ;
			data[92430] <= 8'h10 ;
			data[92431] <= 8'h10 ;
			data[92432] <= 8'h10 ;
			data[92433] <= 8'h10 ;
			data[92434] <= 8'h10 ;
			data[92435] <= 8'h10 ;
			data[92436] <= 8'h10 ;
			data[92437] <= 8'h10 ;
			data[92438] <= 8'h10 ;
			data[92439] <= 8'h10 ;
			data[92440] <= 8'h10 ;
			data[92441] <= 8'h10 ;
			data[92442] <= 8'h10 ;
			data[92443] <= 8'h10 ;
			data[92444] <= 8'h10 ;
			data[92445] <= 8'h10 ;
			data[92446] <= 8'h10 ;
			data[92447] <= 8'h10 ;
			data[92448] <= 8'h10 ;
			data[92449] <= 8'h10 ;
			data[92450] <= 8'h10 ;
			data[92451] <= 8'h10 ;
			data[92452] <= 8'h10 ;
			data[92453] <= 8'h10 ;
			data[92454] <= 8'h10 ;
			data[92455] <= 8'h10 ;
			data[92456] <= 8'h10 ;
			data[92457] <= 8'h10 ;
			data[92458] <= 8'h10 ;
			data[92459] <= 8'h10 ;
			data[92460] <= 8'h10 ;
			data[92461] <= 8'h10 ;
			data[92462] <= 8'h10 ;
			data[92463] <= 8'h10 ;
			data[92464] <= 8'h10 ;
			data[92465] <= 8'h10 ;
			data[92466] <= 8'h10 ;
			data[92467] <= 8'h10 ;
			data[92468] <= 8'h10 ;
			data[92469] <= 8'h10 ;
			data[92470] <= 8'h10 ;
			data[92471] <= 8'h10 ;
			data[92472] <= 8'h10 ;
			data[92473] <= 8'h10 ;
			data[92474] <= 8'h10 ;
			data[92475] <= 8'h10 ;
			data[92476] <= 8'h10 ;
			data[92477] <= 8'h10 ;
			data[92478] <= 8'h10 ;
			data[92479] <= 8'h10 ;
			data[92480] <= 8'h10 ;
			data[92481] <= 8'h10 ;
			data[92482] <= 8'h10 ;
			data[92483] <= 8'h10 ;
			data[92484] <= 8'h10 ;
			data[92485] <= 8'h10 ;
			data[92486] <= 8'h10 ;
			data[92487] <= 8'h10 ;
			data[92488] <= 8'h10 ;
			data[92489] <= 8'h10 ;
			data[92490] <= 8'h10 ;
			data[92491] <= 8'h10 ;
			data[92492] <= 8'h10 ;
			data[92493] <= 8'h10 ;
			data[92494] <= 8'h10 ;
			data[92495] <= 8'h10 ;
			data[92496] <= 8'h10 ;
			data[92497] <= 8'h10 ;
			data[92498] <= 8'h10 ;
			data[92499] <= 8'h10 ;
			data[92500] <= 8'h10 ;
			data[92501] <= 8'h10 ;
			data[92502] <= 8'h10 ;
			data[92503] <= 8'h10 ;
			data[92504] <= 8'h10 ;
			data[92505] <= 8'h10 ;
			data[92506] <= 8'h10 ;
			data[92507] <= 8'h10 ;
			data[92508] <= 8'h10 ;
			data[92509] <= 8'h10 ;
			data[92510] <= 8'h10 ;
			data[92511] <= 8'h10 ;
			data[92512] <= 8'h10 ;
			data[92513] <= 8'h10 ;
			data[92514] <= 8'h10 ;
			data[92515] <= 8'h10 ;
			data[92516] <= 8'h10 ;
			data[92517] <= 8'h10 ;
			data[92518] <= 8'h10 ;
			data[92519] <= 8'h10 ;
			data[92520] <= 8'h10 ;
			data[92521] <= 8'h10 ;
			data[92522] <= 8'h10 ;
			data[92523] <= 8'h10 ;
			data[92524] <= 8'h10 ;
			data[92525] <= 8'h10 ;
			data[92526] <= 8'h10 ;
			data[92527] <= 8'h10 ;
			data[92528] <= 8'h10 ;
			data[92529] <= 8'h10 ;
			data[92530] <= 8'h10 ;
			data[92531] <= 8'h10 ;
			data[92532] <= 8'h10 ;
			data[92533] <= 8'h10 ;
			data[92534] <= 8'h10 ;
			data[92535] <= 8'h10 ;
			data[92536] <= 8'h10 ;
			data[92537] <= 8'h10 ;
			data[92538] <= 8'h10 ;
			data[92539] <= 8'h10 ;
			data[92540] <= 8'h10 ;
			data[92541] <= 8'h10 ;
			data[92542] <= 8'h10 ;
			data[92543] <= 8'h10 ;
			data[92544] <= 8'h10 ;
			data[92545] <= 8'h10 ;
			data[92546] <= 8'h10 ;
			data[92547] <= 8'h10 ;
			data[92548] <= 8'h10 ;
			data[92549] <= 8'h10 ;
			data[92550] <= 8'h10 ;
			data[92551] <= 8'h10 ;
			data[92552] <= 8'h10 ;
			data[92553] <= 8'h10 ;
			data[92554] <= 8'h10 ;
			data[92555] <= 8'h10 ;
			data[92556] <= 8'h10 ;
			data[92557] <= 8'h10 ;
			data[92558] <= 8'h10 ;
			data[92559] <= 8'h10 ;
			data[92560] <= 8'h10 ;
			data[92561] <= 8'h10 ;
			data[92562] <= 8'h10 ;
			data[92563] <= 8'h10 ;
			data[92564] <= 8'h10 ;
			data[92565] <= 8'h10 ;
			data[92566] <= 8'h10 ;
			data[92567] <= 8'h10 ;
			data[92568] <= 8'h10 ;
			data[92569] <= 8'h10 ;
			data[92570] <= 8'h10 ;
			data[92571] <= 8'h10 ;
			data[92572] <= 8'h10 ;
			data[92573] <= 8'h10 ;
			data[92574] <= 8'h10 ;
			data[92575] <= 8'h10 ;
			data[92576] <= 8'h10 ;
			data[92577] <= 8'h10 ;
			data[92578] <= 8'h10 ;
			data[92579] <= 8'h10 ;
			data[92580] <= 8'h10 ;
			data[92581] <= 8'h10 ;
			data[92582] <= 8'h10 ;
			data[92583] <= 8'h10 ;
			data[92584] <= 8'h10 ;
			data[92585] <= 8'h10 ;
			data[92586] <= 8'h10 ;
			data[92587] <= 8'h10 ;
			data[92588] <= 8'h10 ;
			data[92589] <= 8'h10 ;
			data[92590] <= 8'h10 ;
			data[92591] <= 8'h10 ;
			data[92592] <= 8'h10 ;
			data[92593] <= 8'h10 ;
			data[92594] <= 8'h10 ;
			data[92595] <= 8'h10 ;
			data[92596] <= 8'h10 ;
			data[92597] <= 8'h10 ;
			data[92598] <= 8'h10 ;
			data[92599] <= 8'h10 ;
			data[92600] <= 8'h10 ;
			data[92601] <= 8'h10 ;
			data[92602] <= 8'h10 ;
			data[92603] <= 8'h10 ;
			data[92604] <= 8'h10 ;
			data[92605] <= 8'h10 ;
			data[92606] <= 8'h10 ;
			data[92607] <= 8'h10 ;
			data[92608] <= 8'h10 ;
			data[92609] <= 8'h10 ;
			data[92610] <= 8'h10 ;
			data[92611] <= 8'h10 ;
			data[92612] <= 8'h10 ;
			data[92613] <= 8'h10 ;
			data[92614] <= 8'h10 ;
			data[92615] <= 8'h10 ;
			data[92616] <= 8'h10 ;
			data[92617] <= 8'h10 ;
			data[92618] <= 8'h10 ;
			data[92619] <= 8'h10 ;
			data[92620] <= 8'h10 ;
			data[92621] <= 8'h10 ;
			data[92622] <= 8'h10 ;
			data[92623] <= 8'h10 ;
			data[92624] <= 8'h10 ;
			data[92625] <= 8'h10 ;
			data[92626] <= 8'h10 ;
			data[92627] <= 8'h10 ;
			data[92628] <= 8'h10 ;
			data[92629] <= 8'h10 ;
			data[92630] <= 8'h10 ;
			data[92631] <= 8'h10 ;
			data[92632] <= 8'h10 ;
			data[92633] <= 8'h10 ;
			data[92634] <= 8'h10 ;
			data[92635] <= 8'h10 ;
			data[92636] <= 8'h10 ;
			data[92637] <= 8'h10 ;
			data[92638] <= 8'h10 ;
			data[92639] <= 8'h10 ;
			data[92640] <= 8'h10 ;
			data[92641] <= 8'h10 ;
			data[92642] <= 8'h10 ;
			data[92643] <= 8'h10 ;
			data[92644] <= 8'h10 ;
			data[92645] <= 8'h10 ;
			data[92646] <= 8'h10 ;
			data[92647] <= 8'h10 ;
			data[92648] <= 8'h10 ;
			data[92649] <= 8'h10 ;
			data[92650] <= 8'h10 ;
			data[92651] <= 8'h10 ;
			data[92652] <= 8'h10 ;
			data[92653] <= 8'h10 ;
			data[92654] <= 8'h10 ;
			data[92655] <= 8'h10 ;
			data[92656] <= 8'h10 ;
			data[92657] <= 8'h10 ;
			data[92658] <= 8'h10 ;
			data[92659] <= 8'h10 ;
			data[92660] <= 8'h10 ;
			data[92661] <= 8'h10 ;
			data[92662] <= 8'h10 ;
			data[92663] <= 8'h10 ;
			data[92664] <= 8'h10 ;
			data[92665] <= 8'h10 ;
			data[92666] <= 8'h10 ;
			data[92667] <= 8'h10 ;
			data[92668] <= 8'h10 ;
			data[92669] <= 8'h10 ;
			data[92670] <= 8'h10 ;
			data[92671] <= 8'h10 ;
			data[92672] <= 8'h10 ;
			data[92673] <= 8'h10 ;
			data[92674] <= 8'h10 ;
			data[92675] <= 8'h10 ;
			data[92676] <= 8'h10 ;
			data[92677] <= 8'h10 ;
			data[92678] <= 8'h10 ;
			data[92679] <= 8'h10 ;
			data[92680] <= 8'h10 ;
			data[92681] <= 8'h10 ;
			data[92682] <= 8'h10 ;
			data[92683] <= 8'h10 ;
			data[92684] <= 8'h10 ;
			data[92685] <= 8'h10 ;
			data[92686] <= 8'h10 ;
			data[92687] <= 8'h10 ;
			data[92688] <= 8'h10 ;
			data[92689] <= 8'h10 ;
			data[92690] <= 8'h10 ;
			data[92691] <= 8'h10 ;
			data[92692] <= 8'h10 ;
			data[92693] <= 8'h10 ;
			data[92694] <= 8'h10 ;
			data[92695] <= 8'h10 ;
			data[92696] <= 8'h10 ;
			data[92697] <= 8'h10 ;
			data[92698] <= 8'h10 ;
			data[92699] <= 8'h10 ;
			data[92700] <= 8'h10 ;
			data[92701] <= 8'h10 ;
			data[92702] <= 8'h10 ;
			data[92703] <= 8'h10 ;
			data[92704] <= 8'h10 ;
			data[92705] <= 8'h10 ;
			data[92706] <= 8'h10 ;
			data[92707] <= 8'h10 ;
			data[92708] <= 8'h10 ;
			data[92709] <= 8'h10 ;
			data[92710] <= 8'h10 ;
			data[92711] <= 8'h10 ;
			data[92712] <= 8'h10 ;
			data[92713] <= 8'h10 ;
			data[92714] <= 8'h10 ;
			data[92715] <= 8'h10 ;
			data[92716] <= 8'h10 ;
			data[92717] <= 8'h10 ;
			data[92718] <= 8'h10 ;
			data[92719] <= 8'h10 ;
			data[92720] <= 8'h10 ;
			data[92721] <= 8'h10 ;
			data[92722] <= 8'h10 ;
			data[92723] <= 8'h10 ;
			data[92724] <= 8'h10 ;
			data[92725] <= 8'h10 ;
			data[92726] <= 8'h10 ;
			data[92727] <= 8'h10 ;
			data[92728] <= 8'h10 ;
			data[92729] <= 8'h10 ;
			data[92730] <= 8'h10 ;
			data[92731] <= 8'h10 ;
			data[92732] <= 8'h10 ;
			data[92733] <= 8'h10 ;
			data[92734] <= 8'h10 ;
			data[92735] <= 8'h10 ;
			data[92736] <= 8'h10 ;
			data[92737] <= 8'h10 ;
			data[92738] <= 8'h10 ;
			data[92739] <= 8'h10 ;
			data[92740] <= 8'h10 ;
			data[92741] <= 8'h10 ;
			data[92742] <= 8'h10 ;
			data[92743] <= 8'h10 ;
			data[92744] <= 8'h10 ;
			data[92745] <= 8'h10 ;
			data[92746] <= 8'h10 ;
			data[92747] <= 8'h10 ;
			data[92748] <= 8'h10 ;
			data[92749] <= 8'h10 ;
			data[92750] <= 8'h10 ;
			data[92751] <= 8'h10 ;
			data[92752] <= 8'h10 ;
			data[92753] <= 8'h10 ;
			data[92754] <= 8'h10 ;
			data[92755] <= 8'h10 ;
			data[92756] <= 8'h10 ;
			data[92757] <= 8'h10 ;
			data[92758] <= 8'h10 ;
			data[92759] <= 8'h10 ;
			data[92760] <= 8'h10 ;
			data[92761] <= 8'h10 ;
			data[92762] <= 8'h10 ;
			data[92763] <= 8'h10 ;
			data[92764] <= 8'h10 ;
			data[92765] <= 8'h10 ;
			data[92766] <= 8'h10 ;
			data[92767] <= 8'h10 ;
			data[92768] <= 8'h10 ;
			data[92769] <= 8'h10 ;
			data[92770] <= 8'h10 ;
			data[92771] <= 8'h10 ;
			data[92772] <= 8'h10 ;
			data[92773] <= 8'h10 ;
			data[92774] <= 8'h10 ;
			data[92775] <= 8'h10 ;
			data[92776] <= 8'h10 ;
			data[92777] <= 8'h10 ;
			data[92778] <= 8'h10 ;
			data[92779] <= 8'h10 ;
			data[92780] <= 8'h10 ;
			data[92781] <= 8'h10 ;
			data[92782] <= 8'h10 ;
			data[92783] <= 8'h10 ;
			data[92784] <= 8'h10 ;
			data[92785] <= 8'h10 ;
			data[92786] <= 8'h10 ;
			data[92787] <= 8'h10 ;
			data[92788] <= 8'h10 ;
			data[92789] <= 8'h10 ;
			data[92790] <= 8'h10 ;
			data[92791] <= 8'h10 ;
			data[92792] <= 8'h10 ;
			data[92793] <= 8'h10 ;
			data[92794] <= 8'h10 ;
			data[92795] <= 8'h10 ;
			data[92796] <= 8'h10 ;
			data[92797] <= 8'h10 ;
			data[92798] <= 8'h10 ;
			data[92799] <= 8'h10 ;
			data[92800] <= 8'h10 ;
			data[92801] <= 8'h10 ;
			data[92802] <= 8'h10 ;
			data[92803] <= 8'h10 ;
			data[92804] <= 8'h10 ;
			data[92805] <= 8'h10 ;
			data[92806] <= 8'h10 ;
			data[92807] <= 8'h10 ;
			data[92808] <= 8'h10 ;
			data[92809] <= 8'h10 ;
			data[92810] <= 8'h10 ;
			data[92811] <= 8'h10 ;
			data[92812] <= 8'h10 ;
			data[92813] <= 8'h10 ;
			data[92814] <= 8'h10 ;
			data[92815] <= 8'h10 ;
			data[92816] <= 8'h10 ;
			data[92817] <= 8'h10 ;
			data[92818] <= 8'h10 ;
			data[92819] <= 8'h10 ;
			data[92820] <= 8'h10 ;
			data[92821] <= 8'h10 ;
			data[92822] <= 8'h10 ;
			data[92823] <= 8'h10 ;
			data[92824] <= 8'h10 ;
			data[92825] <= 8'h10 ;
			data[92826] <= 8'h10 ;
			data[92827] <= 8'h10 ;
			data[92828] <= 8'h10 ;
			data[92829] <= 8'h10 ;
			data[92830] <= 8'h10 ;
			data[92831] <= 8'h10 ;
			data[92832] <= 8'h10 ;
			data[92833] <= 8'h10 ;
			data[92834] <= 8'h10 ;
			data[92835] <= 8'h10 ;
			data[92836] <= 8'h10 ;
			data[92837] <= 8'h10 ;
			data[92838] <= 8'h10 ;
			data[92839] <= 8'h10 ;
			data[92840] <= 8'h10 ;
			data[92841] <= 8'h10 ;
			data[92842] <= 8'h10 ;
			data[92843] <= 8'h10 ;
			data[92844] <= 8'h10 ;
			data[92845] <= 8'h10 ;
			data[92846] <= 8'h10 ;
			data[92847] <= 8'h10 ;
			data[92848] <= 8'h10 ;
			data[92849] <= 8'h10 ;
			data[92850] <= 8'h10 ;
			data[92851] <= 8'h10 ;
			data[92852] <= 8'h10 ;
			data[92853] <= 8'h10 ;
			data[92854] <= 8'h10 ;
			data[92855] <= 8'h10 ;
			data[92856] <= 8'h10 ;
			data[92857] <= 8'h10 ;
			data[92858] <= 8'h10 ;
			data[92859] <= 8'h10 ;
			data[92860] <= 8'h10 ;
			data[92861] <= 8'h10 ;
			data[92862] <= 8'h10 ;
			data[92863] <= 8'h10 ;
			data[92864] <= 8'h10 ;
			data[92865] <= 8'h10 ;
			data[92866] <= 8'h10 ;
			data[92867] <= 8'h10 ;
			data[92868] <= 8'h10 ;
			data[92869] <= 8'h10 ;
			data[92870] <= 8'h10 ;
			data[92871] <= 8'h10 ;
			data[92872] <= 8'h10 ;
			data[92873] <= 8'h10 ;
			data[92874] <= 8'h10 ;
			data[92875] <= 8'h10 ;
			data[92876] <= 8'h10 ;
			data[92877] <= 8'h10 ;
			data[92878] <= 8'h10 ;
			data[92879] <= 8'h10 ;
			data[92880] <= 8'h10 ;
			data[92881] <= 8'h10 ;
			data[92882] <= 8'h10 ;
			data[92883] <= 8'h10 ;
			data[92884] <= 8'h10 ;
			data[92885] <= 8'h10 ;
			data[92886] <= 8'h10 ;
			data[92887] <= 8'h10 ;
			data[92888] <= 8'h10 ;
			data[92889] <= 8'h10 ;
			data[92890] <= 8'h10 ;
			data[92891] <= 8'h10 ;
			data[92892] <= 8'h10 ;
			data[92893] <= 8'h10 ;
			data[92894] <= 8'h10 ;
			data[92895] <= 8'h10 ;
			data[92896] <= 8'h10 ;
			data[92897] <= 8'h10 ;
			data[92898] <= 8'h10 ;
			data[92899] <= 8'h10 ;
			data[92900] <= 8'h10 ;
			data[92901] <= 8'h10 ;
			data[92902] <= 8'h10 ;
			data[92903] <= 8'h10 ;
			data[92904] <= 8'h10 ;
			data[92905] <= 8'h10 ;
			data[92906] <= 8'h10 ;
			data[92907] <= 8'h10 ;
			data[92908] <= 8'h10 ;
			data[92909] <= 8'h10 ;
			data[92910] <= 8'h10 ;
			data[92911] <= 8'h10 ;
			data[92912] <= 8'h10 ;
			data[92913] <= 8'h10 ;
			data[92914] <= 8'h10 ;
			data[92915] <= 8'h10 ;
			data[92916] <= 8'h10 ;
			data[92917] <= 8'h10 ;
			data[92918] <= 8'h10 ;
			data[92919] <= 8'h10 ;
			data[92920] <= 8'h10 ;
			data[92921] <= 8'h10 ;
			data[92922] <= 8'h10 ;
			data[92923] <= 8'h10 ;
			data[92924] <= 8'h10 ;
			data[92925] <= 8'h10 ;
			data[92926] <= 8'h10 ;
			data[92927] <= 8'h10 ;
			data[92928] <= 8'h10 ;
			data[92929] <= 8'h10 ;
			data[92930] <= 8'h10 ;
			data[92931] <= 8'h10 ;
			data[92932] <= 8'h10 ;
			data[92933] <= 8'h10 ;
			data[92934] <= 8'h10 ;
			data[92935] <= 8'h10 ;
			data[92936] <= 8'h10 ;
			data[92937] <= 8'h10 ;
			data[92938] <= 8'h10 ;
			data[92939] <= 8'h10 ;
			data[92940] <= 8'h10 ;
			data[92941] <= 8'h10 ;
			data[92942] <= 8'h10 ;
			data[92943] <= 8'h10 ;
			data[92944] <= 8'h10 ;
			data[92945] <= 8'h10 ;
			data[92946] <= 8'h10 ;
			data[92947] <= 8'h10 ;
			data[92948] <= 8'h10 ;
			data[92949] <= 8'h10 ;
			data[92950] <= 8'h10 ;
			data[92951] <= 8'h10 ;
			data[92952] <= 8'h10 ;
			data[92953] <= 8'h10 ;
			data[92954] <= 8'h10 ;
			data[92955] <= 8'h10 ;
			data[92956] <= 8'h10 ;
			data[92957] <= 8'h10 ;
			data[92958] <= 8'h10 ;
			data[92959] <= 8'h10 ;
			data[92960] <= 8'h10 ;
			data[92961] <= 8'h10 ;
			data[92962] <= 8'h10 ;
			data[92963] <= 8'h10 ;
			data[92964] <= 8'h10 ;
			data[92965] <= 8'h10 ;
			data[92966] <= 8'h10 ;
			data[92967] <= 8'h10 ;
			data[92968] <= 8'h10 ;
			data[92969] <= 8'h10 ;
			data[92970] <= 8'h10 ;
			data[92971] <= 8'h10 ;
			data[92972] <= 8'h10 ;
			data[92973] <= 8'h10 ;
			data[92974] <= 8'h10 ;
			data[92975] <= 8'h10 ;
			data[92976] <= 8'h10 ;
			data[92977] <= 8'h10 ;
			data[92978] <= 8'h10 ;
			data[92979] <= 8'h10 ;
			data[92980] <= 8'h10 ;
			data[92981] <= 8'h10 ;
			data[92982] <= 8'h10 ;
			data[92983] <= 8'h10 ;
			data[92984] <= 8'h10 ;
			data[92985] <= 8'h10 ;
			data[92986] <= 8'h10 ;
			data[92987] <= 8'h10 ;
			data[92988] <= 8'h10 ;
			data[92989] <= 8'h10 ;
			data[92990] <= 8'h10 ;
			data[92991] <= 8'h10 ;
			data[92992] <= 8'h10 ;
			data[92993] <= 8'h10 ;
			data[92994] <= 8'h10 ;
			data[92995] <= 8'h10 ;
			data[92996] <= 8'h10 ;
			data[92997] <= 8'h10 ;
			data[92998] <= 8'h10 ;
			data[92999] <= 8'h10 ;
			data[93000] <= 8'h10 ;
			data[93001] <= 8'h10 ;
			data[93002] <= 8'h10 ;
			data[93003] <= 8'h10 ;
			data[93004] <= 8'h10 ;
			data[93005] <= 8'h10 ;
			data[93006] <= 8'h10 ;
			data[93007] <= 8'h10 ;
			data[93008] <= 8'h10 ;
			data[93009] <= 8'h10 ;
			data[93010] <= 8'h10 ;
			data[93011] <= 8'h10 ;
			data[93012] <= 8'h10 ;
			data[93013] <= 8'h10 ;
			data[93014] <= 8'h10 ;
			data[93015] <= 8'h10 ;
			data[93016] <= 8'h10 ;
			data[93017] <= 8'h10 ;
			data[93018] <= 8'h10 ;
			data[93019] <= 8'h10 ;
			data[93020] <= 8'h10 ;
			data[93021] <= 8'h10 ;
			data[93022] <= 8'h10 ;
			data[93023] <= 8'h10 ;
			data[93024] <= 8'h10 ;
			data[93025] <= 8'h10 ;
			data[93026] <= 8'h10 ;
			data[93027] <= 8'h10 ;
			data[93028] <= 8'h10 ;
			data[93029] <= 8'h10 ;
			data[93030] <= 8'h10 ;
			data[93031] <= 8'h10 ;
			data[93032] <= 8'h10 ;
			data[93033] <= 8'h10 ;
			data[93034] <= 8'h10 ;
			data[93035] <= 8'h10 ;
			data[93036] <= 8'h10 ;
			data[93037] <= 8'h10 ;
			data[93038] <= 8'h10 ;
			data[93039] <= 8'h10 ;
			data[93040] <= 8'h10 ;
			data[93041] <= 8'h10 ;
			data[93042] <= 8'h10 ;
			data[93043] <= 8'h10 ;
			data[93044] <= 8'h10 ;
			data[93045] <= 8'h10 ;
			data[93046] <= 8'h10 ;
			data[93047] <= 8'h10 ;
			data[93048] <= 8'h10 ;
			data[93049] <= 8'h10 ;
			data[93050] <= 8'h10 ;
			data[93051] <= 8'h10 ;
			data[93052] <= 8'h10 ;
			data[93053] <= 8'h10 ;
			data[93054] <= 8'h10 ;
			data[93055] <= 8'h10 ;
			data[93056] <= 8'h10 ;
			data[93057] <= 8'h10 ;
			data[93058] <= 8'h10 ;
			data[93059] <= 8'h10 ;
			data[93060] <= 8'h10 ;
			data[93061] <= 8'h10 ;
			data[93062] <= 8'h10 ;
			data[93063] <= 8'h10 ;
			data[93064] <= 8'h10 ;
			data[93065] <= 8'h10 ;
			data[93066] <= 8'h10 ;
			data[93067] <= 8'h10 ;
			data[93068] <= 8'h10 ;
			data[93069] <= 8'h10 ;
			data[93070] <= 8'h10 ;
			data[93071] <= 8'h10 ;
			data[93072] <= 8'h10 ;
			data[93073] <= 8'h10 ;
			data[93074] <= 8'h10 ;
			data[93075] <= 8'h10 ;
			data[93076] <= 8'h10 ;
			data[93077] <= 8'h10 ;
			data[93078] <= 8'h10 ;
			data[93079] <= 8'h10 ;
			data[93080] <= 8'h10 ;
			data[93081] <= 8'h10 ;
			data[93082] <= 8'h10 ;
			data[93083] <= 8'h10 ;
			data[93084] <= 8'h10 ;
			data[93085] <= 8'h10 ;
			data[93086] <= 8'h10 ;
			data[93087] <= 8'h10 ;
			data[93088] <= 8'h10 ;
			data[93089] <= 8'h10 ;
			data[93090] <= 8'h10 ;
			data[93091] <= 8'h10 ;
			data[93092] <= 8'h10 ;
			data[93093] <= 8'h10 ;
			data[93094] <= 8'h10 ;
			data[93095] <= 8'h10 ;
			data[93096] <= 8'h10 ;
			data[93097] <= 8'h10 ;
			data[93098] <= 8'h10 ;
			data[93099] <= 8'h10 ;
			data[93100] <= 8'h10 ;
			data[93101] <= 8'h10 ;
			data[93102] <= 8'h10 ;
			data[93103] <= 8'h10 ;
			data[93104] <= 8'h10 ;
			data[93105] <= 8'h10 ;
			data[93106] <= 8'h10 ;
			data[93107] <= 8'h10 ;
			data[93108] <= 8'h10 ;
			data[93109] <= 8'h10 ;
			data[93110] <= 8'h10 ;
			data[93111] <= 8'h10 ;
			data[93112] <= 8'h10 ;
			data[93113] <= 8'h10 ;
			data[93114] <= 8'h10 ;
			data[93115] <= 8'h10 ;
			data[93116] <= 8'h10 ;
			data[93117] <= 8'h10 ;
			data[93118] <= 8'h10 ;
			data[93119] <= 8'h10 ;
			data[93120] <= 8'h10 ;
			data[93121] <= 8'h10 ;
			data[93122] <= 8'h10 ;
			data[93123] <= 8'h10 ;
			data[93124] <= 8'h10 ;
			data[93125] <= 8'h10 ;
			data[93126] <= 8'h10 ;
			data[93127] <= 8'h10 ;
			data[93128] <= 8'h10 ;
			data[93129] <= 8'h10 ;
			data[93130] <= 8'h10 ;
			data[93131] <= 8'h10 ;
			data[93132] <= 8'h10 ;
			data[93133] <= 8'h10 ;
			data[93134] <= 8'h10 ;
			data[93135] <= 8'h10 ;
			data[93136] <= 8'h10 ;
			data[93137] <= 8'h10 ;
			data[93138] <= 8'h10 ;
			data[93139] <= 8'h10 ;
			data[93140] <= 8'h10 ;
			data[93141] <= 8'h10 ;
			data[93142] <= 8'h10 ;
			data[93143] <= 8'h10 ;
			data[93144] <= 8'h10 ;
			data[93145] <= 8'h10 ;
			data[93146] <= 8'h10 ;
			data[93147] <= 8'h10 ;
			data[93148] <= 8'h10 ;
			data[93149] <= 8'h10 ;
			data[93150] <= 8'h10 ;
			data[93151] <= 8'h10 ;
			data[93152] <= 8'h10 ;
			data[93153] <= 8'h10 ;
			data[93154] <= 8'h10 ;
			data[93155] <= 8'h10 ;
			data[93156] <= 8'h10 ;
			data[93157] <= 8'h10 ;
			data[93158] <= 8'h10 ;
			data[93159] <= 8'h10 ;
			data[93160] <= 8'h10 ;
			data[93161] <= 8'h10 ;
			data[93162] <= 8'h10 ;
			data[93163] <= 8'h10 ;
			data[93164] <= 8'h10 ;
			data[93165] <= 8'h10 ;
			data[93166] <= 8'h10 ;
			data[93167] <= 8'h10 ;
			data[93168] <= 8'h10 ;
			data[93169] <= 8'h10 ;
			data[93170] <= 8'h10 ;
			data[93171] <= 8'h10 ;
			data[93172] <= 8'h10 ;
			data[93173] <= 8'h10 ;
			data[93174] <= 8'h10 ;
			data[93175] <= 8'h10 ;
			data[93176] <= 8'h10 ;
			data[93177] <= 8'h10 ;
			data[93178] <= 8'h10 ;
			data[93179] <= 8'h10 ;
			data[93180] <= 8'h10 ;
			data[93181] <= 8'h10 ;
			data[93182] <= 8'h10 ;
			data[93183] <= 8'h10 ;
			data[93184] <= 8'h10 ;
			data[93185] <= 8'h10 ;
			data[93186] <= 8'h10 ;
			data[93187] <= 8'h10 ;
			data[93188] <= 8'h10 ;
			data[93189] <= 8'h10 ;
			data[93190] <= 8'h10 ;
			data[93191] <= 8'h10 ;
			data[93192] <= 8'h10 ;
			data[93193] <= 8'h10 ;
			data[93194] <= 8'h10 ;
			data[93195] <= 8'h10 ;
			data[93196] <= 8'h10 ;
			data[93197] <= 8'h10 ;
			data[93198] <= 8'h10 ;
			data[93199] <= 8'h10 ;
			data[93200] <= 8'h10 ;
			data[93201] <= 8'h10 ;
			data[93202] <= 8'h10 ;
			data[93203] <= 8'h10 ;
			data[93204] <= 8'h10 ;
			data[93205] <= 8'h10 ;
			data[93206] <= 8'h10 ;
			data[93207] <= 8'h10 ;
			data[93208] <= 8'h10 ;
			data[93209] <= 8'h10 ;
			data[93210] <= 8'h10 ;
			data[93211] <= 8'h10 ;
			data[93212] <= 8'h10 ;
			data[93213] <= 8'h10 ;
			data[93214] <= 8'h10 ;
			data[93215] <= 8'h10 ;
			data[93216] <= 8'h10 ;
			data[93217] <= 8'h10 ;
			data[93218] <= 8'h10 ;
			data[93219] <= 8'h10 ;
			data[93220] <= 8'h10 ;
			data[93221] <= 8'h10 ;
			data[93222] <= 8'h10 ;
			data[93223] <= 8'h10 ;
			data[93224] <= 8'h10 ;
			data[93225] <= 8'h10 ;
			data[93226] <= 8'h10 ;
			data[93227] <= 8'h10 ;
			data[93228] <= 8'h10 ;
			data[93229] <= 8'h10 ;
			data[93230] <= 8'h10 ;
			data[93231] <= 8'h10 ;
			data[93232] <= 8'h10 ;
			data[93233] <= 8'h10 ;
			data[93234] <= 8'h10 ;
			data[93235] <= 8'h10 ;
			data[93236] <= 8'h10 ;
			data[93237] <= 8'h10 ;
			data[93238] <= 8'h10 ;
			data[93239] <= 8'h10 ;
			data[93240] <= 8'h10 ;
			data[93241] <= 8'h10 ;
			data[93242] <= 8'h10 ;
			data[93243] <= 8'h10 ;
			data[93244] <= 8'h10 ;
			data[93245] <= 8'h10 ;
			data[93246] <= 8'h10 ;
			data[93247] <= 8'h10 ;
			data[93248] <= 8'h10 ;
			data[93249] <= 8'h10 ;
			data[93250] <= 8'h10 ;
			data[93251] <= 8'h10 ;
			data[93252] <= 8'h10 ;
			data[93253] <= 8'h10 ;
			data[93254] <= 8'h10 ;
			data[93255] <= 8'h10 ;
			data[93256] <= 8'h10 ;
			data[93257] <= 8'h10 ;
			data[93258] <= 8'h10 ;
			data[93259] <= 8'h10 ;
			data[93260] <= 8'h10 ;
			data[93261] <= 8'h10 ;
			data[93262] <= 8'h10 ;
			data[93263] <= 8'h10 ;
			data[93264] <= 8'h10 ;
			data[93265] <= 8'h10 ;
			data[93266] <= 8'h10 ;
			data[93267] <= 8'h10 ;
			data[93268] <= 8'h10 ;
			data[93269] <= 8'h10 ;
			data[93270] <= 8'h10 ;
			data[93271] <= 8'h10 ;
			data[93272] <= 8'h10 ;
			data[93273] <= 8'h10 ;
			data[93274] <= 8'h10 ;
			data[93275] <= 8'h10 ;
			data[93276] <= 8'h10 ;
			data[93277] <= 8'h10 ;
			data[93278] <= 8'h10 ;
			data[93279] <= 8'h10 ;
			data[93280] <= 8'h10 ;
			data[93281] <= 8'h10 ;
			data[93282] <= 8'h10 ;
			data[93283] <= 8'h10 ;
			data[93284] <= 8'h10 ;
			data[93285] <= 8'h10 ;
			data[93286] <= 8'h10 ;
			data[93287] <= 8'h10 ;
			data[93288] <= 8'h10 ;
			data[93289] <= 8'h10 ;
			data[93290] <= 8'h10 ;
			data[93291] <= 8'h10 ;
			data[93292] <= 8'h10 ;
			data[93293] <= 8'h10 ;
			data[93294] <= 8'h10 ;
			data[93295] <= 8'h10 ;
			data[93296] <= 8'h10 ;
			data[93297] <= 8'h10 ;
			data[93298] <= 8'h10 ;
			data[93299] <= 8'h10 ;
			data[93300] <= 8'h10 ;
			data[93301] <= 8'h10 ;
			data[93302] <= 8'h10 ;
			data[93303] <= 8'h10 ;
			data[93304] <= 8'h10 ;
			data[93305] <= 8'h10 ;
			data[93306] <= 8'h10 ;
			data[93307] <= 8'h10 ;
			data[93308] <= 8'h10 ;
			data[93309] <= 8'h10 ;
			data[93310] <= 8'h10 ;
			data[93311] <= 8'h10 ;
			data[93312] <= 8'h10 ;
			data[93313] <= 8'h10 ;
			data[93314] <= 8'h10 ;
			data[93315] <= 8'h10 ;
			data[93316] <= 8'h10 ;
			data[93317] <= 8'h10 ;
			data[93318] <= 8'h10 ;
			data[93319] <= 8'h10 ;
			data[93320] <= 8'h10 ;
			data[93321] <= 8'h10 ;
			data[93322] <= 8'h10 ;
			data[93323] <= 8'h10 ;
			data[93324] <= 8'h10 ;
			data[93325] <= 8'h10 ;
			data[93326] <= 8'h10 ;
			data[93327] <= 8'h10 ;
			data[93328] <= 8'h10 ;
			data[93329] <= 8'h10 ;
			data[93330] <= 8'h10 ;
			data[93331] <= 8'h10 ;
			data[93332] <= 8'h10 ;
			data[93333] <= 8'h10 ;
			data[93334] <= 8'h10 ;
			data[93335] <= 8'h10 ;
			data[93336] <= 8'h10 ;
			data[93337] <= 8'h10 ;
			data[93338] <= 8'h10 ;
			data[93339] <= 8'h10 ;
			data[93340] <= 8'h10 ;
			data[93341] <= 8'h10 ;
			data[93342] <= 8'h10 ;
			data[93343] <= 8'h10 ;
			data[93344] <= 8'h10 ;
			data[93345] <= 8'h10 ;
			data[93346] <= 8'h10 ;
			data[93347] <= 8'h10 ;
			data[93348] <= 8'h10 ;
			data[93349] <= 8'h10 ;
			data[93350] <= 8'h10 ;
			data[93351] <= 8'h10 ;
			data[93352] <= 8'h10 ;
			data[93353] <= 8'h10 ;
			data[93354] <= 8'h10 ;
			data[93355] <= 8'h10 ;
			data[93356] <= 8'h10 ;
			data[93357] <= 8'h10 ;
			data[93358] <= 8'h10 ;
			data[93359] <= 8'h10 ;
			data[93360] <= 8'h10 ;
			data[93361] <= 8'h10 ;
			data[93362] <= 8'h10 ;
			data[93363] <= 8'h10 ;
			data[93364] <= 8'h10 ;
			data[93365] <= 8'h10 ;
			data[93366] <= 8'h10 ;
			data[93367] <= 8'h10 ;
			data[93368] <= 8'h10 ;
			data[93369] <= 8'h10 ;
			data[93370] <= 8'h10 ;
			data[93371] <= 8'h10 ;
			data[93372] <= 8'h10 ;
			data[93373] <= 8'h10 ;
			data[93374] <= 8'h10 ;
			data[93375] <= 8'h10 ;
			data[93376] <= 8'h10 ;
			data[93377] <= 8'h10 ;
			data[93378] <= 8'h10 ;
			data[93379] <= 8'h10 ;
			data[93380] <= 8'h10 ;
			data[93381] <= 8'h10 ;
			data[93382] <= 8'h10 ;
			data[93383] <= 8'h10 ;
			data[93384] <= 8'h10 ;
			data[93385] <= 8'h10 ;
			data[93386] <= 8'h10 ;
			data[93387] <= 8'h10 ;
			data[93388] <= 8'h10 ;
			data[93389] <= 8'h10 ;
			data[93390] <= 8'h10 ;
			data[93391] <= 8'h10 ;
			data[93392] <= 8'h10 ;
			data[93393] <= 8'h10 ;
			data[93394] <= 8'h10 ;
			data[93395] <= 8'h10 ;
			data[93396] <= 8'h10 ;
			data[93397] <= 8'h10 ;
			data[93398] <= 8'h10 ;
			data[93399] <= 8'h10 ;
			data[93400] <= 8'h10 ;
			data[93401] <= 8'h10 ;
			data[93402] <= 8'h10 ;
			data[93403] <= 8'h10 ;
			data[93404] <= 8'h10 ;
			data[93405] <= 8'h10 ;
			data[93406] <= 8'h10 ;
			data[93407] <= 8'h10 ;
			data[93408] <= 8'h10 ;
			data[93409] <= 8'h10 ;
			data[93410] <= 8'h10 ;
			data[93411] <= 8'h10 ;
			data[93412] <= 8'h10 ;
			data[93413] <= 8'h10 ;
			data[93414] <= 8'h10 ;
			data[93415] <= 8'h10 ;
			data[93416] <= 8'h10 ;
			data[93417] <= 8'h10 ;
			data[93418] <= 8'h10 ;
			data[93419] <= 8'h10 ;
			data[93420] <= 8'h10 ;
			data[93421] <= 8'h10 ;
			data[93422] <= 8'h10 ;
			data[93423] <= 8'h10 ;
			data[93424] <= 8'h10 ;
			data[93425] <= 8'h10 ;
			data[93426] <= 8'h10 ;
			data[93427] <= 8'h10 ;
			data[93428] <= 8'h10 ;
			data[93429] <= 8'h10 ;
			data[93430] <= 8'h10 ;
			data[93431] <= 8'h10 ;
			data[93432] <= 8'h10 ;
			data[93433] <= 8'h10 ;
			data[93434] <= 8'h10 ;
			data[93435] <= 8'h10 ;
			data[93436] <= 8'h10 ;
			data[93437] <= 8'h10 ;
			data[93438] <= 8'h10 ;
			data[93439] <= 8'h10 ;
			data[93440] <= 8'h10 ;
			data[93441] <= 8'h10 ;
			data[93442] <= 8'h10 ;
			data[93443] <= 8'h10 ;
			data[93444] <= 8'h10 ;
			data[93445] <= 8'h10 ;
			data[93446] <= 8'h10 ;
			data[93447] <= 8'h10 ;
			data[93448] <= 8'h10 ;
			data[93449] <= 8'h10 ;
			data[93450] <= 8'h10 ;
			data[93451] <= 8'h10 ;
			data[93452] <= 8'h10 ;
			data[93453] <= 8'h10 ;
			data[93454] <= 8'h10 ;
			data[93455] <= 8'h10 ;
			data[93456] <= 8'h10 ;
			data[93457] <= 8'h10 ;
			data[93458] <= 8'h10 ;
			data[93459] <= 8'h10 ;
			data[93460] <= 8'h10 ;
			data[93461] <= 8'h10 ;
			data[93462] <= 8'h10 ;
			data[93463] <= 8'h10 ;
			data[93464] <= 8'h10 ;
			data[93465] <= 8'h10 ;
			data[93466] <= 8'h10 ;
			data[93467] <= 8'h10 ;
			data[93468] <= 8'h10 ;
			data[93469] <= 8'h10 ;
			data[93470] <= 8'h10 ;
			data[93471] <= 8'h10 ;
			data[93472] <= 8'h10 ;
			data[93473] <= 8'h10 ;
			data[93474] <= 8'h10 ;
			data[93475] <= 8'h10 ;
			data[93476] <= 8'h10 ;
			data[93477] <= 8'h10 ;
			data[93478] <= 8'h10 ;
			data[93479] <= 8'h10 ;
			data[93480] <= 8'h10 ;
			data[93481] <= 8'h10 ;
			data[93482] <= 8'h10 ;
			data[93483] <= 8'h10 ;
			data[93484] <= 8'h10 ;
			data[93485] <= 8'h10 ;
			data[93486] <= 8'h10 ;
			data[93487] <= 8'h10 ;
			data[93488] <= 8'h10 ;
			data[93489] <= 8'h10 ;
			data[93490] <= 8'h10 ;
			data[93491] <= 8'h10 ;
			data[93492] <= 8'h10 ;
			data[93493] <= 8'h10 ;
			data[93494] <= 8'h10 ;
			data[93495] <= 8'h10 ;
			data[93496] <= 8'h10 ;
			data[93497] <= 8'h10 ;
			data[93498] <= 8'h10 ;
			data[93499] <= 8'h10 ;
			data[93500] <= 8'h10 ;
			data[93501] <= 8'h10 ;
			data[93502] <= 8'h10 ;
			data[93503] <= 8'h10 ;
			data[93504] <= 8'h10 ;
			data[93505] <= 8'h10 ;
			data[93506] <= 8'h10 ;
			data[93507] <= 8'h10 ;
			data[93508] <= 8'h10 ;
			data[93509] <= 8'h10 ;
			data[93510] <= 8'h10 ;
			data[93511] <= 8'h10 ;
			data[93512] <= 8'h10 ;
			data[93513] <= 8'h10 ;
			data[93514] <= 8'h10 ;
			data[93515] <= 8'h10 ;
			data[93516] <= 8'h10 ;
			data[93517] <= 8'h10 ;
			data[93518] <= 8'h10 ;
			data[93519] <= 8'h10 ;
			data[93520] <= 8'h10 ;
			data[93521] <= 8'h10 ;
			data[93522] <= 8'h10 ;
			data[93523] <= 8'h10 ;
			data[93524] <= 8'h10 ;
			data[93525] <= 8'h10 ;
			data[93526] <= 8'h10 ;
			data[93527] <= 8'h10 ;
			data[93528] <= 8'h10 ;
			data[93529] <= 8'h10 ;
			data[93530] <= 8'h10 ;
			data[93531] <= 8'h10 ;
			data[93532] <= 8'h10 ;
			data[93533] <= 8'h10 ;
			data[93534] <= 8'h10 ;
			data[93535] <= 8'h10 ;
			data[93536] <= 8'h10 ;
			data[93537] <= 8'h10 ;
			data[93538] <= 8'h10 ;
			data[93539] <= 8'h10 ;
			data[93540] <= 8'h10 ;
			data[93541] <= 8'h10 ;
			data[93542] <= 8'h10 ;
			data[93543] <= 8'h10 ;
			data[93544] <= 8'h10 ;
			data[93545] <= 8'h10 ;
			data[93546] <= 8'h10 ;
			data[93547] <= 8'h10 ;
			data[93548] <= 8'h10 ;
			data[93549] <= 8'h10 ;
			data[93550] <= 8'h10 ;
			data[93551] <= 8'h10 ;
			data[93552] <= 8'h10 ;
			data[93553] <= 8'h10 ;
			data[93554] <= 8'h10 ;
			data[93555] <= 8'h10 ;
			data[93556] <= 8'h10 ;
			data[93557] <= 8'h10 ;
			data[93558] <= 8'h10 ;
			data[93559] <= 8'h10 ;
			data[93560] <= 8'h10 ;
			data[93561] <= 8'h10 ;
			data[93562] <= 8'h10 ;
			data[93563] <= 8'h10 ;
			data[93564] <= 8'h10 ;
			data[93565] <= 8'h10 ;
			data[93566] <= 8'h10 ;
			data[93567] <= 8'h10 ;
			data[93568] <= 8'h10 ;
			data[93569] <= 8'h10 ;
			data[93570] <= 8'h10 ;
			data[93571] <= 8'h10 ;
			data[93572] <= 8'h10 ;
			data[93573] <= 8'h10 ;
			data[93574] <= 8'h10 ;
			data[93575] <= 8'h10 ;
			data[93576] <= 8'h10 ;
			data[93577] <= 8'h10 ;
			data[93578] <= 8'h10 ;
			data[93579] <= 8'h10 ;
			data[93580] <= 8'h10 ;
			data[93581] <= 8'h10 ;
			data[93582] <= 8'h10 ;
			data[93583] <= 8'h10 ;
			data[93584] <= 8'h10 ;
			data[93585] <= 8'h10 ;
			data[93586] <= 8'h10 ;
			data[93587] <= 8'h10 ;
			data[93588] <= 8'h10 ;
			data[93589] <= 8'h10 ;
			data[93590] <= 8'h10 ;
			data[93591] <= 8'h10 ;
			data[93592] <= 8'h10 ;
			data[93593] <= 8'h10 ;
			data[93594] <= 8'h10 ;
			data[93595] <= 8'h10 ;
			data[93596] <= 8'h10 ;
			data[93597] <= 8'h10 ;
			data[93598] <= 8'h10 ;
			data[93599] <= 8'h10 ;
			data[93600] <= 8'h10 ;
			data[93601] <= 8'h10 ;
			data[93602] <= 8'h10 ;
			data[93603] <= 8'h10 ;
			data[93604] <= 8'h10 ;
			data[93605] <= 8'h10 ;
			data[93606] <= 8'h10 ;
			data[93607] <= 8'h10 ;
			data[93608] <= 8'h10 ;
			data[93609] <= 8'h10 ;
			data[93610] <= 8'h10 ;
			data[93611] <= 8'h10 ;
			data[93612] <= 8'h10 ;
			data[93613] <= 8'h10 ;
			data[93614] <= 8'h10 ;
			data[93615] <= 8'h10 ;
			data[93616] <= 8'h10 ;
			data[93617] <= 8'h10 ;
			data[93618] <= 8'h10 ;
			data[93619] <= 8'h10 ;
			data[93620] <= 8'h10 ;
			data[93621] <= 8'h10 ;
			data[93622] <= 8'h10 ;
			data[93623] <= 8'h10 ;
			data[93624] <= 8'h10 ;
			data[93625] <= 8'h10 ;
			data[93626] <= 8'h10 ;
			data[93627] <= 8'h10 ;
			data[93628] <= 8'h10 ;
			data[93629] <= 8'h10 ;
			data[93630] <= 8'h10 ;
			data[93631] <= 8'h10 ;
			data[93632] <= 8'h10 ;
			data[93633] <= 8'h10 ;
			data[93634] <= 8'h10 ;
			data[93635] <= 8'h10 ;
			data[93636] <= 8'h10 ;
			data[93637] <= 8'h10 ;
			data[93638] <= 8'h10 ;
			data[93639] <= 8'h10 ;
			data[93640] <= 8'h10 ;
			data[93641] <= 8'h10 ;
			data[93642] <= 8'h10 ;
			data[93643] <= 8'h10 ;
			data[93644] <= 8'h10 ;
			data[93645] <= 8'h10 ;
			data[93646] <= 8'h10 ;
			data[93647] <= 8'h10 ;
			data[93648] <= 8'h10 ;
			data[93649] <= 8'h10 ;
			data[93650] <= 8'h10 ;
			data[93651] <= 8'h10 ;
			data[93652] <= 8'h10 ;
			data[93653] <= 8'h10 ;
			data[93654] <= 8'h10 ;
			data[93655] <= 8'h10 ;
			data[93656] <= 8'h10 ;
			data[93657] <= 8'h10 ;
			data[93658] <= 8'h10 ;
			data[93659] <= 8'h10 ;
			data[93660] <= 8'h10 ;
			data[93661] <= 8'h10 ;
			data[93662] <= 8'h10 ;
			data[93663] <= 8'h10 ;
			data[93664] <= 8'h10 ;
			data[93665] <= 8'h10 ;
			data[93666] <= 8'h10 ;
			data[93667] <= 8'h10 ;
			data[93668] <= 8'h10 ;
			data[93669] <= 8'h10 ;
			data[93670] <= 8'h10 ;
			data[93671] <= 8'h10 ;
			data[93672] <= 8'h10 ;
			data[93673] <= 8'h10 ;
			data[93674] <= 8'h10 ;
			data[93675] <= 8'h10 ;
			data[93676] <= 8'h10 ;
			data[93677] <= 8'h10 ;
			data[93678] <= 8'h10 ;
			data[93679] <= 8'h10 ;
			data[93680] <= 8'h10 ;
			data[93681] <= 8'h10 ;
			data[93682] <= 8'h10 ;
			data[93683] <= 8'h10 ;
			data[93684] <= 8'h10 ;
			data[93685] <= 8'h10 ;
			data[93686] <= 8'h10 ;
			data[93687] <= 8'h10 ;
			data[93688] <= 8'h10 ;
			data[93689] <= 8'h10 ;
			data[93690] <= 8'h10 ;
			data[93691] <= 8'h10 ;
			data[93692] <= 8'h10 ;
			data[93693] <= 8'h10 ;
			data[93694] <= 8'h10 ;
			data[93695] <= 8'h10 ;
			data[93696] <= 8'h10 ;
			data[93697] <= 8'h10 ;
			data[93698] <= 8'h10 ;
			data[93699] <= 8'h10 ;
			data[93700] <= 8'h10 ;
			data[93701] <= 8'h10 ;
			data[93702] <= 8'h10 ;
			data[93703] <= 8'h10 ;
			data[93704] <= 8'h10 ;
			data[93705] <= 8'h10 ;
			data[93706] <= 8'h10 ;
			data[93707] <= 8'h10 ;
			data[93708] <= 8'h10 ;
			data[93709] <= 8'h10 ;
			data[93710] <= 8'h10 ;
			data[93711] <= 8'h10 ;
			data[93712] <= 8'h10 ;
			data[93713] <= 8'h10 ;
			data[93714] <= 8'h10 ;
			data[93715] <= 8'h10 ;
			data[93716] <= 8'h10 ;
			data[93717] <= 8'h10 ;
			data[93718] <= 8'h10 ;
			data[93719] <= 8'h10 ;
			data[93720] <= 8'h10 ;
			data[93721] <= 8'h10 ;
			data[93722] <= 8'h10 ;
			data[93723] <= 8'h10 ;
			data[93724] <= 8'h10 ;
			data[93725] <= 8'h10 ;
			data[93726] <= 8'h10 ;
			data[93727] <= 8'h10 ;
			data[93728] <= 8'h10 ;
			data[93729] <= 8'h10 ;
			data[93730] <= 8'h10 ;
			data[93731] <= 8'h10 ;
			data[93732] <= 8'h10 ;
			data[93733] <= 8'h10 ;
			data[93734] <= 8'h10 ;
			data[93735] <= 8'h10 ;
			data[93736] <= 8'h10 ;
			data[93737] <= 8'h10 ;
			data[93738] <= 8'h10 ;
			data[93739] <= 8'h10 ;
			data[93740] <= 8'h10 ;
			data[93741] <= 8'h10 ;
			data[93742] <= 8'h10 ;
			data[93743] <= 8'h10 ;
			data[93744] <= 8'h10 ;
			data[93745] <= 8'h10 ;
			data[93746] <= 8'h10 ;
			data[93747] <= 8'h10 ;
			data[93748] <= 8'h10 ;
			data[93749] <= 8'h10 ;
			data[93750] <= 8'h10 ;
			data[93751] <= 8'h10 ;
			data[93752] <= 8'h10 ;
			data[93753] <= 8'h10 ;
			data[93754] <= 8'h10 ;
			data[93755] <= 8'h10 ;
			data[93756] <= 8'h10 ;
			data[93757] <= 8'h10 ;
			data[93758] <= 8'h10 ;
			data[93759] <= 8'h10 ;
			data[93760] <= 8'h10 ;
			data[93761] <= 8'h10 ;
			data[93762] <= 8'h10 ;
			data[93763] <= 8'h10 ;
			data[93764] <= 8'h10 ;
			data[93765] <= 8'h10 ;
			data[93766] <= 8'h10 ;
			data[93767] <= 8'h10 ;
			data[93768] <= 8'h10 ;
			data[93769] <= 8'h10 ;
			data[93770] <= 8'h10 ;
			data[93771] <= 8'h10 ;
			data[93772] <= 8'h10 ;
			data[93773] <= 8'h10 ;
			data[93774] <= 8'h10 ;
			data[93775] <= 8'h10 ;
			data[93776] <= 8'h10 ;
			data[93777] <= 8'h10 ;
			data[93778] <= 8'h10 ;
			data[93779] <= 8'h10 ;
			data[93780] <= 8'h10 ;
			data[93781] <= 8'h10 ;
			data[93782] <= 8'h10 ;
			data[93783] <= 8'h10 ;
			data[93784] <= 8'h10 ;
			data[93785] <= 8'h10 ;
			data[93786] <= 8'h10 ;
			data[93787] <= 8'h10 ;
			data[93788] <= 8'h10 ;
			data[93789] <= 8'h10 ;
			data[93790] <= 8'h10 ;
			data[93791] <= 8'h10 ;
			data[93792] <= 8'h10 ;
			data[93793] <= 8'h10 ;
			data[93794] <= 8'h10 ;
			data[93795] <= 8'h10 ;
			data[93796] <= 8'h10 ;
			data[93797] <= 8'h10 ;
			data[93798] <= 8'h10 ;
			data[93799] <= 8'h10 ;
			data[93800] <= 8'h10 ;
			data[93801] <= 8'h10 ;
			data[93802] <= 8'h10 ;
			data[93803] <= 8'h10 ;
			data[93804] <= 8'h10 ;
			data[93805] <= 8'h10 ;
			data[93806] <= 8'h10 ;
			data[93807] <= 8'h10 ;
			data[93808] <= 8'h10 ;
			data[93809] <= 8'h10 ;
			data[93810] <= 8'h10 ;
			data[93811] <= 8'h10 ;
			data[93812] <= 8'h10 ;
			data[93813] <= 8'h10 ;
			data[93814] <= 8'h10 ;
			data[93815] <= 8'h10 ;
			data[93816] <= 8'h10 ;
			data[93817] <= 8'h10 ;
			data[93818] <= 8'h10 ;
			data[93819] <= 8'h10 ;
			data[93820] <= 8'h10 ;
			data[93821] <= 8'h10 ;
			data[93822] <= 8'h10 ;
			data[93823] <= 8'h10 ;
			data[93824] <= 8'h10 ;
			data[93825] <= 8'h10 ;
			data[93826] <= 8'h10 ;
			data[93827] <= 8'h10 ;
			data[93828] <= 8'h10 ;
			data[93829] <= 8'h10 ;
			data[93830] <= 8'h10 ;
			data[93831] <= 8'h10 ;
			data[93832] <= 8'h10 ;
			data[93833] <= 8'h10 ;
			data[93834] <= 8'h10 ;
			data[93835] <= 8'h10 ;
			data[93836] <= 8'h10 ;
			data[93837] <= 8'h10 ;
			data[93838] <= 8'h10 ;
			data[93839] <= 8'h10 ;
			data[93840] <= 8'h10 ;
			data[93841] <= 8'h10 ;
			data[93842] <= 8'h10 ;
			data[93843] <= 8'h10 ;
			data[93844] <= 8'h10 ;
			data[93845] <= 8'h10 ;
			data[93846] <= 8'h10 ;
			data[93847] <= 8'h10 ;
			data[93848] <= 8'h10 ;
			data[93849] <= 8'h10 ;
			data[93850] <= 8'h10 ;
			data[93851] <= 8'h10 ;
			data[93852] <= 8'h10 ;
			data[93853] <= 8'h10 ;
			data[93854] <= 8'h10 ;
			data[93855] <= 8'h10 ;
			data[93856] <= 8'h10 ;
			data[93857] <= 8'h10 ;
			data[93858] <= 8'h10 ;
			data[93859] <= 8'h10 ;
			data[93860] <= 8'h10 ;
			data[93861] <= 8'h10 ;
			data[93862] <= 8'h10 ;
			data[93863] <= 8'h10 ;
			data[93864] <= 8'h10 ;
			data[93865] <= 8'h10 ;
			data[93866] <= 8'h10 ;
			data[93867] <= 8'h10 ;
			data[93868] <= 8'h10 ;
			data[93869] <= 8'h10 ;
			data[93870] <= 8'h10 ;
			data[93871] <= 8'h10 ;
			data[93872] <= 8'h10 ;
			data[93873] <= 8'h10 ;
			data[93874] <= 8'h10 ;
			data[93875] <= 8'h10 ;
			data[93876] <= 8'h10 ;
			data[93877] <= 8'h10 ;
			data[93878] <= 8'h10 ;
			data[93879] <= 8'h10 ;
			data[93880] <= 8'h10 ;
			data[93881] <= 8'h10 ;
			data[93882] <= 8'h10 ;
			data[93883] <= 8'h10 ;
			data[93884] <= 8'h10 ;
			data[93885] <= 8'h10 ;
			data[93886] <= 8'h10 ;
			data[93887] <= 8'h10 ;
			data[93888] <= 8'h10 ;
			data[93889] <= 8'h10 ;
			data[93890] <= 8'h10 ;
			data[93891] <= 8'h10 ;
			data[93892] <= 8'h10 ;
			data[93893] <= 8'h10 ;
			data[93894] <= 8'h10 ;
			data[93895] <= 8'h10 ;
			data[93896] <= 8'h10 ;
			data[93897] <= 8'h10 ;
			data[93898] <= 8'h10 ;
			data[93899] <= 8'h10 ;
			data[93900] <= 8'h10 ;
			data[93901] <= 8'h10 ;
			data[93902] <= 8'h10 ;
			data[93903] <= 8'h10 ;
			data[93904] <= 8'h10 ;
			data[93905] <= 8'h10 ;
			data[93906] <= 8'h10 ;
			data[93907] <= 8'h10 ;
			data[93908] <= 8'h10 ;
			data[93909] <= 8'h10 ;
			data[93910] <= 8'h10 ;
			data[93911] <= 8'h10 ;
			data[93912] <= 8'h10 ;
			data[93913] <= 8'h10 ;
			data[93914] <= 8'h10 ;
			data[93915] <= 8'h10 ;
			data[93916] <= 8'h10 ;
			data[93917] <= 8'h10 ;
			data[93918] <= 8'h10 ;
			data[93919] <= 8'h10 ;
			data[93920] <= 8'h10 ;
			data[93921] <= 8'h10 ;
			data[93922] <= 8'h10 ;
			data[93923] <= 8'h10 ;
			data[93924] <= 8'h10 ;
			data[93925] <= 8'h10 ;
			data[93926] <= 8'h10 ;
			data[93927] <= 8'h10 ;
			data[93928] <= 8'h10 ;
			data[93929] <= 8'h10 ;
			data[93930] <= 8'h10 ;
			data[93931] <= 8'h10 ;
			data[93932] <= 8'h10 ;
			data[93933] <= 8'h10 ;
			data[93934] <= 8'h10 ;
			data[93935] <= 8'h10 ;
			data[93936] <= 8'h10 ;
			data[93937] <= 8'h10 ;
			data[93938] <= 8'h10 ;
			data[93939] <= 8'h10 ;
			data[93940] <= 8'h10 ;
			data[93941] <= 8'h10 ;
			data[93942] <= 8'h10 ;
			data[93943] <= 8'h10 ;
			data[93944] <= 8'h10 ;
			data[93945] <= 8'h10 ;
			data[93946] <= 8'h10 ;
			data[93947] <= 8'h10 ;
			data[93948] <= 8'h10 ;
			data[93949] <= 8'h10 ;
			data[93950] <= 8'h10 ;
			data[93951] <= 8'h10 ;
			data[93952] <= 8'h10 ;
			data[93953] <= 8'h10 ;
			data[93954] <= 8'h10 ;
			data[93955] <= 8'h10 ;
			data[93956] <= 8'h10 ;
			data[93957] <= 8'h10 ;
			data[93958] <= 8'h10 ;
			data[93959] <= 8'h10 ;
			data[93960] <= 8'h10 ;
			data[93961] <= 8'h10 ;
			data[93962] <= 8'h10 ;
			data[93963] <= 8'h10 ;
			data[93964] <= 8'h10 ;
			data[93965] <= 8'h10 ;
			data[93966] <= 8'h10 ;
			data[93967] <= 8'h10 ;
			data[93968] <= 8'h10 ;
			data[93969] <= 8'h10 ;
			data[93970] <= 8'h10 ;
			data[93971] <= 8'h10 ;
			data[93972] <= 8'h10 ;
			data[93973] <= 8'h10 ;
			data[93974] <= 8'h10 ;
			data[93975] <= 8'h10 ;
			data[93976] <= 8'h10 ;
			data[93977] <= 8'h10 ;
			data[93978] <= 8'h10 ;
			data[93979] <= 8'h10 ;
			data[93980] <= 8'h10 ;
			data[93981] <= 8'h10 ;
			data[93982] <= 8'h10 ;
			data[93983] <= 8'h10 ;
			data[93984] <= 8'h10 ;
			data[93985] <= 8'h10 ;
			data[93986] <= 8'h10 ;
			data[93987] <= 8'h10 ;
			data[93988] <= 8'h10 ;
			data[93989] <= 8'h10 ;
			data[93990] <= 8'h10 ;
			data[93991] <= 8'h10 ;
			data[93992] <= 8'h10 ;
			data[93993] <= 8'h10 ;
			data[93994] <= 8'h10 ;
			data[93995] <= 8'h10 ;
			data[93996] <= 8'h10 ;
			data[93997] <= 8'h10 ;
			data[93998] <= 8'h10 ;
			data[93999] <= 8'h10 ;
			data[94000] <= 8'h10 ;
			data[94001] <= 8'h10 ;
			data[94002] <= 8'h10 ;
			data[94003] <= 8'h10 ;
			data[94004] <= 8'h10 ;
			data[94005] <= 8'h10 ;
			data[94006] <= 8'h10 ;
			data[94007] <= 8'h10 ;
			data[94008] <= 8'h10 ;
			data[94009] <= 8'h10 ;
			data[94010] <= 8'h10 ;
			data[94011] <= 8'h10 ;
			data[94012] <= 8'h10 ;
			data[94013] <= 8'h10 ;
			data[94014] <= 8'h10 ;
			data[94015] <= 8'h10 ;
			data[94016] <= 8'h10 ;
			data[94017] <= 8'h10 ;
			data[94018] <= 8'h10 ;
			data[94019] <= 8'h10 ;
			data[94020] <= 8'h10 ;
			data[94021] <= 8'h10 ;
			data[94022] <= 8'h10 ;
			data[94023] <= 8'h10 ;
			data[94024] <= 8'h10 ;
			data[94025] <= 8'h10 ;
			data[94026] <= 8'h10 ;
			data[94027] <= 8'h10 ;
			data[94028] <= 8'h10 ;
			data[94029] <= 8'h10 ;
			data[94030] <= 8'h10 ;
			data[94031] <= 8'h10 ;
			data[94032] <= 8'h10 ;
			data[94033] <= 8'h10 ;
			data[94034] <= 8'h10 ;
			data[94035] <= 8'h10 ;
			data[94036] <= 8'h10 ;
			data[94037] <= 8'h10 ;
			data[94038] <= 8'h10 ;
			data[94039] <= 8'h10 ;
			data[94040] <= 8'h10 ;
			data[94041] <= 8'h10 ;
			data[94042] <= 8'h10 ;
			data[94043] <= 8'h10 ;
			data[94044] <= 8'h10 ;
			data[94045] <= 8'h10 ;
			data[94046] <= 8'h10 ;
			data[94047] <= 8'h10 ;
			data[94048] <= 8'h10 ;
			data[94049] <= 8'h10 ;
			data[94050] <= 8'h10 ;
			data[94051] <= 8'h10 ;
			data[94052] <= 8'h10 ;
			data[94053] <= 8'h10 ;
			data[94054] <= 8'h10 ;
			data[94055] <= 8'h10 ;
			data[94056] <= 8'h10 ;
			data[94057] <= 8'h10 ;
			data[94058] <= 8'h10 ;
			data[94059] <= 8'h10 ;
			data[94060] <= 8'h10 ;
			data[94061] <= 8'h10 ;
			data[94062] <= 8'h10 ;
			data[94063] <= 8'h10 ;
			data[94064] <= 8'h10 ;
			data[94065] <= 8'h10 ;
			data[94066] <= 8'h10 ;
			data[94067] <= 8'h10 ;
			data[94068] <= 8'h10 ;
			data[94069] <= 8'h10 ;
			data[94070] <= 8'h10 ;
			data[94071] <= 8'h10 ;
			data[94072] <= 8'h10 ;
			data[94073] <= 8'h10 ;
			data[94074] <= 8'h10 ;
			data[94075] <= 8'h10 ;
			data[94076] <= 8'h10 ;
			data[94077] <= 8'h10 ;
			data[94078] <= 8'h10 ;
			data[94079] <= 8'h10 ;
			data[94080] <= 8'h10 ;
			data[94081] <= 8'h10 ;
			data[94082] <= 8'h10 ;
			data[94083] <= 8'h10 ;
			data[94084] <= 8'h10 ;
			data[94085] <= 8'h10 ;
			data[94086] <= 8'h10 ;
			data[94087] <= 8'h10 ;
			data[94088] <= 8'h10 ;
			data[94089] <= 8'h10 ;
			data[94090] <= 8'h10 ;
			data[94091] <= 8'h10 ;
			data[94092] <= 8'h10 ;
			data[94093] <= 8'h10 ;
			data[94094] <= 8'h10 ;
			data[94095] <= 8'h10 ;
			data[94096] <= 8'h10 ;
			data[94097] <= 8'h10 ;
			data[94098] <= 8'h10 ;
			data[94099] <= 8'h10 ;
			data[94100] <= 8'h10 ;
			data[94101] <= 8'h10 ;
			data[94102] <= 8'h10 ;
			data[94103] <= 8'h10 ;
			data[94104] <= 8'h10 ;
			data[94105] <= 8'h10 ;
			data[94106] <= 8'h10 ;
			data[94107] <= 8'h10 ;
			data[94108] <= 8'h10 ;
			data[94109] <= 8'h10 ;
			data[94110] <= 8'h10 ;
			data[94111] <= 8'h10 ;
			data[94112] <= 8'h10 ;
			data[94113] <= 8'h10 ;
			data[94114] <= 8'h10 ;
			data[94115] <= 8'h10 ;
			data[94116] <= 8'h10 ;
			data[94117] <= 8'h10 ;
			data[94118] <= 8'h10 ;
			data[94119] <= 8'h10 ;
			data[94120] <= 8'h10 ;
			data[94121] <= 8'h10 ;
			data[94122] <= 8'h10 ;
			data[94123] <= 8'h10 ;
			data[94124] <= 8'h10 ;
			data[94125] <= 8'h10 ;
			data[94126] <= 8'h10 ;
			data[94127] <= 8'h10 ;
			data[94128] <= 8'h10 ;
			data[94129] <= 8'h10 ;
			data[94130] <= 8'h10 ;
			data[94131] <= 8'h10 ;
			data[94132] <= 8'h10 ;
			data[94133] <= 8'h10 ;
			data[94134] <= 8'h10 ;
			data[94135] <= 8'h10 ;
			data[94136] <= 8'h10 ;
			data[94137] <= 8'h10 ;
			data[94138] <= 8'h10 ;
			data[94139] <= 8'h10 ;
			data[94140] <= 8'h10 ;
			data[94141] <= 8'h10 ;
			data[94142] <= 8'h10 ;
			data[94143] <= 8'h10 ;
			data[94144] <= 8'h10 ;
			data[94145] <= 8'h10 ;
			data[94146] <= 8'h10 ;
			data[94147] <= 8'h10 ;
			data[94148] <= 8'h10 ;
			data[94149] <= 8'h10 ;
			data[94150] <= 8'h10 ;
			data[94151] <= 8'h10 ;
			data[94152] <= 8'h10 ;
			data[94153] <= 8'h10 ;
			data[94154] <= 8'h10 ;
			data[94155] <= 8'h10 ;
			data[94156] <= 8'h10 ;
			data[94157] <= 8'h10 ;
			data[94158] <= 8'h10 ;
			data[94159] <= 8'h10 ;
			data[94160] <= 8'h10 ;
			data[94161] <= 8'h10 ;
			data[94162] <= 8'h10 ;
			data[94163] <= 8'h10 ;
			data[94164] <= 8'h10 ;
			data[94165] <= 8'h10 ;
			data[94166] <= 8'h10 ;
			data[94167] <= 8'h10 ;
			data[94168] <= 8'h10 ;
			data[94169] <= 8'h10 ;
			data[94170] <= 8'h10 ;
			data[94171] <= 8'h10 ;
			data[94172] <= 8'h10 ;
			data[94173] <= 8'h10 ;
			data[94174] <= 8'h10 ;
			data[94175] <= 8'h10 ;
			data[94176] <= 8'h10 ;
			data[94177] <= 8'h10 ;
			data[94178] <= 8'h10 ;
			data[94179] <= 8'h10 ;
			data[94180] <= 8'h10 ;
			data[94181] <= 8'h10 ;
			data[94182] <= 8'h10 ;
			data[94183] <= 8'h10 ;
			data[94184] <= 8'h10 ;
			data[94185] <= 8'h10 ;
			data[94186] <= 8'h10 ;
			data[94187] <= 8'h10 ;
			data[94188] <= 8'h10 ;
			data[94189] <= 8'h10 ;
			data[94190] <= 8'h10 ;
			data[94191] <= 8'h10 ;
			data[94192] <= 8'h10 ;
			data[94193] <= 8'h10 ;
			data[94194] <= 8'h10 ;
			data[94195] <= 8'h10 ;
			data[94196] <= 8'h10 ;
			data[94197] <= 8'h10 ;
			data[94198] <= 8'h10 ;
			data[94199] <= 8'h10 ;
			data[94200] <= 8'h10 ;
			data[94201] <= 8'h10 ;
			data[94202] <= 8'h10 ;
			data[94203] <= 8'h10 ;
			data[94204] <= 8'h10 ;
			data[94205] <= 8'h10 ;
			data[94206] <= 8'h10 ;
			data[94207] <= 8'h10 ;
			data[94208] <= 8'h10 ;
			data[94209] <= 8'h10 ;
			data[94210] <= 8'h10 ;
			data[94211] <= 8'h10 ;
			data[94212] <= 8'h10 ;
			data[94213] <= 8'h10 ;
			data[94214] <= 8'h10 ;
			data[94215] <= 8'h10 ;
			data[94216] <= 8'h10 ;
			data[94217] <= 8'h10 ;
			data[94218] <= 8'h10 ;
			data[94219] <= 8'h10 ;
			data[94220] <= 8'h10 ;
			data[94221] <= 8'h10 ;
			data[94222] <= 8'h10 ;
			data[94223] <= 8'h10 ;
			data[94224] <= 8'h10 ;
			data[94225] <= 8'h10 ;
			data[94226] <= 8'h10 ;
			data[94227] <= 8'h10 ;
			data[94228] <= 8'h10 ;
			data[94229] <= 8'h10 ;
			data[94230] <= 8'h10 ;
			data[94231] <= 8'h10 ;
			data[94232] <= 8'h10 ;
			data[94233] <= 8'h10 ;
			data[94234] <= 8'h10 ;
			data[94235] <= 8'h10 ;
			data[94236] <= 8'h10 ;
			data[94237] <= 8'h10 ;
			data[94238] <= 8'h10 ;
			data[94239] <= 8'h10 ;
			data[94240] <= 8'h10 ;
			data[94241] <= 8'h10 ;
			data[94242] <= 8'h10 ;
			data[94243] <= 8'h10 ;
			data[94244] <= 8'h10 ;
			data[94245] <= 8'h10 ;
			data[94246] <= 8'h10 ;
			data[94247] <= 8'h10 ;
			data[94248] <= 8'h10 ;
			data[94249] <= 8'h10 ;
			data[94250] <= 8'h10 ;
			data[94251] <= 8'h10 ;
			data[94252] <= 8'h10 ;
			data[94253] <= 8'h10 ;
			data[94254] <= 8'h10 ;
			data[94255] <= 8'h10 ;
			data[94256] <= 8'h10 ;
			data[94257] <= 8'h10 ;
			data[94258] <= 8'h10 ;
			data[94259] <= 8'h10 ;
			data[94260] <= 8'h10 ;
			data[94261] <= 8'h10 ;
			data[94262] <= 8'h10 ;
			data[94263] <= 8'h10 ;
			data[94264] <= 8'h10 ;
			data[94265] <= 8'h10 ;
			data[94266] <= 8'h10 ;
			data[94267] <= 8'h10 ;
			data[94268] <= 8'h10 ;
			data[94269] <= 8'h10 ;
			data[94270] <= 8'h10 ;
			data[94271] <= 8'h10 ;
			data[94272] <= 8'h10 ;
			data[94273] <= 8'h10 ;
			data[94274] <= 8'h10 ;
			data[94275] <= 8'h10 ;
			data[94276] <= 8'h10 ;
			data[94277] <= 8'h10 ;
			data[94278] <= 8'h10 ;
			data[94279] <= 8'h10 ;
			data[94280] <= 8'h10 ;
			data[94281] <= 8'h10 ;
			data[94282] <= 8'h10 ;
			data[94283] <= 8'h10 ;
			data[94284] <= 8'h10 ;
			data[94285] <= 8'h10 ;
			data[94286] <= 8'h10 ;
			data[94287] <= 8'h10 ;
			data[94288] <= 8'h10 ;
			data[94289] <= 8'h10 ;
			data[94290] <= 8'h10 ;
			data[94291] <= 8'h10 ;
			data[94292] <= 8'h10 ;
			data[94293] <= 8'h10 ;
			data[94294] <= 8'h10 ;
			data[94295] <= 8'h10 ;
			data[94296] <= 8'h10 ;
			data[94297] <= 8'h10 ;
			data[94298] <= 8'h10 ;
			data[94299] <= 8'h10 ;
			data[94300] <= 8'h10 ;
			data[94301] <= 8'h10 ;
			data[94302] <= 8'h10 ;
			data[94303] <= 8'h10 ;
			data[94304] <= 8'h10 ;
			data[94305] <= 8'h10 ;
			data[94306] <= 8'h10 ;
			data[94307] <= 8'h10 ;
			data[94308] <= 8'h10 ;
			data[94309] <= 8'h10 ;
			data[94310] <= 8'h10 ;
			data[94311] <= 8'h10 ;
			data[94312] <= 8'h10 ;
			data[94313] <= 8'h10 ;
			data[94314] <= 8'h10 ;
			data[94315] <= 8'h10 ;
			data[94316] <= 8'h10 ;
			data[94317] <= 8'h10 ;
			data[94318] <= 8'h10 ;
			data[94319] <= 8'h10 ;
			data[94320] <= 8'h10 ;
			data[94321] <= 8'h10 ;
			data[94322] <= 8'h10 ;
			data[94323] <= 8'h10 ;
			data[94324] <= 8'h10 ;
			data[94325] <= 8'h10 ;
			data[94326] <= 8'h10 ;
			data[94327] <= 8'h10 ;
			data[94328] <= 8'h10 ;
			data[94329] <= 8'h10 ;
			data[94330] <= 8'h10 ;
			data[94331] <= 8'h10 ;
			data[94332] <= 8'h10 ;
			data[94333] <= 8'h10 ;
			data[94334] <= 8'h10 ;
			data[94335] <= 8'h10 ;
			data[94336] <= 8'h10 ;
			data[94337] <= 8'h10 ;
			data[94338] <= 8'h10 ;
			data[94339] <= 8'h10 ;
			data[94340] <= 8'h10 ;
			data[94341] <= 8'h10 ;
			data[94342] <= 8'h10 ;
			data[94343] <= 8'h10 ;
			data[94344] <= 8'h10 ;
			data[94345] <= 8'h10 ;
			data[94346] <= 8'h10 ;
			data[94347] <= 8'h10 ;
			data[94348] <= 8'h10 ;
			data[94349] <= 8'h10 ;
			data[94350] <= 8'h10 ;
			data[94351] <= 8'h10 ;
			data[94352] <= 8'h10 ;
			data[94353] <= 8'h10 ;
			data[94354] <= 8'h10 ;
			data[94355] <= 8'h10 ;
			data[94356] <= 8'h10 ;
			data[94357] <= 8'h10 ;
			data[94358] <= 8'h10 ;
			data[94359] <= 8'h10 ;
			data[94360] <= 8'h10 ;
			data[94361] <= 8'h10 ;
			data[94362] <= 8'h10 ;
			data[94363] <= 8'h10 ;
			data[94364] <= 8'h10 ;
			data[94365] <= 8'h10 ;
			data[94366] <= 8'h10 ;
			data[94367] <= 8'h10 ;
			data[94368] <= 8'h10 ;
			data[94369] <= 8'h10 ;
			data[94370] <= 8'h10 ;
			data[94371] <= 8'h10 ;
			data[94372] <= 8'h10 ;
			data[94373] <= 8'h10 ;
			data[94374] <= 8'h10 ;
			data[94375] <= 8'h10 ;
			data[94376] <= 8'h10 ;
			data[94377] <= 8'h10 ;
			data[94378] <= 8'h10 ;
			data[94379] <= 8'h10 ;
			data[94380] <= 8'h10 ;
			data[94381] <= 8'h10 ;
			data[94382] <= 8'h10 ;
			data[94383] <= 8'h10 ;
			data[94384] <= 8'h10 ;
			data[94385] <= 8'h10 ;
			data[94386] <= 8'h10 ;
			data[94387] <= 8'h10 ;
			data[94388] <= 8'h10 ;
			data[94389] <= 8'h10 ;
			data[94390] <= 8'h10 ;
			data[94391] <= 8'h10 ;
			data[94392] <= 8'h10 ;
			data[94393] <= 8'h10 ;
			data[94394] <= 8'h10 ;
			data[94395] <= 8'h10 ;
			data[94396] <= 8'h10 ;
			data[94397] <= 8'h10 ;
			data[94398] <= 8'h10 ;
			data[94399] <= 8'h10 ;
			data[94400] <= 8'h10 ;
			data[94401] <= 8'h10 ;
			data[94402] <= 8'h10 ;
			data[94403] <= 8'h10 ;
			data[94404] <= 8'h10 ;
			data[94405] <= 8'h10 ;
			data[94406] <= 8'h10 ;
			data[94407] <= 8'h10 ;
			data[94408] <= 8'h10 ;
			data[94409] <= 8'h10 ;
			data[94410] <= 8'h10 ;
			data[94411] <= 8'h10 ;
			data[94412] <= 8'h10 ;
			data[94413] <= 8'h10 ;
			data[94414] <= 8'h10 ;
			data[94415] <= 8'h10 ;
			data[94416] <= 8'h10 ;
			data[94417] <= 8'h10 ;
			data[94418] <= 8'h10 ;
			data[94419] <= 8'h10 ;
			data[94420] <= 8'h10 ;
			data[94421] <= 8'h10 ;
			data[94422] <= 8'h10 ;
			data[94423] <= 8'h10 ;
			data[94424] <= 8'h10 ;
			data[94425] <= 8'h10 ;
			data[94426] <= 8'h10 ;
			data[94427] <= 8'h10 ;
			data[94428] <= 8'h10 ;
			data[94429] <= 8'h10 ;
			data[94430] <= 8'h10 ;
			data[94431] <= 8'h10 ;
			data[94432] <= 8'h10 ;
			data[94433] <= 8'h10 ;
			data[94434] <= 8'h10 ;
			data[94435] <= 8'h10 ;
			data[94436] <= 8'h10 ;
			data[94437] <= 8'h10 ;
			data[94438] <= 8'h10 ;
			data[94439] <= 8'h10 ;
			data[94440] <= 8'h10 ;
			data[94441] <= 8'h10 ;
			data[94442] <= 8'h10 ;
			data[94443] <= 8'h10 ;
			data[94444] <= 8'h10 ;
			data[94445] <= 8'h10 ;
			data[94446] <= 8'h10 ;
			data[94447] <= 8'h10 ;
			data[94448] <= 8'h10 ;
			data[94449] <= 8'h10 ;
			data[94450] <= 8'h10 ;
			data[94451] <= 8'h10 ;
			data[94452] <= 8'h10 ;
			data[94453] <= 8'h10 ;
			data[94454] <= 8'h10 ;
			data[94455] <= 8'h10 ;
			data[94456] <= 8'h10 ;
			data[94457] <= 8'h10 ;
			data[94458] <= 8'h10 ;
			data[94459] <= 8'h10 ;
			data[94460] <= 8'h10 ;
			data[94461] <= 8'h10 ;
			data[94462] <= 8'h10 ;
			data[94463] <= 8'h10 ;
			data[94464] <= 8'h10 ;
			data[94465] <= 8'h10 ;
			data[94466] <= 8'h10 ;
			data[94467] <= 8'h10 ;
			data[94468] <= 8'h10 ;
			data[94469] <= 8'h10 ;
			data[94470] <= 8'h10 ;
			data[94471] <= 8'h10 ;
			data[94472] <= 8'h10 ;
			data[94473] <= 8'h10 ;
			data[94474] <= 8'h10 ;
			data[94475] <= 8'h10 ;
			data[94476] <= 8'h10 ;
			data[94477] <= 8'h10 ;
			data[94478] <= 8'h10 ;
			data[94479] <= 8'h10 ;
			data[94480] <= 8'h10 ;
			data[94481] <= 8'h10 ;
			data[94482] <= 8'h10 ;
			data[94483] <= 8'h10 ;
			data[94484] <= 8'h10 ;
			data[94485] <= 8'h10 ;
			data[94486] <= 8'h10 ;
			data[94487] <= 8'h10 ;
			data[94488] <= 8'h10 ;
			data[94489] <= 8'h10 ;
			data[94490] <= 8'h10 ;
			data[94491] <= 8'h10 ;
			data[94492] <= 8'h10 ;
			data[94493] <= 8'h10 ;
			data[94494] <= 8'h10 ;
			data[94495] <= 8'h10 ;
			data[94496] <= 8'h10 ;
			data[94497] <= 8'h10 ;
			data[94498] <= 8'h10 ;
			data[94499] <= 8'h10 ;
			data[94500] <= 8'h10 ;
			data[94501] <= 8'h10 ;
			data[94502] <= 8'h10 ;
			data[94503] <= 8'h10 ;
			data[94504] <= 8'h10 ;
			data[94505] <= 8'h10 ;
			data[94506] <= 8'h10 ;
			data[94507] <= 8'h10 ;
			data[94508] <= 8'h10 ;
			data[94509] <= 8'h10 ;
			data[94510] <= 8'h10 ;
			data[94511] <= 8'h10 ;
			data[94512] <= 8'h10 ;
			data[94513] <= 8'h10 ;
			data[94514] <= 8'h10 ;
			data[94515] <= 8'h10 ;
			data[94516] <= 8'h10 ;
			data[94517] <= 8'h10 ;
			data[94518] <= 8'h10 ;
			data[94519] <= 8'h10 ;
			data[94520] <= 8'h10 ;
			data[94521] <= 8'h10 ;
			data[94522] <= 8'h10 ;
			data[94523] <= 8'h10 ;
			data[94524] <= 8'h10 ;
			data[94525] <= 8'h10 ;
			data[94526] <= 8'h10 ;
			data[94527] <= 8'h10 ;
			data[94528] <= 8'h10 ;
			data[94529] <= 8'h10 ;
			data[94530] <= 8'h10 ;
			data[94531] <= 8'h10 ;
			data[94532] <= 8'h10 ;
			data[94533] <= 8'h10 ;
			data[94534] <= 8'h10 ;
			data[94535] <= 8'h10 ;
			data[94536] <= 8'h10 ;
			data[94537] <= 8'h10 ;
			data[94538] <= 8'h10 ;
			data[94539] <= 8'h10 ;
			data[94540] <= 8'h10 ;
			data[94541] <= 8'h10 ;
			data[94542] <= 8'h10 ;
			data[94543] <= 8'h10 ;
			data[94544] <= 8'h10 ;
			data[94545] <= 8'h10 ;
			data[94546] <= 8'h10 ;
			data[94547] <= 8'h10 ;
			data[94548] <= 8'h10 ;
			data[94549] <= 8'h10 ;
			data[94550] <= 8'h10 ;
			data[94551] <= 8'h10 ;
			data[94552] <= 8'h10 ;
			data[94553] <= 8'h10 ;
			data[94554] <= 8'h10 ;
			data[94555] <= 8'h10 ;
			data[94556] <= 8'h10 ;
			data[94557] <= 8'h10 ;
			data[94558] <= 8'h10 ;
			data[94559] <= 8'h10 ;
			data[94560] <= 8'h10 ;
			data[94561] <= 8'h10 ;
			data[94562] <= 8'h10 ;
			data[94563] <= 8'h10 ;
			data[94564] <= 8'h10 ;
			data[94565] <= 8'h10 ;
			data[94566] <= 8'h10 ;
			data[94567] <= 8'h10 ;
			data[94568] <= 8'h10 ;
			data[94569] <= 8'h10 ;
			data[94570] <= 8'h10 ;
			data[94571] <= 8'h10 ;
			data[94572] <= 8'h10 ;
			data[94573] <= 8'h10 ;
			data[94574] <= 8'h10 ;
			data[94575] <= 8'h10 ;
			data[94576] <= 8'h10 ;
			data[94577] <= 8'h10 ;
			data[94578] <= 8'h10 ;
			data[94579] <= 8'h10 ;
			data[94580] <= 8'h10 ;
			data[94581] <= 8'h10 ;
			data[94582] <= 8'h10 ;
			data[94583] <= 8'h10 ;
			data[94584] <= 8'h10 ;
			data[94585] <= 8'h10 ;
			data[94586] <= 8'h10 ;
			data[94587] <= 8'h10 ;
			data[94588] <= 8'h10 ;
			data[94589] <= 8'h10 ;
			data[94590] <= 8'h10 ;
			data[94591] <= 8'h10 ;
			data[94592] <= 8'h10 ;
			data[94593] <= 8'h10 ;
			data[94594] <= 8'h10 ;
			data[94595] <= 8'h10 ;
			data[94596] <= 8'h10 ;
			data[94597] <= 8'h10 ;
			data[94598] <= 8'h10 ;
			data[94599] <= 8'h10 ;
			data[94600] <= 8'h10 ;
			data[94601] <= 8'h10 ;
			data[94602] <= 8'h10 ;
			data[94603] <= 8'h10 ;
			data[94604] <= 8'h10 ;
			data[94605] <= 8'h10 ;
			data[94606] <= 8'h10 ;
			data[94607] <= 8'h10 ;
			data[94608] <= 8'h10 ;
			data[94609] <= 8'h10 ;
			data[94610] <= 8'h10 ;
			data[94611] <= 8'h10 ;
			data[94612] <= 8'h10 ;
			data[94613] <= 8'h10 ;
			data[94614] <= 8'h10 ;
			data[94615] <= 8'h10 ;
			data[94616] <= 8'h10 ;
			data[94617] <= 8'h10 ;
			data[94618] <= 8'h10 ;
			data[94619] <= 8'h10 ;
			data[94620] <= 8'h10 ;
			data[94621] <= 8'h10 ;
			data[94622] <= 8'h10 ;
			data[94623] <= 8'h10 ;
			data[94624] <= 8'h10 ;
			data[94625] <= 8'h10 ;
			data[94626] <= 8'h10 ;
			data[94627] <= 8'h10 ;
			data[94628] <= 8'h10 ;
			data[94629] <= 8'h10 ;
			data[94630] <= 8'h10 ;
			data[94631] <= 8'h10 ;
			data[94632] <= 8'h10 ;
			data[94633] <= 8'h10 ;
			data[94634] <= 8'h10 ;
			data[94635] <= 8'h10 ;
			data[94636] <= 8'h10 ;
			data[94637] <= 8'h10 ;
			data[94638] <= 8'h10 ;
			data[94639] <= 8'h10 ;
			data[94640] <= 8'h10 ;
			data[94641] <= 8'h10 ;
			data[94642] <= 8'h10 ;
			data[94643] <= 8'h10 ;
			data[94644] <= 8'h10 ;
			data[94645] <= 8'h10 ;
			data[94646] <= 8'h10 ;
			data[94647] <= 8'h10 ;
			data[94648] <= 8'h10 ;
			data[94649] <= 8'h10 ;
			data[94650] <= 8'h10 ;
			data[94651] <= 8'h10 ;
			data[94652] <= 8'h10 ;
			data[94653] <= 8'h10 ;
			data[94654] <= 8'h10 ;
			data[94655] <= 8'h10 ;
			data[94656] <= 8'h10 ;
			data[94657] <= 8'h10 ;
			data[94658] <= 8'h10 ;
			data[94659] <= 8'h10 ;
			data[94660] <= 8'h10 ;
			data[94661] <= 8'h10 ;
			data[94662] <= 8'h10 ;
			data[94663] <= 8'h10 ;
			data[94664] <= 8'h10 ;
			data[94665] <= 8'h10 ;
			data[94666] <= 8'h10 ;
			data[94667] <= 8'h10 ;
			data[94668] <= 8'h10 ;
			data[94669] <= 8'h10 ;
			data[94670] <= 8'h10 ;
			data[94671] <= 8'h10 ;
			data[94672] <= 8'h10 ;
			data[94673] <= 8'h10 ;
			data[94674] <= 8'h10 ;
			data[94675] <= 8'h10 ;
			data[94676] <= 8'h10 ;
			data[94677] <= 8'h10 ;
			data[94678] <= 8'h10 ;
			data[94679] <= 8'h10 ;
			data[94680] <= 8'h10 ;
			data[94681] <= 8'h10 ;
			data[94682] <= 8'h10 ;
			data[94683] <= 8'h10 ;
			data[94684] <= 8'h10 ;
			data[94685] <= 8'h10 ;
			data[94686] <= 8'h10 ;
			data[94687] <= 8'h10 ;
			data[94688] <= 8'h10 ;
			data[94689] <= 8'h10 ;
			data[94690] <= 8'h10 ;
			data[94691] <= 8'h10 ;
			data[94692] <= 8'h10 ;
			data[94693] <= 8'h10 ;
			data[94694] <= 8'h10 ;
			data[94695] <= 8'h10 ;
			data[94696] <= 8'h10 ;
			data[94697] <= 8'h10 ;
			data[94698] <= 8'h10 ;
			data[94699] <= 8'h10 ;
			data[94700] <= 8'h10 ;
			data[94701] <= 8'h10 ;
			data[94702] <= 8'h10 ;
			data[94703] <= 8'h10 ;
			data[94704] <= 8'h10 ;
			data[94705] <= 8'h10 ;
			data[94706] <= 8'h10 ;
			data[94707] <= 8'h10 ;
			data[94708] <= 8'h10 ;
			data[94709] <= 8'h10 ;
			data[94710] <= 8'h10 ;
			data[94711] <= 8'h10 ;
			data[94712] <= 8'h10 ;
			data[94713] <= 8'h10 ;
			data[94714] <= 8'h10 ;
			data[94715] <= 8'h10 ;
			data[94716] <= 8'h10 ;
			data[94717] <= 8'h10 ;
			data[94718] <= 8'h10 ;
			data[94719] <= 8'h10 ;
			data[94720] <= 8'h10 ;
			data[94721] <= 8'h10 ;
			data[94722] <= 8'h10 ;
			data[94723] <= 8'h10 ;
			data[94724] <= 8'h10 ;
			data[94725] <= 8'h10 ;
			data[94726] <= 8'h10 ;
			data[94727] <= 8'h10 ;
			data[94728] <= 8'h10 ;
			data[94729] <= 8'h10 ;
			data[94730] <= 8'h10 ;
			data[94731] <= 8'h10 ;
			data[94732] <= 8'h10 ;
			data[94733] <= 8'h10 ;
			data[94734] <= 8'h10 ;
			data[94735] <= 8'h10 ;
			data[94736] <= 8'h10 ;
			data[94737] <= 8'h10 ;
			data[94738] <= 8'h10 ;
			data[94739] <= 8'h10 ;
			data[94740] <= 8'h10 ;
			data[94741] <= 8'h10 ;
			data[94742] <= 8'h10 ;
			data[94743] <= 8'h10 ;
			data[94744] <= 8'h10 ;
			data[94745] <= 8'h10 ;
			data[94746] <= 8'h10 ;
			data[94747] <= 8'h10 ;
			data[94748] <= 8'h10 ;
			data[94749] <= 8'h10 ;
			data[94750] <= 8'h10 ;
			data[94751] <= 8'h10 ;
			data[94752] <= 8'h10 ;
			data[94753] <= 8'h10 ;
			data[94754] <= 8'h10 ;
			data[94755] <= 8'h10 ;
			data[94756] <= 8'h10 ;
			data[94757] <= 8'h10 ;
			data[94758] <= 8'h10 ;
			data[94759] <= 8'h10 ;
			data[94760] <= 8'h10 ;
			data[94761] <= 8'h10 ;
			data[94762] <= 8'h10 ;
			data[94763] <= 8'h10 ;
			data[94764] <= 8'h10 ;
			data[94765] <= 8'h10 ;
			data[94766] <= 8'h10 ;
			data[94767] <= 8'h10 ;
			data[94768] <= 8'h10 ;
			data[94769] <= 8'h10 ;
			data[94770] <= 8'h10 ;
			data[94771] <= 8'h10 ;
			data[94772] <= 8'h10 ;
			data[94773] <= 8'h10 ;
			data[94774] <= 8'h10 ;
			data[94775] <= 8'h10 ;
			data[94776] <= 8'h10 ;
			data[94777] <= 8'h10 ;
			data[94778] <= 8'h10 ;
			data[94779] <= 8'h10 ;
			data[94780] <= 8'h10 ;
			data[94781] <= 8'h10 ;
			data[94782] <= 8'h10 ;
			data[94783] <= 8'h10 ;
			data[94784] <= 8'h10 ;
			data[94785] <= 8'h10 ;
			data[94786] <= 8'h10 ;
			data[94787] <= 8'h10 ;
			data[94788] <= 8'h10 ;
			data[94789] <= 8'h10 ;
			data[94790] <= 8'h10 ;
			data[94791] <= 8'h10 ;
			data[94792] <= 8'h10 ;
			data[94793] <= 8'h10 ;
			data[94794] <= 8'h10 ;
			data[94795] <= 8'h10 ;
			data[94796] <= 8'h10 ;
			data[94797] <= 8'h10 ;
			data[94798] <= 8'h10 ;
			data[94799] <= 8'h10 ;
			data[94800] <= 8'h10 ;
			data[94801] <= 8'h10 ;
			data[94802] <= 8'h10 ;
			data[94803] <= 8'h10 ;
			data[94804] <= 8'h10 ;
			data[94805] <= 8'h10 ;
			data[94806] <= 8'h10 ;
			data[94807] <= 8'h10 ;
			data[94808] <= 8'h10 ;
			data[94809] <= 8'h10 ;
			data[94810] <= 8'h10 ;
			data[94811] <= 8'h10 ;
			data[94812] <= 8'h10 ;
			data[94813] <= 8'h10 ;
			data[94814] <= 8'h10 ;
			data[94815] <= 8'h10 ;
			data[94816] <= 8'h10 ;
			data[94817] <= 8'h10 ;
			data[94818] <= 8'h10 ;
			data[94819] <= 8'h10 ;
			data[94820] <= 8'h10 ;
			data[94821] <= 8'h10 ;
			data[94822] <= 8'h10 ;
			data[94823] <= 8'h10 ;
			data[94824] <= 8'h10 ;
			data[94825] <= 8'h10 ;
			data[94826] <= 8'h10 ;
			data[94827] <= 8'h10 ;
			data[94828] <= 8'h10 ;
			data[94829] <= 8'h10 ;
			data[94830] <= 8'h10 ;
			data[94831] <= 8'h10 ;
			data[94832] <= 8'h10 ;
			data[94833] <= 8'h10 ;
			data[94834] <= 8'h10 ;
			data[94835] <= 8'h10 ;
			data[94836] <= 8'h10 ;
			data[94837] <= 8'h10 ;
			data[94838] <= 8'h10 ;
			data[94839] <= 8'h10 ;
			data[94840] <= 8'h10 ;
			data[94841] <= 8'h10 ;
			data[94842] <= 8'h10 ;
			data[94843] <= 8'h10 ;
			data[94844] <= 8'h10 ;
			data[94845] <= 8'h10 ;
			data[94846] <= 8'h10 ;
			data[94847] <= 8'h10 ;
			data[94848] <= 8'h10 ;
			data[94849] <= 8'h10 ;
			data[94850] <= 8'h10 ;
			data[94851] <= 8'h10 ;
			data[94852] <= 8'h10 ;
			data[94853] <= 8'h10 ;
			data[94854] <= 8'h10 ;
			data[94855] <= 8'h10 ;
			data[94856] <= 8'h10 ;
			data[94857] <= 8'h10 ;
			data[94858] <= 8'h10 ;
			data[94859] <= 8'h10 ;
			data[94860] <= 8'h10 ;
			data[94861] <= 8'h10 ;
			data[94862] <= 8'h10 ;
			data[94863] <= 8'h10 ;
			data[94864] <= 8'h10 ;
			data[94865] <= 8'h10 ;
			data[94866] <= 8'h10 ;
			data[94867] <= 8'h10 ;
			data[94868] <= 8'h10 ;
			data[94869] <= 8'h10 ;
			data[94870] <= 8'h10 ;
			data[94871] <= 8'h10 ;
			data[94872] <= 8'h10 ;
			data[94873] <= 8'h10 ;
			data[94874] <= 8'h10 ;
			data[94875] <= 8'h10 ;
			data[94876] <= 8'h10 ;
			data[94877] <= 8'h10 ;
			data[94878] <= 8'h10 ;
			data[94879] <= 8'h10 ;
			data[94880] <= 8'h10 ;
			data[94881] <= 8'h10 ;
			data[94882] <= 8'h10 ;
			data[94883] <= 8'h10 ;
			data[94884] <= 8'h10 ;
			data[94885] <= 8'h10 ;
			data[94886] <= 8'h10 ;
			data[94887] <= 8'h10 ;
			data[94888] <= 8'h10 ;
			data[94889] <= 8'h10 ;
			data[94890] <= 8'h10 ;
			data[94891] <= 8'h10 ;
			data[94892] <= 8'h10 ;
			data[94893] <= 8'h10 ;
			data[94894] <= 8'h10 ;
			data[94895] <= 8'h10 ;
			data[94896] <= 8'h10 ;
			data[94897] <= 8'h10 ;
			data[94898] <= 8'h10 ;
			data[94899] <= 8'h10 ;
			data[94900] <= 8'h10 ;
			data[94901] <= 8'h10 ;
			data[94902] <= 8'h10 ;
			data[94903] <= 8'h10 ;
			data[94904] <= 8'h10 ;
			data[94905] <= 8'h10 ;
			data[94906] <= 8'h10 ;
			data[94907] <= 8'h10 ;
			data[94908] <= 8'h10 ;
			data[94909] <= 8'h10 ;
			data[94910] <= 8'h10 ;
			data[94911] <= 8'h10 ;
			data[94912] <= 8'h10 ;
			data[94913] <= 8'h10 ;
			data[94914] <= 8'h10 ;
			data[94915] <= 8'h10 ;
			data[94916] <= 8'h10 ;
			data[94917] <= 8'h10 ;
			data[94918] <= 8'h10 ;
			data[94919] <= 8'h10 ;
			data[94920] <= 8'h10 ;
			data[94921] <= 8'h10 ;
			data[94922] <= 8'h10 ;
			data[94923] <= 8'h10 ;
			data[94924] <= 8'h10 ;
			data[94925] <= 8'h10 ;
			data[94926] <= 8'h10 ;
			data[94927] <= 8'h10 ;
			data[94928] <= 8'h10 ;
			data[94929] <= 8'h10 ;
			data[94930] <= 8'h10 ;
			data[94931] <= 8'h10 ;
			data[94932] <= 8'h10 ;
			data[94933] <= 8'h10 ;
			data[94934] <= 8'h10 ;
			data[94935] <= 8'h10 ;
			data[94936] <= 8'h10 ;
			data[94937] <= 8'h10 ;
			data[94938] <= 8'h10 ;
			data[94939] <= 8'h10 ;
			data[94940] <= 8'h10 ;
			data[94941] <= 8'h10 ;
			data[94942] <= 8'h10 ;
			data[94943] <= 8'h10 ;
			data[94944] <= 8'h10 ;
			data[94945] <= 8'h10 ;
			data[94946] <= 8'h10 ;
			data[94947] <= 8'h10 ;
			data[94948] <= 8'h10 ;
			data[94949] <= 8'h10 ;
			data[94950] <= 8'h10 ;
			data[94951] <= 8'h10 ;
			data[94952] <= 8'h10 ;
			data[94953] <= 8'h10 ;
			data[94954] <= 8'h10 ;
			data[94955] <= 8'h10 ;
			data[94956] <= 8'h10 ;
			data[94957] <= 8'h10 ;
			data[94958] <= 8'h10 ;
			data[94959] <= 8'h10 ;
			data[94960] <= 8'h10 ;
			data[94961] <= 8'h10 ;
			data[94962] <= 8'h10 ;
			data[94963] <= 8'h10 ;
			data[94964] <= 8'h10 ;
			data[94965] <= 8'h10 ;
			data[94966] <= 8'h10 ;
			data[94967] <= 8'h10 ;
			data[94968] <= 8'h10 ;
			data[94969] <= 8'h10 ;
			data[94970] <= 8'h10 ;
			data[94971] <= 8'h10 ;
			data[94972] <= 8'h10 ;
			data[94973] <= 8'h10 ;
			data[94974] <= 8'h10 ;
			data[94975] <= 8'h10 ;
			data[94976] <= 8'h10 ;
			data[94977] <= 8'h10 ;
			data[94978] <= 8'h10 ;
			data[94979] <= 8'h10 ;
			data[94980] <= 8'h10 ;
			data[94981] <= 8'h10 ;
			data[94982] <= 8'h10 ;
			data[94983] <= 8'h10 ;
			data[94984] <= 8'h10 ;
			data[94985] <= 8'h10 ;
			data[94986] <= 8'h10 ;
			data[94987] <= 8'h10 ;
			data[94988] <= 8'h10 ;
			data[94989] <= 8'h10 ;
			data[94990] <= 8'h10 ;
			data[94991] <= 8'h10 ;
			data[94992] <= 8'h10 ;
			data[94993] <= 8'h10 ;
			data[94994] <= 8'h10 ;
			data[94995] <= 8'h10 ;
			data[94996] <= 8'h10 ;
			data[94997] <= 8'h10 ;
			data[94998] <= 8'h10 ;
			data[94999] <= 8'h10 ;
			data[95000] <= 8'h10 ;
			data[95001] <= 8'h10 ;
			data[95002] <= 8'h10 ;
			data[95003] <= 8'h10 ;
			data[95004] <= 8'h10 ;
			data[95005] <= 8'h10 ;
			data[95006] <= 8'h10 ;
			data[95007] <= 8'h10 ;
			data[95008] <= 8'h10 ;
			data[95009] <= 8'h10 ;
			data[95010] <= 8'h10 ;
			data[95011] <= 8'h10 ;
			data[95012] <= 8'h10 ;
			data[95013] <= 8'h10 ;
			data[95014] <= 8'h10 ;
			data[95015] <= 8'h10 ;
			data[95016] <= 8'h10 ;
			data[95017] <= 8'h10 ;
			data[95018] <= 8'h10 ;
			data[95019] <= 8'h10 ;
			data[95020] <= 8'h10 ;
			data[95021] <= 8'h10 ;
			data[95022] <= 8'h10 ;
			data[95023] <= 8'h10 ;
			data[95024] <= 8'h10 ;
			data[95025] <= 8'h10 ;
			data[95026] <= 8'h10 ;
			data[95027] <= 8'h10 ;
			data[95028] <= 8'h10 ;
			data[95029] <= 8'h10 ;
			data[95030] <= 8'h10 ;
			data[95031] <= 8'h10 ;
			data[95032] <= 8'h10 ;
			data[95033] <= 8'h10 ;
			data[95034] <= 8'h10 ;
			data[95035] <= 8'h10 ;
			data[95036] <= 8'h10 ;
			data[95037] <= 8'h10 ;
			data[95038] <= 8'h10 ;
			data[95039] <= 8'h10 ;
			data[95040] <= 8'h10 ;
			data[95041] <= 8'h10 ;
			data[95042] <= 8'h10 ;
			data[95043] <= 8'h10 ;
			data[95044] <= 8'h10 ;
			data[95045] <= 8'h10 ;
			data[95046] <= 8'h10 ;
			data[95047] <= 8'h10 ;
			data[95048] <= 8'h10 ;
			data[95049] <= 8'h10 ;
			data[95050] <= 8'h10 ;
			data[95051] <= 8'h10 ;
			data[95052] <= 8'h10 ;
			data[95053] <= 8'h10 ;
			data[95054] <= 8'h10 ;
			data[95055] <= 8'h10 ;
			data[95056] <= 8'h10 ;
			data[95057] <= 8'h10 ;
			data[95058] <= 8'h10 ;
			data[95059] <= 8'h10 ;
			data[95060] <= 8'h10 ;
			data[95061] <= 8'h10 ;
			data[95062] <= 8'h10 ;
			data[95063] <= 8'h10 ;
			data[95064] <= 8'h10 ;
			data[95065] <= 8'h10 ;
			data[95066] <= 8'h10 ;
			data[95067] <= 8'h10 ;
			data[95068] <= 8'h10 ;
			data[95069] <= 8'h10 ;
			data[95070] <= 8'h10 ;
			data[95071] <= 8'h10 ;
			data[95072] <= 8'h10 ;
			data[95073] <= 8'h10 ;
			data[95074] <= 8'h10 ;
			data[95075] <= 8'h10 ;
			data[95076] <= 8'h10 ;
			data[95077] <= 8'h10 ;
			data[95078] <= 8'h10 ;
			data[95079] <= 8'h10 ;
			data[95080] <= 8'h10 ;
			data[95081] <= 8'h10 ;
			data[95082] <= 8'h10 ;
			data[95083] <= 8'h10 ;
			data[95084] <= 8'h10 ;
			data[95085] <= 8'h10 ;
			data[95086] <= 8'h10 ;
			data[95087] <= 8'h10 ;
			data[95088] <= 8'h10 ;
			data[95089] <= 8'h10 ;
			data[95090] <= 8'h10 ;
			data[95091] <= 8'h10 ;
			data[95092] <= 8'h10 ;
			data[95093] <= 8'h10 ;
			data[95094] <= 8'h10 ;
			data[95095] <= 8'h10 ;
			data[95096] <= 8'h10 ;
			data[95097] <= 8'h10 ;
			data[95098] <= 8'h10 ;
			data[95099] <= 8'h10 ;
			data[95100] <= 8'h10 ;
			data[95101] <= 8'h10 ;
			data[95102] <= 8'h10 ;
			data[95103] <= 8'h10 ;
			data[95104] <= 8'h10 ;
			data[95105] <= 8'h10 ;
			data[95106] <= 8'h10 ;
			data[95107] <= 8'h10 ;
			data[95108] <= 8'h10 ;
			data[95109] <= 8'h10 ;
			data[95110] <= 8'h10 ;
			data[95111] <= 8'h10 ;
			data[95112] <= 8'h10 ;
			data[95113] <= 8'h10 ;
			data[95114] <= 8'h10 ;
			data[95115] <= 8'h10 ;
			data[95116] <= 8'h10 ;
			data[95117] <= 8'h10 ;
			data[95118] <= 8'h10 ;
			data[95119] <= 8'h10 ;
			data[95120] <= 8'h10 ;
			data[95121] <= 8'h10 ;
			data[95122] <= 8'h10 ;
			data[95123] <= 8'h10 ;
			data[95124] <= 8'h10 ;
			data[95125] <= 8'h10 ;
			data[95126] <= 8'h10 ;
			data[95127] <= 8'h10 ;
			data[95128] <= 8'h10 ;
			data[95129] <= 8'h10 ;
			data[95130] <= 8'h10 ;
			data[95131] <= 8'h10 ;
			data[95132] <= 8'h10 ;
			data[95133] <= 8'h10 ;
			data[95134] <= 8'h10 ;
			data[95135] <= 8'h10 ;
			data[95136] <= 8'h10 ;
			data[95137] <= 8'h10 ;
			data[95138] <= 8'h10 ;
			data[95139] <= 8'h10 ;
			data[95140] <= 8'h10 ;
			data[95141] <= 8'h10 ;
			data[95142] <= 8'h10 ;
			data[95143] <= 8'h10 ;
			data[95144] <= 8'h10 ;
			data[95145] <= 8'h10 ;
			data[95146] <= 8'h10 ;
			data[95147] <= 8'h10 ;
			data[95148] <= 8'h10 ;
			data[95149] <= 8'h10 ;
			data[95150] <= 8'h10 ;
			data[95151] <= 8'h10 ;
			data[95152] <= 8'h10 ;
			data[95153] <= 8'h10 ;
			data[95154] <= 8'h10 ;
			data[95155] <= 8'h10 ;
			data[95156] <= 8'h10 ;
			data[95157] <= 8'h10 ;
			data[95158] <= 8'h10 ;
			data[95159] <= 8'h10 ;
			data[95160] <= 8'h10 ;
			data[95161] <= 8'h10 ;
			data[95162] <= 8'h10 ;
			data[95163] <= 8'h10 ;
			data[95164] <= 8'h10 ;
			data[95165] <= 8'h10 ;
			data[95166] <= 8'h10 ;
			data[95167] <= 8'h10 ;
			data[95168] <= 8'h10 ;
			data[95169] <= 8'h10 ;
			data[95170] <= 8'h10 ;
			data[95171] <= 8'h10 ;
			data[95172] <= 8'h10 ;
			data[95173] <= 8'h10 ;
			data[95174] <= 8'h10 ;
			data[95175] <= 8'h10 ;
			data[95176] <= 8'h10 ;
			data[95177] <= 8'h10 ;
			data[95178] <= 8'h10 ;
			data[95179] <= 8'h10 ;
			data[95180] <= 8'h10 ;
			data[95181] <= 8'h10 ;
			data[95182] <= 8'h10 ;
			data[95183] <= 8'h10 ;
			data[95184] <= 8'h10 ;
			data[95185] <= 8'h10 ;
			data[95186] <= 8'h10 ;
			data[95187] <= 8'h10 ;
			data[95188] <= 8'h10 ;
			data[95189] <= 8'h10 ;
			data[95190] <= 8'h10 ;
			data[95191] <= 8'h10 ;
			data[95192] <= 8'h10 ;
			data[95193] <= 8'h10 ;
			data[95194] <= 8'h10 ;
			data[95195] <= 8'h10 ;
			data[95196] <= 8'h10 ;
			data[95197] <= 8'h10 ;
			data[95198] <= 8'h10 ;
			data[95199] <= 8'h10 ;
			data[95200] <= 8'h10 ;
			data[95201] <= 8'h10 ;
			data[95202] <= 8'h10 ;
			data[95203] <= 8'h10 ;
			data[95204] <= 8'h10 ;
			data[95205] <= 8'h10 ;
			data[95206] <= 8'h10 ;
			data[95207] <= 8'h10 ;
			data[95208] <= 8'h10 ;
			data[95209] <= 8'h10 ;
			data[95210] <= 8'h10 ;
			data[95211] <= 8'h10 ;
			data[95212] <= 8'h10 ;
			data[95213] <= 8'h10 ;
			data[95214] <= 8'h10 ;
			data[95215] <= 8'h10 ;
			data[95216] <= 8'h10 ;
			data[95217] <= 8'h10 ;
			data[95218] <= 8'h10 ;
			data[95219] <= 8'h10 ;
			data[95220] <= 8'h10 ;
			data[95221] <= 8'h10 ;
			data[95222] <= 8'h10 ;
			data[95223] <= 8'h10 ;
			data[95224] <= 8'h10 ;
			data[95225] <= 8'h10 ;
			data[95226] <= 8'h10 ;
			data[95227] <= 8'h10 ;
			data[95228] <= 8'h10 ;
			data[95229] <= 8'h10 ;
			data[95230] <= 8'h10 ;
			data[95231] <= 8'h10 ;
			data[95232] <= 8'h10 ;
			data[95233] <= 8'h10 ;
			data[95234] <= 8'h10 ;
			data[95235] <= 8'h10 ;
			data[95236] <= 8'h10 ;
			data[95237] <= 8'h10 ;
			data[95238] <= 8'h10 ;
			data[95239] <= 8'h10 ;
			data[95240] <= 8'h10 ;
			data[95241] <= 8'h10 ;
			data[95242] <= 8'h10 ;
			data[95243] <= 8'h10 ;
			data[95244] <= 8'h10 ;
			data[95245] <= 8'h10 ;
			data[95246] <= 8'h10 ;
			data[95247] <= 8'h10 ;
			data[95248] <= 8'h10 ;
			data[95249] <= 8'h10 ;
			data[95250] <= 8'h10 ;
			data[95251] <= 8'h10 ;
			data[95252] <= 8'h10 ;
			data[95253] <= 8'h10 ;
			data[95254] <= 8'h10 ;
			data[95255] <= 8'h10 ;
			data[95256] <= 8'h10 ;
			data[95257] <= 8'h10 ;
			data[95258] <= 8'h10 ;
			data[95259] <= 8'h10 ;
			data[95260] <= 8'h10 ;
			data[95261] <= 8'h10 ;
			data[95262] <= 8'h10 ;
			data[95263] <= 8'h10 ;
			data[95264] <= 8'h10 ;
			data[95265] <= 8'h10 ;
			data[95266] <= 8'h10 ;
			data[95267] <= 8'h10 ;
			data[95268] <= 8'h10 ;
			data[95269] <= 8'h10 ;
			data[95270] <= 8'h10 ;
			data[95271] <= 8'h10 ;
			data[95272] <= 8'h10 ;
			data[95273] <= 8'h10 ;
			data[95274] <= 8'h10 ;
			data[95275] <= 8'h10 ;
			data[95276] <= 8'h10 ;
			data[95277] <= 8'h10 ;
			data[95278] <= 8'h10 ;
			data[95279] <= 8'h10 ;
			data[95280] <= 8'h10 ;
			data[95281] <= 8'h10 ;
			data[95282] <= 8'h10 ;
			data[95283] <= 8'h10 ;
			data[95284] <= 8'h10 ;
			data[95285] <= 8'h10 ;
			data[95286] <= 8'h10 ;
			data[95287] <= 8'h10 ;
			data[95288] <= 8'h10 ;
			data[95289] <= 8'h10 ;
			data[95290] <= 8'h10 ;
			data[95291] <= 8'h10 ;
			data[95292] <= 8'h10 ;
			data[95293] <= 8'h10 ;
			data[95294] <= 8'h10 ;
			data[95295] <= 8'h10 ;
			data[95296] <= 8'h10 ;
			data[95297] <= 8'h10 ;
			data[95298] <= 8'h10 ;
			data[95299] <= 8'h10 ;
			data[95300] <= 8'h10 ;
			data[95301] <= 8'h10 ;
			data[95302] <= 8'h10 ;
			data[95303] <= 8'h10 ;
			data[95304] <= 8'h10 ;
			data[95305] <= 8'h10 ;
			data[95306] <= 8'h10 ;
			data[95307] <= 8'h10 ;
			data[95308] <= 8'h10 ;
			data[95309] <= 8'h10 ;
			data[95310] <= 8'h10 ;
			data[95311] <= 8'h10 ;
			data[95312] <= 8'h10 ;
			data[95313] <= 8'h10 ;
			data[95314] <= 8'h10 ;
			data[95315] <= 8'h10 ;
			data[95316] <= 8'h10 ;
			data[95317] <= 8'h10 ;
			data[95318] <= 8'h10 ;
			data[95319] <= 8'h10 ;
			data[95320] <= 8'h10 ;
			data[95321] <= 8'h10 ;
			data[95322] <= 8'h10 ;
			data[95323] <= 8'h10 ;
			data[95324] <= 8'h10 ;
			data[95325] <= 8'h10 ;
			data[95326] <= 8'h10 ;
			data[95327] <= 8'h10 ;
			data[95328] <= 8'h10 ;
			data[95329] <= 8'h10 ;
			data[95330] <= 8'h10 ;
			data[95331] <= 8'h10 ;
			data[95332] <= 8'h10 ;
			data[95333] <= 8'h10 ;
			data[95334] <= 8'h10 ;
			data[95335] <= 8'h10 ;
			data[95336] <= 8'h10 ;
			data[95337] <= 8'h10 ;
			data[95338] <= 8'h10 ;
			data[95339] <= 8'h10 ;
			data[95340] <= 8'h10 ;
			data[95341] <= 8'h10 ;
			data[95342] <= 8'h10 ;
			data[95343] <= 8'h10 ;
			data[95344] <= 8'h10 ;
			data[95345] <= 8'h10 ;
			data[95346] <= 8'h10 ;
			data[95347] <= 8'h10 ;
			data[95348] <= 8'h10 ;
			data[95349] <= 8'h10 ;
			data[95350] <= 8'h10 ;
			data[95351] <= 8'h10 ;
			data[95352] <= 8'h10 ;
			data[95353] <= 8'h10 ;
			data[95354] <= 8'h10 ;
			data[95355] <= 8'h10 ;
			data[95356] <= 8'h10 ;
			data[95357] <= 8'h10 ;
			data[95358] <= 8'h10 ;
			data[95359] <= 8'h10 ;
			data[95360] <= 8'h10 ;
			data[95361] <= 8'h10 ;
			data[95362] <= 8'h10 ;
			data[95363] <= 8'h10 ;
			data[95364] <= 8'h10 ;
			data[95365] <= 8'h10 ;
			data[95366] <= 8'h10 ;
			data[95367] <= 8'h10 ;
			data[95368] <= 8'h10 ;
			data[95369] <= 8'h10 ;
			data[95370] <= 8'h10 ;
			data[95371] <= 8'h10 ;
			data[95372] <= 8'h10 ;
			data[95373] <= 8'h10 ;
			data[95374] <= 8'h10 ;
			data[95375] <= 8'h10 ;
			data[95376] <= 8'h10 ;
			data[95377] <= 8'h10 ;
			data[95378] <= 8'h10 ;
			data[95379] <= 8'h10 ;
			data[95380] <= 8'h10 ;
			data[95381] <= 8'h10 ;
			data[95382] <= 8'h10 ;
			data[95383] <= 8'h10 ;
			data[95384] <= 8'h10 ;
			data[95385] <= 8'h10 ;
			data[95386] <= 8'h10 ;
			data[95387] <= 8'h10 ;
			data[95388] <= 8'h10 ;
			data[95389] <= 8'h10 ;
			data[95390] <= 8'h10 ;
			data[95391] <= 8'h10 ;
			data[95392] <= 8'h10 ;
			data[95393] <= 8'h10 ;
			data[95394] <= 8'h10 ;
			data[95395] <= 8'h10 ;
			data[95396] <= 8'h10 ;
			data[95397] <= 8'h10 ;
			data[95398] <= 8'h10 ;
			data[95399] <= 8'h10 ;
			data[95400] <= 8'h10 ;
			data[95401] <= 8'h10 ;
			data[95402] <= 8'h10 ;
			data[95403] <= 8'h10 ;
			data[95404] <= 8'h10 ;
			data[95405] <= 8'h10 ;
			data[95406] <= 8'h10 ;
			data[95407] <= 8'h10 ;
			data[95408] <= 8'h10 ;
			data[95409] <= 8'h10 ;
			data[95410] <= 8'h10 ;
			data[95411] <= 8'h10 ;
			data[95412] <= 8'h10 ;
			data[95413] <= 8'h10 ;
			data[95414] <= 8'h10 ;
			data[95415] <= 8'h10 ;
			data[95416] <= 8'h10 ;
			data[95417] <= 8'h10 ;
			data[95418] <= 8'h10 ;
			data[95419] <= 8'h10 ;
			data[95420] <= 8'h10 ;
			data[95421] <= 8'h10 ;
			data[95422] <= 8'h10 ;
			data[95423] <= 8'h10 ;
			data[95424] <= 8'h10 ;
			data[95425] <= 8'h10 ;
			data[95426] <= 8'h10 ;
			data[95427] <= 8'h10 ;
			data[95428] <= 8'h10 ;
			data[95429] <= 8'h10 ;
			data[95430] <= 8'h10 ;
			data[95431] <= 8'h10 ;
			data[95432] <= 8'h10 ;
			data[95433] <= 8'h10 ;
			data[95434] <= 8'h10 ;
			data[95435] <= 8'h10 ;
			data[95436] <= 8'h10 ;
			data[95437] <= 8'h10 ;
			data[95438] <= 8'h10 ;
			data[95439] <= 8'h10 ;
			data[95440] <= 8'h10 ;
			data[95441] <= 8'h10 ;
			data[95442] <= 8'h10 ;
			data[95443] <= 8'h10 ;
			data[95444] <= 8'h10 ;
			data[95445] <= 8'h10 ;
			data[95446] <= 8'h10 ;
			data[95447] <= 8'h10 ;
			data[95448] <= 8'h10 ;
			data[95449] <= 8'h10 ;
			data[95450] <= 8'h10 ;
			data[95451] <= 8'h10 ;
			data[95452] <= 8'h10 ;
			data[95453] <= 8'h10 ;
			data[95454] <= 8'h10 ;
			data[95455] <= 8'h10 ;
			data[95456] <= 8'h10 ;
			data[95457] <= 8'h10 ;
			data[95458] <= 8'h10 ;
			data[95459] <= 8'h10 ;
			data[95460] <= 8'h10 ;
			data[95461] <= 8'h10 ;
			data[95462] <= 8'h10 ;
			data[95463] <= 8'h10 ;
			data[95464] <= 8'h10 ;
			data[95465] <= 8'h10 ;
			data[95466] <= 8'h10 ;
			data[95467] <= 8'h10 ;
			data[95468] <= 8'h10 ;
			data[95469] <= 8'h10 ;
			data[95470] <= 8'h10 ;
			data[95471] <= 8'h10 ;
			data[95472] <= 8'h10 ;
			data[95473] <= 8'h10 ;
			data[95474] <= 8'h10 ;
			data[95475] <= 8'h10 ;
			data[95476] <= 8'h10 ;
			data[95477] <= 8'h10 ;
			data[95478] <= 8'h10 ;
			data[95479] <= 8'h10 ;
			data[95480] <= 8'h10 ;
			data[95481] <= 8'h10 ;
			data[95482] <= 8'h10 ;
			data[95483] <= 8'h10 ;
			data[95484] <= 8'h10 ;
			data[95485] <= 8'h10 ;
			data[95486] <= 8'h10 ;
			data[95487] <= 8'h10 ;
			data[95488] <= 8'h10 ;
			data[95489] <= 8'h10 ;
			data[95490] <= 8'h10 ;
			data[95491] <= 8'h10 ;
			data[95492] <= 8'h10 ;
			data[95493] <= 8'h10 ;
			data[95494] <= 8'h10 ;
			data[95495] <= 8'h10 ;
			data[95496] <= 8'h10 ;
			data[95497] <= 8'h10 ;
			data[95498] <= 8'h10 ;
			data[95499] <= 8'h10 ;
			data[95500] <= 8'h10 ;
			data[95501] <= 8'h10 ;
			data[95502] <= 8'h10 ;
			data[95503] <= 8'h10 ;
			data[95504] <= 8'h10 ;
			data[95505] <= 8'h10 ;
			data[95506] <= 8'h10 ;
			data[95507] <= 8'h10 ;
			data[95508] <= 8'h10 ;
			data[95509] <= 8'h10 ;
			data[95510] <= 8'h10 ;
			data[95511] <= 8'h10 ;
			data[95512] <= 8'h10 ;
			data[95513] <= 8'h10 ;
			data[95514] <= 8'h10 ;
			data[95515] <= 8'h10 ;
			data[95516] <= 8'h10 ;
			data[95517] <= 8'h10 ;
			data[95518] <= 8'h10 ;
			data[95519] <= 8'h10 ;
			data[95520] <= 8'h10 ;
			data[95521] <= 8'h10 ;
			data[95522] <= 8'h10 ;
			data[95523] <= 8'h10 ;
			data[95524] <= 8'h10 ;
			data[95525] <= 8'h10 ;
			data[95526] <= 8'h10 ;
			data[95527] <= 8'h10 ;
			data[95528] <= 8'h10 ;
			data[95529] <= 8'h10 ;
			data[95530] <= 8'h10 ;
			data[95531] <= 8'h10 ;
			data[95532] <= 8'h10 ;
			data[95533] <= 8'h10 ;
			data[95534] <= 8'h10 ;
			data[95535] <= 8'h10 ;
			data[95536] <= 8'h10 ;
			data[95537] <= 8'h10 ;
			data[95538] <= 8'h10 ;
			data[95539] <= 8'h10 ;
			data[95540] <= 8'h10 ;
			data[95541] <= 8'h10 ;
			data[95542] <= 8'h10 ;
			data[95543] <= 8'h10 ;
			data[95544] <= 8'h10 ;
			data[95545] <= 8'h10 ;
			data[95546] <= 8'h10 ;
			data[95547] <= 8'h10 ;
			data[95548] <= 8'h10 ;
			data[95549] <= 8'h10 ;
			data[95550] <= 8'h10 ;
			data[95551] <= 8'h10 ;
			data[95552] <= 8'h10 ;
			data[95553] <= 8'h10 ;
			data[95554] <= 8'h10 ;
			data[95555] <= 8'h10 ;
			data[95556] <= 8'h10 ;
			data[95557] <= 8'h10 ;
			data[95558] <= 8'h10 ;
			data[95559] <= 8'h10 ;
			data[95560] <= 8'h10 ;
			data[95561] <= 8'h10 ;
			data[95562] <= 8'h10 ;
			data[95563] <= 8'h10 ;
			data[95564] <= 8'h10 ;
			data[95565] <= 8'h10 ;
			data[95566] <= 8'h10 ;
			data[95567] <= 8'h10 ;
			data[95568] <= 8'h10 ;
			data[95569] <= 8'h10 ;
			data[95570] <= 8'h10 ;
			data[95571] <= 8'h10 ;
			data[95572] <= 8'h10 ;
			data[95573] <= 8'h10 ;
			data[95574] <= 8'h10 ;
			data[95575] <= 8'h10 ;
			data[95576] <= 8'h10 ;
			data[95577] <= 8'h10 ;
			data[95578] <= 8'h10 ;
			data[95579] <= 8'h10 ;
			data[95580] <= 8'h10 ;
			data[95581] <= 8'h10 ;
			data[95582] <= 8'h10 ;
			data[95583] <= 8'h10 ;
			data[95584] <= 8'h10 ;
			data[95585] <= 8'h10 ;
			data[95586] <= 8'h10 ;
			data[95587] <= 8'h10 ;
			data[95588] <= 8'h10 ;
			data[95589] <= 8'h10 ;
			data[95590] <= 8'h10 ;
			data[95591] <= 8'h10 ;
			data[95592] <= 8'h10 ;
			data[95593] <= 8'h10 ;
			data[95594] <= 8'h10 ;
			data[95595] <= 8'h10 ;
			data[95596] <= 8'h10 ;
			data[95597] <= 8'h10 ;
			data[95598] <= 8'h10 ;
			data[95599] <= 8'h10 ;
			data[95600] <= 8'h10 ;
			data[95601] <= 8'h10 ;
			data[95602] <= 8'h10 ;
			data[95603] <= 8'h10 ;
			data[95604] <= 8'h10 ;
			data[95605] <= 8'h10 ;
			data[95606] <= 8'h10 ;
			data[95607] <= 8'h10 ;
			data[95608] <= 8'h10 ;
			data[95609] <= 8'h10 ;
			data[95610] <= 8'h10 ;
			data[95611] <= 8'h10 ;
			data[95612] <= 8'h10 ;
			data[95613] <= 8'h10 ;
			data[95614] <= 8'h10 ;
			data[95615] <= 8'h10 ;
			data[95616] <= 8'h10 ;
			data[95617] <= 8'h10 ;
			data[95618] <= 8'h10 ;
			data[95619] <= 8'h10 ;
			data[95620] <= 8'h10 ;
			data[95621] <= 8'h10 ;
			data[95622] <= 8'h10 ;
			data[95623] <= 8'h10 ;
			data[95624] <= 8'h10 ;
			data[95625] <= 8'h10 ;
			data[95626] <= 8'h10 ;
			data[95627] <= 8'h10 ;
			data[95628] <= 8'h10 ;
			data[95629] <= 8'h10 ;
			data[95630] <= 8'h10 ;
			data[95631] <= 8'h10 ;
			data[95632] <= 8'h10 ;
			data[95633] <= 8'h10 ;
			data[95634] <= 8'h10 ;
			data[95635] <= 8'h10 ;
			data[95636] <= 8'h10 ;
			data[95637] <= 8'h10 ;
			data[95638] <= 8'h10 ;
			data[95639] <= 8'h10 ;
			data[95640] <= 8'h10 ;
			data[95641] <= 8'h10 ;
			data[95642] <= 8'h10 ;
			data[95643] <= 8'h10 ;
			data[95644] <= 8'h10 ;
			data[95645] <= 8'h10 ;
			data[95646] <= 8'h10 ;
			data[95647] <= 8'h10 ;
			data[95648] <= 8'h10 ;
			data[95649] <= 8'h10 ;
			data[95650] <= 8'h10 ;
			data[95651] <= 8'h10 ;
			data[95652] <= 8'h10 ;
			data[95653] <= 8'h10 ;
			data[95654] <= 8'h10 ;
			data[95655] <= 8'h10 ;
			data[95656] <= 8'h10 ;
			data[95657] <= 8'h10 ;
			data[95658] <= 8'h10 ;
			data[95659] <= 8'h10 ;
			data[95660] <= 8'h10 ;
			data[95661] <= 8'h10 ;
			data[95662] <= 8'h10 ;
			data[95663] <= 8'h10 ;
			data[95664] <= 8'h10 ;
			data[95665] <= 8'h10 ;
			data[95666] <= 8'h10 ;
			data[95667] <= 8'h10 ;
			data[95668] <= 8'h10 ;
			data[95669] <= 8'h10 ;
			data[95670] <= 8'h10 ;
			data[95671] <= 8'h10 ;
			data[95672] <= 8'h10 ;
			data[95673] <= 8'h10 ;
			data[95674] <= 8'h10 ;
			data[95675] <= 8'h10 ;
			data[95676] <= 8'h10 ;
			data[95677] <= 8'h10 ;
			data[95678] <= 8'h10 ;
			data[95679] <= 8'h10 ;
			data[95680] <= 8'h10 ;
			data[95681] <= 8'h10 ;
			data[95682] <= 8'h10 ;
			data[95683] <= 8'h10 ;
			data[95684] <= 8'h10 ;
			data[95685] <= 8'h10 ;
			data[95686] <= 8'h10 ;
			data[95687] <= 8'h10 ;
			data[95688] <= 8'h10 ;
			data[95689] <= 8'h10 ;
			data[95690] <= 8'h10 ;
			data[95691] <= 8'h10 ;
			data[95692] <= 8'h10 ;
			data[95693] <= 8'h10 ;
			data[95694] <= 8'h10 ;
			data[95695] <= 8'h10 ;
			data[95696] <= 8'h10 ;
			data[95697] <= 8'h10 ;
			data[95698] <= 8'h10 ;
			data[95699] <= 8'h10 ;
			data[95700] <= 8'h10 ;
			data[95701] <= 8'h10 ;
			data[95702] <= 8'h10 ;
			data[95703] <= 8'h10 ;
			data[95704] <= 8'h10 ;
			data[95705] <= 8'h10 ;
			data[95706] <= 8'h10 ;
			data[95707] <= 8'h10 ;
			data[95708] <= 8'h10 ;
			data[95709] <= 8'h10 ;
			data[95710] <= 8'h10 ;
			data[95711] <= 8'h10 ;
			data[95712] <= 8'h10 ;
			data[95713] <= 8'h10 ;
			data[95714] <= 8'h10 ;
			data[95715] <= 8'h10 ;
			data[95716] <= 8'h10 ;
			data[95717] <= 8'h10 ;
			data[95718] <= 8'h10 ;
			data[95719] <= 8'h10 ;
			data[95720] <= 8'h10 ;
			data[95721] <= 8'h10 ;
			data[95722] <= 8'h10 ;
			data[95723] <= 8'h10 ;
			data[95724] <= 8'h10 ;
			data[95725] <= 8'h10 ;
			data[95726] <= 8'h10 ;
			data[95727] <= 8'h10 ;
			data[95728] <= 8'h10 ;
			data[95729] <= 8'h10 ;
			data[95730] <= 8'h10 ;
			data[95731] <= 8'h10 ;
			data[95732] <= 8'h10 ;
			data[95733] <= 8'h10 ;
			data[95734] <= 8'h10 ;
			data[95735] <= 8'h10 ;
			data[95736] <= 8'h10 ;
			data[95737] <= 8'h10 ;
			data[95738] <= 8'h10 ;
			data[95739] <= 8'h10 ;
			data[95740] <= 8'h10 ;
			data[95741] <= 8'h10 ;
			data[95742] <= 8'h10 ;
			data[95743] <= 8'h10 ;
			data[95744] <= 8'h10 ;
			data[95745] <= 8'h10 ;
			data[95746] <= 8'h10 ;
			data[95747] <= 8'h10 ;
			data[95748] <= 8'h10 ;
			data[95749] <= 8'h10 ;
			data[95750] <= 8'h10 ;
			data[95751] <= 8'h10 ;
			data[95752] <= 8'h10 ;
			data[95753] <= 8'h10 ;
			data[95754] <= 8'h10 ;
			data[95755] <= 8'h10 ;
			data[95756] <= 8'h10 ;
			data[95757] <= 8'h10 ;
			data[95758] <= 8'h10 ;
			data[95759] <= 8'h10 ;
			data[95760] <= 8'h10 ;
			data[95761] <= 8'h10 ;
			data[95762] <= 8'h10 ;
			data[95763] <= 8'h10 ;
			data[95764] <= 8'h10 ;
			data[95765] <= 8'h10 ;
			data[95766] <= 8'h10 ;
			data[95767] <= 8'h10 ;
			data[95768] <= 8'h10 ;
			data[95769] <= 8'h10 ;
			data[95770] <= 8'h10 ;
			data[95771] <= 8'h10 ;
			data[95772] <= 8'h10 ;
			data[95773] <= 8'h10 ;
			data[95774] <= 8'h10 ;
			data[95775] <= 8'h10 ;
			data[95776] <= 8'h10 ;
			data[95777] <= 8'h10 ;
			data[95778] <= 8'h10 ;
			data[95779] <= 8'h10 ;
			data[95780] <= 8'h10 ;
			data[95781] <= 8'h10 ;
			data[95782] <= 8'h10 ;
			data[95783] <= 8'h10 ;
			data[95784] <= 8'h10 ;
			data[95785] <= 8'h10 ;
			data[95786] <= 8'h10 ;
			data[95787] <= 8'h10 ;
			data[95788] <= 8'h10 ;
			data[95789] <= 8'h10 ;
			data[95790] <= 8'h10 ;
			data[95791] <= 8'h10 ;
			data[95792] <= 8'h10 ;
			data[95793] <= 8'h10 ;
			data[95794] <= 8'h10 ;
			data[95795] <= 8'h10 ;
			data[95796] <= 8'h10 ;
			data[95797] <= 8'h10 ;
			data[95798] <= 8'h10 ;
			data[95799] <= 8'h10 ;
			data[95800] <= 8'h10 ;
			data[95801] <= 8'h10 ;
			data[95802] <= 8'h10 ;
			data[95803] <= 8'h10 ;
			data[95804] <= 8'h10 ;
			data[95805] <= 8'h10 ;
			data[95806] <= 8'h10 ;
			data[95807] <= 8'h10 ;
			data[95808] <= 8'h10 ;
			data[95809] <= 8'h10 ;
			data[95810] <= 8'h10 ;
			data[95811] <= 8'h10 ;
			data[95812] <= 8'h10 ;
			data[95813] <= 8'h10 ;
			data[95814] <= 8'h10 ;
			data[95815] <= 8'h10 ;
			data[95816] <= 8'h10 ;
			data[95817] <= 8'h10 ;
			data[95818] <= 8'h10 ;
			data[95819] <= 8'h10 ;
			data[95820] <= 8'h10 ;
			data[95821] <= 8'h10 ;
			data[95822] <= 8'h10 ;
			data[95823] <= 8'h10 ;
			data[95824] <= 8'h10 ;
			data[95825] <= 8'h10 ;
			data[95826] <= 8'h10 ;
			data[95827] <= 8'h10 ;
			data[95828] <= 8'h10 ;
			data[95829] <= 8'h10 ;
			data[95830] <= 8'h10 ;
			data[95831] <= 8'h10 ;
			data[95832] <= 8'h10 ;
			data[95833] <= 8'h10 ;
			data[95834] <= 8'h10 ;
			data[95835] <= 8'h10 ;
			data[95836] <= 8'h10 ;
			data[95837] <= 8'h10 ;
			data[95838] <= 8'h10 ;
			data[95839] <= 8'h10 ;
			data[95840] <= 8'h10 ;
			data[95841] <= 8'h10 ;
			data[95842] <= 8'h10 ;
			data[95843] <= 8'h10 ;
			data[95844] <= 8'h10 ;
			data[95845] <= 8'h10 ;
			data[95846] <= 8'h10 ;
			data[95847] <= 8'h10 ;
			data[95848] <= 8'h10 ;
			data[95849] <= 8'h10 ;
			data[95850] <= 8'h10 ;
			data[95851] <= 8'h10 ;
			data[95852] <= 8'h10 ;
			data[95853] <= 8'h10 ;
			data[95854] <= 8'h10 ;
			data[95855] <= 8'h10 ;
			data[95856] <= 8'h10 ;
			data[95857] <= 8'h10 ;
			data[95858] <= 8'h10 ;
			data[95859] <= 8'h10 ;
			data[95860] <= 8'h10 ;
			data[95861] <= 8'h10 ;
			data[95862] <= 8'h10 ;
			data[95863] <= 8'h10 ;
			data[95864] <= 8'h10 ;
			data[95865] <= 8'h10 ;
			data[95866] <= 8'h10 ;
			data[95867] <= 8'h10 ;
			data[95868] <= 8'h10 ;
			data[95869] <= 8'h10 ;
			data[95870] <= 8'h10 ;
			data[95871] <= 8'h10 ;
			data[95872] <= 8'h10 ;
			data[95873] <= 8'h10 ;
			data[95874] <= 8'h10 ;
			data[95875] <= 8'h10 ;
			data[95876] <= 8'h10 ;
			data[95877] <= 8'h10 ;
			data[95878] <= 8'h10 ;
			data[95879] <= 8'h10 ;
			data[95880] <= 8'h10 ;
			data[95881] <= 8'h10 ;
			data[95882] <= 8'h10 ;
			data[95883] <= 8'h10 ;
			data[95884] <= 8'h10 ;
			data[95885] <= 8'h10 ;
			data[95886] <= 8'h10 ;
			data[95887] <= 8'h10 ;
			data[95888] <= 8'h10 ;
			data[95889] <= 8'h10 ;
			data[95890] <= 8'h10 ;
			data[95891] <= 8'h10 ;
			data[95892] <= 8'h10 ;
			data[95893] <= 8'h10 ;
			data[95894] <= 8'h10 ;
			data[95895] <= 8'h10 ;
			data[95896] <= 8'h10 ;
			data[95897] <= 8'h10 ;
			data[95898] <= 8'h10 ;
			data[95899] <= 8'h10 ;
			data[95900] <= 8'h10 ;
			data[95901] <= 8'h10 ;
			data[95902] <= 8'h10 ;
			data[95903] <= 8'h10 ;
			data[95904] <= 8'h10 ;
			data[95905] <= 8'h10 ;
			data[95906] <= 8'h10 ;
			data[95907] <= 8'h10 ;
			data[95908] <= 8'h10 ;
			data[95909] <= 8'h10 ;
			data[95910] <= 8'h10 ;
			data[95911] <= 8'h10 ;
			data[95912] <= 8'h10 ;
			data[95913] <= 8'h10 ;
			data[95914] <= 8'h10 ;
			data[95915] <= 8'h10 ;
			data[95916] <= 8'h10 ;
			data[95917] <= 8'h10 ;
			data[95918] <= 8'h10 ;
			data[95919] <= 8'h10 ;
			data[95920] <= 8'h10 ;
			data[95921] <= 8'h10 ;
			data[95922] <= 8'h10 ;
			data[95923] <= 8'h10 ;
			data[95924] <= 8'h10 ;
			data[95925] <= 8'h10 ;
			data[95926] <= 8'h10 ;
			data[95927] <= 8'h10 ;
			data[95928] <= 8'h10 ;
			data[95929] <= 8'h10 ;
			data[95930] <= 8'h10 ;
			data[95931] <= 8'h10 ;
			data[95932] <= 8'h10 ;
			data[95933] <= 8'h10 ;
			data[95934] <= 8'h10 ;
			data[95935] <= 8'h10 ;
			data[95936] <= 8'h10 ;
			data[95937] <= 8'h10 ;
			data[95938] <= 8'h10 ;
			data[95939] <= 8'h10 ;
			data[95940] <= 8'h10 ;
			data[95941] <= 8'h10 ;
			data[95942] <= 8'h10 ;
			data[95943] <= 8'h10 ;
			data[95944] <= 8'h10 ;
			data[95945] <= 8'h10 ;
			data[95946] <= 8'h10 ;
			data[95947] <= 8'h10 ;
			data[95948] <= 8'h10 ;
			data[95949] <= 8'h10 ;
			data[95950] <= 8'h10 ;
			data[95951] <= 8'h10 ;
			data[95952] <= 8'h10 ;
			data[95953] <= 8'h10 ;
			data[95954] <= 8'h10 ;
			data[95955] <= 8'h10 ;
			data[95956] <= 8'h10 ;
			data[95957] <= 8'h10 ;
			data[95958] <= 8'h10 ;
			data[95959] <= 8'h10 ;
			data[95960] <= 8'h10 ;
			data[95961] <= 8'h10 ;
			data[95962] <= 8'h10 ;
			data[95963] <= 8'h10 ;
			data[95964] <= 8'h10 ;
			data[95965] <= 8'h10 ;
			data[95966] <= 8'h10 ;
			data[95967] <= 8'h10 ;
			data[95968] <= 8'h10 ;
			data[95969] <= 8'h10 ;
			data[95970] <= 8'h10 ;
			data[95971] <= 8'h10 ;
			data[95972] <= 8'h10 ;
			data[95973] <= 8'h10 ;
			data[95974] <= 8'h10 ;
			data[95975] <= 8'h10 ;
			data[95976] <= 8'h10 ;
			data[95977] <= 8'h10 ;
			data[95978] <= 8'h10 ;
			data[95979] <= 8'h10 ;
			data[95980] <= 8'h10 ;
			data[95981] <= 8'h10 ;
			data[95982] <= 8'h10 ;
			data[95983] <= 8'h10 ;
			data[95984] <= 8'h10 ;
			data[95985] <= 8'h10 ;
			data[95986] <= 8'h10 ;
			data[95987] <= 8'h10 ;
			data[95988] <= 8'h10 ;
			data[95989] <= 8'h10 ;
			data[95990] <= 8'h10 ;
			data[95991] <= 8'h10 ;
			data[95992] <= 8'h10 ;
			data[95993] <= 8'h10 ;
			data[95994] <= 8'h10 ;
			data[95995] <= 8'h10 ;
			data[95996] <= 8'h10 ;
			data[95997] <= 8'h10 ;
			data[95998] <= 8'h10 ;
			data[95999] <= 8'h10 ;
			data[96000] <= 8'h10 ;
			data[96001] <= 8'h10 ;
			data[96002] <= 8'h10 ;
			data[96003] <= 8'h10 ;
			data[96004] <= 8'h10 ;
			data[96005] <= 8'h10 ;
			data[96006] <= 8'h10 ;
			data[96007] <= 8'h10 ;
			data[96008] <= 8'h10 ;
			data[96009] <= 8'h10 ;
			data[96010] <= 8'h10 ;
			data[96011] <= 8'h10 ;
			data[96012] <= 8'h10 ;
			data[96013] <= 8'h10 ;
			data[96014] <= 8'h10 ;
			data[96015] <= 8'h10 ;
			data[96016] <= 8'h10 ;
			data[96017] <= 8'h10 ;
			data[96018] <= 8'h10 ;
			data[96019] <= 8'h10 ;
			data[96020] <= 8'h10 ;
			data[96021] <= 8'h10 ;
			data[96022] <= 8'h10 ;
			data[96023] <= 8'h10 ;
			data[96024] <= 8'h10 ;
			data[96025] <= 8'h10 ;
			data[96026] <= 8'h10 ;
			data[96027] <= 8'h10 ;
			data[96028] <= 8'h10 ;
			data[96029] <= 8'h10 ;
			data[96030] <= 8'h10 ;
			data[96031] <= 8'h10 ;
			data[96032] <= 8'h10 ;
			data[96033] <= 8'h10 ;
			data[96034] <= 8'h10 ;
			data[96035] <= 8'h10 ;
			data[96036] <= 8'h10 ;
			data[96037] <= 8'h10 ;
			data[96038] <= 8'h10 ;
			data[96039] <= 8'h10 ;
			data[96040] <= 8'h10 ;
			data[96041] <= 8'h10 ;
			data[96042] <= 8'h10 ;
			data[96043] <= 8'h10 ;
			data[96044] <= 8'h10 ;
			data[96045] <= 8'h10 ;
			data[96046] <= 8'h10 ;
			data[96047] <= 8'h10 ;
			data[96048] <= 8'h10 ;
			data[96049] <= 8'h10 ;
			data[96050] <= 8'h10 ;
			data[96051] <= 8'h10 ;
			data[96052] <= 8'h10 ;
			data[96053] <= 8'h10 ;
			data[96054] <= 8'h10 ;
			data[96055] <= 8'h10 ;
			data[96056] <= 8'h10 ;
			data[96057] <= 8'h10 ;
			data[96058] <= 8'h10 ;
			data[96059] <= 8'h10 ;
			data[96060] <= 8'h10 ;
			data[96061] <= 8'h10 ;
			data[96062] <= 8'h10 ;
			data[96063] <= 8'h10 ;
			data[96064] <= 8'h10 ;
			data[96065] <= 8'h10 ;
			data[96066] <= 8'h10 ;
			data[96067] <= 8'h10 ;
			data[96068] <= 8'h10 ;
			data[96069] <= 8'h10 ;
			data[96070] <= 8'h10 ;
			data[96071] <= 8'h10 ;
			data[96072] <= 8'h10 ;
			data[96073] <= 8'h10 ;
			data[96074] <= 8'h10 ;
			data[96075] <= 8'h10 ;
			data[96076] <= 8'h10 ;
			data[96077] <= 8'h10 ;
			data[96078] <= 8'h10 ;
			data[96079] <= 8'h10 ;
			data[96080] <= 8'h10 ;
			data[96081] <= 8'h10 ;
			data[96082] <= 8'h10 ;
			data[96083] <= 8'h10 ;
			data[96084] <= 8'h10 ;
			data[96085] <= 8'h10 ;
			data[96086] <= 8'h10 ;
			data[96087] <= 8'h10 ;
			data[96088] <= 8'h10 ;
			data[96089] <= 8'h10 ;
			data[96090] <= 8'h10 ;
			data[96091] <= 8'h10 ;
			data[96092] <= 8'h10 ;
			data[96093] <= 8'h10 ;
			data[96094] <= 8'h10 ;
			data[96095] <= 8'h10 ;
			data[96096] <= 8'h10 ;
			data[96097] <= 8'h10 ;
			data[96098] <= 8'h10 ;
			data[96099] <= 8'h10 ;
			data[96100] <= 8'h10 ;
			data[96101] <= 8'h10 ;
			data[96102] <= 8'h10 ;
			data[96103] <= 8'h10 ;
			data[96104] <= 8'h10 ;
			data[96105] <= 8'h10 ;
			data[96106] <= 8'h10 ;
			data[96107] <= 8'h10 ;
			data[96108] <= 8'h10 ;
			data[96109] <= 8'h10 ;
			data[96110] <= 8'h10 ;
			data[96111] <= 8'h10 ;
			data[96112] <= 8'h10 ;
			data[96113] <= 8'h10 ;
			data[96114] <= 8'h10 ;
			data[96115] <= 8'h10 ;
			data[96116] <= 8'h10 ;
			data[96117] <= 8'h10 ;
			data[96118] <= 8'h10 ;
			data[96119] <= 8'h10 ;
			data[96120] <= 8'h10 ;
			data[96121] <= 8'h10 ;
			data[96122] <= 8'h10 ;
			data[96123] <= 8'h10 ;
			data[96124] <= 8'h10 ;
			data[96125] <= 8'h10 ;
			data[96126] <= 8'h10 ;
			data[96127] <= 8'h10 ;
			data[96128] <= 8'h10 ;
			data[96129] <= 8'h10 ;
			data[96130] <= 8'h10 ;
			data[96131] <= 8'h10 ;
			data[96132] <= 8'h10 ;
			data[96133] <= 8'h10 ;
			data[96134] <= 8'h10 ;
			data[96135] <= 8'h10 ;
			data[96136] <= 8'h10 ;
			data[96137] <= 8'h10 ;
			data[96138] <= 8'h10 ;
			data[96139] <= 8'h10 ;
			data[96140] <= 8'h10 ;
			data[96141] <= 8'h10 ;
			data[96142] <= 8'h10 ;
			data[96143] <= 8'h10 ;
			data[96144] <= 8'h10 ;
			data[96145] <= 8'h10 ;
			data[96146] <= 8'h10 ;
			data[96147] <= 8'h10 ;
			data[96148] <= 8'h10 ;
			data[96149] <= 8'h10 ;
			data[96150] <= 8'h10 ;
			data[96151] <= 8'h10 ;
			data[96152] <= 8'h10 ;
			data[96153] <= 8'h10 ;
			data[96154] <= 8'h10 ;
			data[96155] <= 8'h10 ;
			data[96156] <= 8'h10 ;
			data[96157] <= 8'h10 ;
			data[96158] <= 8'h10 ;
			data[96159] <= 8'h10 ;
			data[96160] <= 8'h10 ;
			data[96161] <= 8'h10 ;
			data[96162] <= 8'h10 ;
			data[96163] <= 8'h10 ;
			data[96164] <= 8'h10 ;
			data[96165] <= 8'h10 ;
			data[96166] <= 8'h10 ;
			data[96167] <= 8'h10 ;
			data[96168] <= 8'h10 ;
			data[96169] <= 8'h10 ;
			data[96170] <= 8'h10 ;
			data[96171] <= 8'h10 ;
			data[96172] <= 8'h10 ;
			data[96173] <= 8'h10 ;
			data[96174] <= 8'h10 ;
			data[96175] <= 8'h10 ;
			data[96176] <= 8'h10 ;
			data[96177] <= 8'h10 ;
			data[96178] <= 8'h10 ;
			data[96179] <= 8'h10 ;
			data[96180] <= 8'h10 ;
			data[96181] <= 8'h10 ;
			data[96182] <= 8'h10 ;
			data[96183] <= 8'h10 ;
			data[96184] <= 8'h10 ;
			data[96185] <= 8'h10 ;
			data[96186] <= 8'h10 ;
			data[96187] <= 8'h10 ;
			data[96188] <= 8'h10 ;
			data[96189] <= 8'h10 ;
			data[96190] <= 8'h10 ;
			data[96191] <= 8'h10 ;
			data[96192] <= 8'h10 ;
			data[96193] <= 8'h10 ;
			data[96194] <= 8'h10 ;
			data[96195] <= 8'h10 ;
			data[96196] <= 8'h10 ;
			data[96197] <= 8'h10 ;
			data[96198] <= 8'h10 ;
			data[96199] <= 8'h10 ;
			data[96200] <= 8'h10 ;
			data[96201] <= 8'h10 ;
			data[96202] <= 8'h10 ;
			data[96203] <= 8'h10 ;
			data[96204] <= 8'h10 ;
			data[96205] <= 8'h10 ;
			data[96206] <= 8'h10 ;
			data[96207] <= 8'h10 ;
			data[96208] <= 8'h10 ;
			data[96209] <= 8'h10 ;
			data[96210] <= 8'h10 ;
			data[96211] <= 8'h10 ;
			data[96212] <= 8'h10 ;
			data[96213] <= 8'h10 ;
			data[96214] <= 8'h10 ;
			data[96215] <= 8'h10 ;
			data[96216] <= 8'h10 ;
			data[96217] <= 8'h10 ;
			data[96218] <= 8'h10 ;
			data[96219] <= 8'h10 ;
			data[96220] <= 8'h10 ;
			data[96221] <= 8'h10 ;
			data[96222] <= 8'h10 ;
			data[96223] <= 8'h10 ;
			data[96224] <= 8'h10 ;
			data[96225] <= 8'h10 ;
			data[96226] <= 8'h10 ;
			data[96227] <= 8'h10 ;
			data[96228] <= 8'h10 ;
			data[96229] <= 8'h10 ;
			data[96230] <= 8'h10 ;
			data[96231] <= 8'h10 ;
			data[96232] <= 8'h10 ;
			data[96233] <= 8'h10 ;
			data[96234] <= 8'h10 ;
			data[96235] <= 8'h10 ;
			data[96236] <= 8'h10 ;
			data[96237] <= 8'h10 ;
			data[96238] <= 8'h10 ;
			data[96239] <= 8'h10 ;
			data[96240] <= 8'h10 ;
			data[96241] <= 8'h10 ;
			data[96242] <= 8'h10 ;
			data[96243] <= 8'h10 ;
			data[96244] <= 8'h10 ;
			data[96245] <= 8'h10 ;
			data[96246] <= 8'h10 ;
			data[96247] <= 8'h10 ;
			data[96248] <= 8'h10 ;
			data[96249] <= 8'h10 ;
			data[96250] <= 8'h10 ;
			data[96251] <= 8'h10 ;
			data[96252] <= 8'h10 ;
			data[96253] <= 8'h10 ;
			data[96254] <= 8'h10 ;
			data[96255] <= 8'h10 ;
			data[96256] <= 8'h10 ;
			data[96257] <= 8'h10 ;
			data[96258] <= 8'h10 ;
			data[96259] <= 8'h10 ;
			data[96260] <= 8'h10 ;
			data[96261] <= 8'h10 ;
			data[96262] <= 8'h10 ;
			data[96263] <= 8'h10 ;
			data[96264] <= 8'h10 ;
			data[96265] <= 8'h10 ;
			data[96266] <= 8'h10 ;
			data[96267] <= 8'h10 ;
			data[96268] <= 8'h10 ;
			data[96269] <= 8'h10 ;
			data[96270] <= 8'h10 ;
			data[96271] <= 8'h10 ;
			data[96272] <= 8'h10 ;
			data[96273] <= 8'h10 ;
			data[96274] <= 8'h10 ;
			data[96275] <= 8'h10 ;
			data[96276] <= 8'h10 ;
			data[96277] <= 8'h10 ;
			data[96278] <= 8'h10 ;
			data[96279] <= 8'h10 ;
			data[96280] <= 8'h10 ;
			data[96281] <= 8'h10 ;
			data[96282] <= 8'h10 ;
			data[96283] <= 8'h10 ;
			data[96284] <= 8'h10 ;
			data[96285] <= 8'h10 ;
			data[96286] <= 8'h10 ;
			data[96287] <= 8'h10 ;
			data[96288] <= 8'h10 ;
			data[96289] <= 8'h10 ;
			data[96290] <= 8'h10 ;
			data[96291] <= 8'h10 ;
			data[96292] <= 8'h10 ;
			data[96293] <= 8'h10 ;
			data[96294] <= 8'h10 ;
			data[96295] <= 8'h10 ;
			data[96296] <= 8'h10 ;
			data[96297] <= 8'h10 ;
			data[96298] <= 8'h10 ;
			data[96299] <= 8'h10 ;
			data[96300] <= 8'h10 ;
			data[96301] <= 8'h10 ;
			data[96302] <= 8'h10 ;
			data[96303] <= 8'h10 ;
			data[96304] <= 8'h10 ;
			data[96305] <= 8'h10 ;
			data[96306] <= 8'h10 ;
			data[96307] <= 8'h10 ;
			data[96308] <= 8'h10 ;
			data[96309] <= 8'h10 ;
			data[96310] <= 8'h10 ;
			data[96311] <= 8'h10 ;
			data[96312] <= 8'h10 ;
			data[96313] <= 8'h10 ;
			data[96314] <= 8'h10 ;
			data[96315] <= 8'h10 ;
			data[96316] <= 8'h10 ;
			data[96317] <= 8'h10 ;
			data[96318] <= 8'h10 ;
			data[96319] <= 8'h10 ;
			data[96320] <= 8'h10 ;
			data[96321] <= 8'h10 ;
			data[96322] <= 8'h10 ;
			data[96323] <= 8'h10 ;
			data[96324] <= 8'h10 ;
			data[96325] <= 8'h10 ;
			data[96326] <= 8'h10 ;
			data[96327] <= 8'h10 ;
			data[96328] <= 8'h10 ;
			data[96329] <= 8'h10 ;
			data[96330] <= 8'h10 ;
			data[96331] <= 8'h10 ;
			data[96332] <= 8'h10 ;
			data[96333] <= 8'h10 ;
			data[96334] <= 8'h10 ;
			data[96335] <= 8'h10 ;
			data[96336] <= 8'h10 ;
			data[96337] <= 8'h10 ;
			data[96338] <= 8'h10 ;
			data[96339] <= 8'h10 ;
			data[96340] <= 8'h10 ;
			data[96341] <= 8'h10 ;
			data[96342] <= 8'h10 ;
			data[96343] <= 8'h10 ;
			data[96344] <= 8'h10 ;
			data[96345] <= 8'h10 ;
			data[96346] <= 8'h10 ;
			data[96347] <= 8'h10 ;
			data[96348] <= 8'h10 ;
			data[96349] <= 8'h10 ;
			data[96350] <= 8'h10 ;
			data[96351] <= 8'h10 ;
			data[96352] <= 8'h10 ;
			data[96353] <= 8'h10 ;
			data[96354] <= 8'h10 ;
			data[96355] <= 8'h10 ;
			data[96356] <= 8'h10 ;
			data[96357] <= 8'h10 ;
			data[96358] <= 8'h10 ;
			data[96359] <= 8'h10 ;
			data[96360] <= 8'h10 ;
			data[96361] <= 8'h10 ;
			data[96362] <= 8'h10 ;
			data[96363] <= 8'h10 ;
			data[96364] <= 8'h10 ;
			data[96365] <= 8'h10 ;
			data[96366] <= 8'h10 ;
			data[96367] <= 8'h10 ;
			data[96368] <= 8'h10 ;
			data[96369] <= 8'h10 ;
			data[96370] <= 8'h10 ;
			data[96371] <= 8'h10 ;
			data[96372] <= 8'h10 ;
			data[96373] <= 8'h10 ;
			data[96374] <= 8'h10 ;
			data[96375] <= 8'h10 ;
			data[96376] <= 8'h10 ;
			data[96377] <= 8'h10 ;
			data[96378] <= 8'h10 ;
			data[96379] <= 8'h10 ;
			data[96380] <= 8'h10 ;
			data[96381] <= 8'h10 ;
			data[96382] <= 8'h10 ;
			data[96383] <= 8'h10 ;
			data[96384] <= 8'h10 ;
			data[96385] <= 8'h10 ;
			data[96386] <= 8'h10 ;
			data[96387] <= 8'h10 ;
			data[96388] <= 8'h10 ;
			data[96389] <= 8'h10 ;
			data[96390] <= 8'h10 ;
			data[96391] <= 8'h10 ;
			data[96392] <= 8'h10 ;
			data[96393] <= 8'h10 ;
			data[96394] <= 8'h10 ;
			data[96395] <= 8'h10 ;
			data[96396] <= 8'h10 ;
			data[96397] <= 8'h10 ;
			data[96398] <= 8'h10 ;
			data[96399] <= 8'h10 ;
			data[96400] <= 8'h10 ;
			data[96401] <= 8'h10 ;
			data[96402] <= 8'h10 ;
			data[96403] <= 8'h10 ;
			data[96404] <= 8'h10 ;
			data[96405] <= 8'h10 ;
			data[96406] <= 8'h10 ;
			data[96407] <= 8'h10 ;
			data[96408] <= 8'h10 ;
			data[96409] <= 8'h10 ;
			data[96410] <= 8'h10 ;
			data[96411] <= 8'h10 ;
			data[96412] <= 8'h10 ;
			data[96413] <= 8'h10 ;
			data[96414] <= 8'h10 ;
			data[96415] <= 8'h10 ;
			data[96416] <= 8'h10 ;
			data[96417] <= 8'h10 ;
			data[96418] <= 8'h10 ;
			data[96419] <= 8'h10 ;
			data[96420] <= 8'h10 ;
			data[96421] <= 8'h10 ;
			data[96422] <= 8'h10 ;
			data[96423] <= 8'h10 ;
			data[96424] <= 8'h10 ;
			data[96425] <= 8'h10 ;
			data[96426] <= 8'h10 ;
			data[96427] <= 8'h10 ;
			data[96428] <= 8'h10 ;
			data[96429] <= 8'h10 ;
			data[96430] <= 8'h10 ;
			data[96431] <= 8'h10 ;
			data[96432] <= 8'h10 ;
			data[96433] <= 8'h10 ;
			data[96434] <= 8'h10 ;
			data[96435] <= 8'h10 ;
			data[96436] <= 8'h10 ;
			data[96437] <= 8'h10 ;
			data[96438] <= 8'h10 ;
			data[96439] <= 8'h10 ;
			data[96440] <= 8'h10 ;
			data[96441] <= 8'h10 ;
			data[96442] <= 8'h10 ;
			data[96443] <= 8'h10 ;
			data[96444] <= 8'h10 ;
			data[96445] <= 8'h10 ;
			data[96446] <= 8'h10 ;
			data[96447] <= 8'h10 ;
			data[96448] <= 8'h10 ;
			data[96449] <= 8'h10 ;
			data[96450] <= 8'h10 ;
			data[96451] <= 8'h10 ;
			data[96452] <= 8'h10 ;
			data[96453] <= 8'h10 ;
			data[96454] <= 8'h10 ;
			data[96455] <= 8'h10 ;
			data[96456] <= 8'h10 ;
			data[96457] <= 8'h10 ;
			data[96458] <= 8'h10 ;
			data[96459] <= 8'h10 ;
			data[96460] <= 8'h10 ;
			data[96461] <= 8'h10 ;
			data[96462] <= 8'h10 ;
			data[96463] <= 8'h10 ;
			data[96464] <= 8'h10 ;
			data[96465] <= 8'h10 ;
			data[96466] <= 8'h10 ;
			data[96467] <= 8'h10 ;
			data[96468] <= 8'h10 ;
			data[96469] <= 8'h10 ;
			data[96470] <= 8'h10 ;
			data[96471] <= 8'h10 ;
			data[96472] <= 8'h10 ;
			data[96473] <= 8'h10 ;
			data[96474] <= 8'h10 ;
			data[96475] <= 8'h10 ;
			data[96476] <= 8'h10 ;
			data[96477] <= 8'h10 ;
			data[96478] <= 8'h10 ;
			data[96479] <= 8'h10 ;
			data[96480] <= 8'h10 ;
			data[96481] <= 8'h10 ;
			data[96482] <= 8'h10 ;
			data[96483] <= 8'h10 ;
			data[96484] <= 8'h10 ;
			data[96485] <= 8'h10 ;
			data[96486] <= 8'h10 ;
			data[96487] <= 8'h10 ;
			data[96488] <= 8'h10 ;
			data[96489] <= 8'h10 ;
			data[96490] <= 8'h10 ;
			data[96491] <= 8'h10 ;
			data[96492] <= 8'h10 ;
			data[96493] <= 8'h10 ;
			data[96494] <= 8'h10 ;
			data[96495] <= 8'h10 ;
			data[96496] <= 8'h10 ;
			data[96497] <= 8'h10 ;
			data[96498] <= 8'h10 ;
			data[96499] <= 8'h10 ;
			data[96500] <= 8'h10 ;
			data[96501] <= 8'h10 ;
			data[96502] <= 8'h10 ;
			data[96503] <= 8'h10 ;
			data[96504] <= 8'h10 ;
			data[96505] <= 8'h10 ;
			data[96506] <= 8'h10 ;
			data[96507] <= 8'h10 ;
			data[96508] <= 8'h10 ;
			data[96509] <= 8'h10 ;
			data[96510] <= 8'h10 ;
			data[96511] <= 8'h10 ;
			data[96512] <= 8'h10 ;
			data[96513] <= 8'h10 ;
			data[96514] <= 8'h10 ;
			data[96515] <= 8'h10 ;
			data[96516] <= 8'h10 ;
			data[96517] <= 8'h10 ;
			data[96518] <= 8'h10 ;
			data[96519] <= 8'h10 ;
			data[96520] <= 8'h10 ;
			data[96521] <= 8'h10 ;
			data[96522] <= 8'h10 ;
			data[96523] <= 8'h10 ;
			data[96524] <= 8'h10 ;
			data[96525] <= 8'h10 ;
			data[96526] <= 8'h10 ;
			data[96527] <= 8'h10 ;
			data[96528] <= 8'h10 ;
			data[96529] <= 8'h10 ;
			data[96530] <= 8'h10 ;
			data[96531] <= 8'h10 ;
			data[96532] <= 8'h10 ;
			data[96533] <= 8'h10 ;
			data[96534] <= 8'h10 ;
			data[96535] <= 8'h10 ;
			data[96536] <= 8'h10 ;
			data[96537] <= 8'h10 ;
			data[96538] <= 8'h10 ;
			data[96539] <= 8'h10 ;
			data[96540] <= 8'h10 ;
			data[96541] <= 8'h10 ;
			data[96542] <= 8'h10 ;
			data[96543] <= 8'h10 ;
			data[96544] <= 8'h10 ;
			data[96545] <= 8'h10 ;
			data[96546] <= 8'h10 ;
			data[96547] <= 8'h10 ;
			data[96548] <= 8'h10 ;
			data[96549] <= 8'h10 ;
			data[96550] <= 8'h10 ;
			data[96551] <= 8'h10 ;
			data[96552] <= 8'h10 ;
			data[96553] <= 8'h10 ;
			data[96554] <= 8'h10 ;
			data[96555] <= 8'h10 ;
			data[96556] <= 8'h10 ;
			data[96557] <= 8'h10 ;
			data[96558] <= 8'h10 ;
			data[96559] <= 8'h10 ;
			data[96560] <= 8'h10 ;
			data[96561] <= 8'h10 ;
			data[96562] <= 8'h10 ;
			data[96563] <= 8'h10 ;
			data[96564] <= 8'h10 ;
			data[96565] <= 8'h10 ;
			data[96566] <= 8'h10 ;
			data[96567] <= 8'h10 ;
			data[96568] <= 8'h10 ;
			data[96569] <= 8'h10 ;
			data[96570] <= 8'h10 ;
			data[96571] <= 8'h10 ;
			data[96572] <= 8'h10 ;
			data[96573] <= 8'h10 ;
			data[96574] <= 8'h10 ;
			data[96575] <= 8'h10 ;
			data[96576] <= 8'h10 ;
			data[96577] <= 8'h10 ;
			data[96578] <= 8'h10 ;
			data[96579] <= 8'h10 ;
			data[96580] <= 8'h10 ;
			data[96581] <= 8'h10 ;
			data[96582] <= 8'h10 ;
			data[96583] <= 8'h10 ;
			data[96584] <= 8'h10 ;
			data[96585] <= 8'h10 ;
			data[96586] <= 8'h10 ;
			data[96587] <= 8'h10 ;
			data[96588] <= 8'h10 ;
			data[96589] <= 8'h10 ;
			data[96590] <= 8'h10 ;
			data[96591] <= 8'h10 ;
			data[96592] <= 8'h10 ;
			data[96593] <= 8'h10 ;
			data[96594] <= 8'h10 ;
			data[96595] <= 8'h10 ;
			data[96596] <= 8'h10 ;
			data[96597] <= 8'h10 ;
			data[96598] <= 8'h10 ;
			data[96599] <= 8'h10 ;
			data[96600] <= 8'h10 ;
			data[96601] <= 8'h10 ;
			data[96602] <= 8'h10 ;
			data[96603] <= 8'h10 ;
			data[96604] <= 8'h10 ;
			data[96605] <= 8'h10 ;
			data[96606] <= 8'h10 ;
			data[96607] <= 8'h10 ;
			data[96608] <= 8'h10 ;
			data[96609] <= 8'h10 ;
			data[96610] <= 8'h10 ;
			data[96611] <= 8'h10 ;
			data[96612] <= 8'h10 ;
			data[96613] <= 8'h10 ;
			data[96614] <= 8'h10 ;
			data[96615] <= 8'h10 ;
			data[96616] <= 8'h10 ;
			data[96617] <= 8'h10 ;
			data[96618] <= 8'h10 ;
			data[96619] <= 8'h10 ;
			data[96620] <= 8'h10 ;
			data[96621] <= 8'h10 ;
			data[96622] <= 8'h10 ;
			data[96623] <= 8'h10 ;
			data[96624] <= 8'h10 ;
			data[96625] <= 8'h10 ;
			data[96626] <= 8'h10 ;
			data[96627] <= 8'h10 ;
			data[96628] <= 8'h10 ;
			data[96629] <= 8'h10 ;
			data[96630] <= 8'h10 ;
			data[96631] <= 8'h10 ;
			data[96632] <= 8'h10 ;
			data[96633] <= 8'h10 ;
			data[96634] <= 8'h10 ;
			data[96635] <= 8'h10 ;
			data[96636] <= 8'h10 ;
			data[96637] <= 8'h10 ;
			data[96638] <= 8'h10 ;
			data[96639] <= 8'h10 ;
			data[96640] <= 8'h10 ;
			data[96641] <= 8'h10 ;
			data[96642] <= 8'h10 ;
			data[96643] <= 8'h10 ;
			data[96644] <= 8'h10 ;
			data[96645] <= 8'h10 ;
			data[96646] <= 8'h10 ;
			data[96647] <= 8'h10 ;
			data[96648] <= 8'h10 ;
			data[96649] <= 8'h10 ;
			data[96650] <= 8'h10 ;
			data[96651] <= 8'h10 ;
			data[96652] <= 8'h10 ;
			data[96653] <= 8'h10 ;
			data[96654] <= 8'h10 ;
			data[96655] <= 8'h10 ;
			data[96656] <= 8'h10 ;
			data[96657] <= 8'h10 ;
			data[96658] <= 8'h10 ;
			data[96659] <= 8'h10 ;
			data[96660] <= 8'h10 ;
			data[96661] <= 8'h10 ;
			data[96662] <= 8'h10 ;
			data[96663] <= 8'h10 ;
			data[96664] <= 8'h10 ;
			data[96665] <= 8'h10 ;
			data[96666] <= 8'h10 ;
			data[96667] <= 8'h10 ;
			data[96668] <= 8'h10 ;
			data[96669] <= 8'h10 ;
			data[96670] <= 8'h10 ;
			data[96671] <= 8'h10 ;
			data[96672] <= 8'h10 ;
			data[96673] <= 8'h10 ;
			data[96674] <= 8'h10 ;
			data[96675] <= 8'h10 ;
			data[96676] <= 8'h10 ;
			data[96677] <= 8'h10 ;
			data[96678] <= 8'h10 ;
			data[96679] <= 8'h10 ;
			data[96680] <= 8'h10 ;
			data[96681] <= 8'h10 ;
			data[96682] <= 8'h10 ;
			data[96683] <= 8'h10 ;
			data[96684] <= 8'h10 ;
			data[96685] <= 8'h10 ;
			data[96686] <= 8'h10 ;
			data[96687] <= 8'h10 ;
			data[96688] <= 8'h10 ;
			data[96689] <= 8'h10 ;
			data[96690] <= 8'h10 ;
			data[96691] <= 8'h10 ;
			data[96692] <= 8'h10 ;
			data[96693] <= 8'h10 ;
			data[96694] <= 8'h10 ;
			data[96695] <= 8'h10 ;
			data[96696] <= 8'h10 ;
			data[96697] <= 8'h10 ;
			data[96698] <= 8'h10 ;
			data[96699] <= 8'h10 ;
			data[96700] <= 8'h10 ;
			data[96701] <= 8'h10 ;
			data[96702] <= 8'h10 ;
			data[96703] <= 8'h10 ;
			data[96704] <= 8'h10 ;
			data[96705] <= 8'h10 ;
			data[96706] <= 8'h10 ;
			data[96707] <= 8'h10 ;
			data[96708] <= 8'h10 ;
			data[96709] <= 8'h10 ;
			data[96710] <= 8'h10 ;
			data[96711] <= 8'h10 ;
			data[96712] <= 8'h10 ;
			data[96713] <= 8'h10 ;
			data[96714] <= 8'h10 ;
			data[96715] <= 8'h10 ;
			data[96716] <= 8'h10 ;
			data[96717] <= 8'h10 ;
			data[96718] <= 8'h10 ;
			data[96719] <= 8'h10 ;
			data[96720] <= 8'h10 ;
			data[96721] <= 8'h10 ;
			data[96722] <= 8'h10 ;
			data[96723] <= 8'h10 ;
			data[96724] <= 8'h10 ;
			data[96725] <= 8'h10 ;
			data[96726] <= 8'h10 ;
			data[96727] <= 8'h10 ;
			data[96728] <= 8'h10 ;
			data[96729] <= 8'h10 ;
			data[96730] <= 8'h10 ;
			data[96731] <= 8'h10 ;
			data[96732] <= 8'h10 ;
			data[96733] <= 8'h10 ;
			data[96734] <= 8'h10 ;
			data[96735] <= 8'h10 ;
			data[96736] <= 8'h10 ;
			data[96737] <= 8'h10 ;
			data[96738] <= 8'h10 ;
			data[96739] <= 8'h10 ;
			data[96740] <= 8'h10 ;
			data[96741] <= 8'h10 ;
			data[96742] <= 8'h10 ;
			data[96743] <= 8'h10 ;
			data[96744] <= 8'h10 ;
			data[96745] <= 8'h10 ;
			data[96746] <= 8'h10 ;
			data[96747] <= 8'h10 ;
			data[96748] <= 8'h10 ;
			data[96749] <= 8'h10 ;
			data[96750] <= 8'h10 ;
			data[96751] <= 8'h10 ;
			data[96752] <= 8'h10 ;
			data[96753] <= 8'h10 ;
			data[96754] <= 8'h10 ;
			data[96755] <= 8'h10 ;
			data[96756] <= 8'h10 ;
			data[96757] <= 8'h10 ;
			data[96758] <= 8'h10 ;
			data[96759] <= 8'h10 ;
			data[96760] <= 8'h10 ;
			data[96761] <= 8'h10 ;
			data[96762] <= 8'h10 ;
			data[96763] <= 8'h10 ;
			data[96764] <= 8'h10 ;
			data[96765] <= 8'h10 ;
			data[96766] <= 8'h10 ;
			data[96767] <= 8'h10 ;
			data[96768] <= 8'h10 ;
			data[96769] <= 8'h10 ;
			data[96770] <= 8'h10 ;
			data[96771] <= 8'h10 ;
			data[96772] <= 8'h10 ;
			data[96773] <= 8'h10 ;
			data[96774] <= 8'h10 ;
			data[96775] <= 8'h10 ;
			data[96776] <= 8'h10 ;
			data[96777] <= 8'h10 ;
			data[96778] <= 8'h10 ;
			data[96779] <= 8'h10 ;
			data[96780] <= 8'h10 ;
			data[96781] <= 8'h10 ;
			data[96782] <= 8'h10 ;
			data[96783] <= 8'h10 ;
			data[96784] <= 8'h10 ;
			data[96785] <= 8'h10 ;
			data[96786] <= 8'h10 ;
			data[96787] <= 8'h10 ;
			data[96788] <= 8'h10 ;
			data[96789] <= 8'h10 ;
			data[96790] <= 8'h10 ;
			data[96791] <= 8'h10 ;
			data[96792] <= 8'h10 ;
			data[96793] <= 8'h10 ;
			data[96794] <= 8'h10 ;
			data[96795] <= 8'h10 ;
			data[96796] <= 8'h10 ;
			data[96797] <= 8'h10 ;
			data[96798] <= 8'h10 ;
			data[96799] <= 8'h10 ;
			data[96800] <= 8'h10 ;
			data[96801] <= 8'h10 ;
			data[96802] <= 8'h10 ;
			data[96803] <= 8'h10 ;
			data[96804] <= 8'h10 ;
			data[96805] <= 8'h10 ;
			data[96806] <= 8'h10 ;
			data[96807] <= 8'h10 ;
			data[96808] <= 8'h10 ;
			data[96809] <= 8'h10 ;
			data[96810] <= 8'h10 ;
			data[96811] <= 8'h10 ;
			data[96812] <= 8'h10 ;
			data[96813] <= 8'h10 ;
			data[96814] <= 8'h10 ;
			data[96815] <= 8'h10 ;
			data[96816] <= 8'h10 ;
			data[96817] <= 8'h10 ;
			data[96818] <= 8'h10 ;
			data[96819] <= 8'h10 ;
			data[96820] <= 8'h10 ;
			data[96821] <= 8'h10 ;
			data[96822] <= 8'h10 ;
			data[96823] <= 8'h10 ;
			data[96824] <= 8'h10 ;
			data[96825] <= 8'h10 ;
			data[96826] <= 8'h10 ;
			data[96827] <= 8'h10 ;
			data[96828] <= 8'h10 ;
			data[96829] <= 8'h10 ;
			data[96830] <= 8'h10 ;
			data[96831] <= 8'h10 ;
			data[96832] <= 8'h10 ;
			data[96833] <= 8'h10 ;
			data[96834] <= 8'h10 ;
			data[96835] <= 8'h10 ;
			data[96836] <= 8'h10 ;
			data[96837] <= 8'h10 ;
			data[96838] <= 8'h10 ;
			data[96839] <= 8'h10 ;
			data[96840] <= 8'h10 ;
			data[96841] <= 8'h10 ;
			data[96842] <= 8'h10 ;
			data[96843] <= 8'h10 ;
			data[96844] <= 8'h10 ;
			data[96845] <= 8'h10 ;
			data[96846] <= 8'h10 ;
			data[96847] <= 8'h10 ;
			data[96848] <= 8'h10 ;
			data[96849] <= 8'h10 ;
			data[96850] <= 8'h10 ;
			data[96851] <= 8'h10 ;
			data[96852] <= 8'h10 ;
			data[96853] <= 8'h10 ;
			data[96854] <= 8'h10 ;
			data[96855] <= 8'h10 ;
			data[96856] <= 8'h10 ;
			data[96857] <= 8'h10 ;
			data[96858] <= 8'h10 ;
			data[96859] <= 8'h10 ;
			data[96860] <= 8'h10 ;
			data[96861] <= 8'h10 ;
			data[96862] <= 8'h10 ;
			data[96863] <= 8'h10 ;
			data[96864] <= 8'h10 ;
			data[96865] <= 8'h10 ;
			data[96866] <= 8'h10 ;
			data[96867] <= 8'h10 ;
			data[96868] <= 8'h10 ;
			data[96869] <= 8'h10 ;
			data[96870] <= 8'h10 ;
			data[96871] <= 8'h10 ;
			data[96872] <= 8'h10 ;
			data[96873] <= 8'h10 ;
			data[96874] <= 8'h10 ;
			data[96875] <= 8'h10 ;
			data[96876] <= 8'h10 ;
			data[96877] <= 8'h10 ;
			data[96878] <= 8'h10 ;
			data[96879] <= 8'h10 ;
			data[96880] <= 8'h10 ;
			data[96881] <= 8'h10 ;
			data[96882] <= 8'h10 ;
			data[96883] <= 8'h10 ;
			data[96884] <= 8'h10 ;
			data[96885] <= 8'h10 ;
			data[96886] <= 8'h10 ;
			data[96887] <= 8'h10 ;
			data[96888] <= 8'h10 ;
			data[96889] <= 8'h10 ;
			data[96890] <= 8'h10 ;
			data[96891] <= 8'h10 ;
			data[96892] <= 8'h10 ;
			data[96893] <= 8'h10 ;
			data[96894] <= 8'h10 ;
			data[96895] <= 8'h10 ;
			data[96896] <= 8'h10 ;
			data[96897] <= 8'h10 ;
			data[96898] <= 8'h10 ;
			data[96899] <= 8'h10 ;
			data[96900] <= 8'h10 ;
			data[96901] <= 8'h10 ;
			data[96902] <= 8'h10 ;
			data[96903] <= 8'h10 ;
			data[96904] <= 8'h10 ;
			data[96905] <= 8'h10 ;
			data[96906] <= 8'h10 ;
			data[96907] <= 8'h10 ;
			data[96908] <= 8'h10 ;
			data[96909] <= 8'h10 ;
			data[96910] <= 8'h10 ;
			data[96911] <= 8'h10 ;
			data[96912] <= 8'h10 ;
			data[96913] <= 8'h10 ;
			data[96914] <= 8'h10 ;
			data[96915] <= 8'h10 ;
			data[96916] <= 8'h10 ;
			data[96917] <= 8'h10 ;
			data[96918] <= 8'h10 ;
			data[96919] <= 8'h10 ;
			data[96920] <= 8'h10 ;
			data[96921] <= 8'h10 ;
			data[96922] <= 8'h10 ;
			data[96923] <= 8'h10 ;
			data[96924] <= 8'h10 ;
			data[96925] <= 8'h10 ;
			data[96926] <= 8'h10 ;
			data[96927] <= 8'h10 ;
			data[96928] <= 8'h10 ;
			data[96929] <= 8'h10 ;
			data[96930] <= 8'h10 ;
			data[96931] <= 8'h10 ;
			data[96932] <= 8'h10 ;
			data[96933] <= 8'h10 ;
			data[96934] <= 8'h10 ;
			data[96935] <= 8'h10 ;
			data[96936] <= 8'h10 ;
			data[96937] <= 8'h10 ;
			data[96938] <= 8'h10 ;
			data[96939] <= 8'h10 ;
			data[96940] <= 8'h10 ;
			data[96941] <= 8'h10 ;
			data[96942] <= 8'h10 ;
			data[96943] <= 8'h10 ;
			data[96944] <= 8'h10 ;
			data[96945] <= 8'h10 ;
			data[96946] <= 8'h10 ;
			data[96947] <= 8'h10 ;
			data[96948] <= 8'h10 ;
			data[96949] <= 8'h10 ;
			data[96950] <= 8'h10 ;
			data[96951] <= 8'h10 ;
			data[96952] <= 8'h10 ;
			data[96953] <= 8'h10 ;
			data[96954] <= 8'h10 ;
			data[96955] <= 8'h10 ;
			data[96956] <= 8'h10 ;
			data[96957] <= 8'h10 ;
			data[96958] <= 8'h10 ;
			data[96959] <= 8'h10 ;
			data[96960] <= 8'h10 ;
			data[96961] <= 8'h10 ;
			data[96962] <= 8'h10 ;
			data[96963] <= 8'h10 ;
			data[96964] <= 8'h10 ;
			data[96965] <= 8'h10 ;
			data[96966] <= 8'h10 ;
			data[96967] <= 8'h10 ;
			data[96968] <= 8'h10 ;
			data[96969] <= 8'h10 ;
			data[96970] <= 8'h10 ;
			data[96971] <= 8'h10 ;
			data[96972] <= 8'h10 ;
			data[96973] <= 8'h10 ;
			data[96974] <= 8'h10 ;
			data[96975] <= 8'h10 ;
			data[96976] <= 8'h10 ;
			data[96977] <= 8'h10 ;
			data[96978] <= 8'h10 ;
			data[96979] <= 8'h10 ;
			data[96980] <= 8'h10 ;
			data[96981] <= 8'h10 ;
			data[96982] <= 8'h10 ;
			data[96983] <= 8'h10 ;
			data[96984] <= 8'h10 ;
			data[96985] <= 8'h10 ;
			data[96986] <= 8'h10 ;
			data[96987] <= 8'h10 ;
			data[96988] <= 8'h10 ;
			data[96989] <= 8'h10 ;
			data[96990] <= 8'h10 ;
			data[96991] <= 8'h10 ;
			data[96992] <= 8'h10 ;
			data[96993] <= 8'h10 ;
			data[96994] <= 8'h10 ;
			data[96995] <= 8'h10 ;
			data[96996] <= 8'h10 ;
			data[96997] <= 8'h10 ;
			data[96998] <= 8'h10 ;
			data[96999] <= 8'h10 ;
			data[97000] <= 8'h10 ;
			data[97001] <= 8'h10 ;
			data[97002] <= 8'h10 ;
			data[97003] <= 8'h10 ;
			data[97004] <= 8'h10 ;
			data[97005] <= 8'h10 ;
			data[97006] <= 8'h10 ;
			data[97007] <= 8'h10 ;
			data[97008] <= 8'h10 ;
			data[97009] <= 8'h10 ;
			data[97010] <= 8'h10 ;
			data[97011] <= 8'h10 ;
			data[97012] <= 8'h10 ;
			data[97013] <= 8'h10 ;
			data[97014] <= 8'h10 ;
			data[97015] <= 8'h10 ;
			data[97016] <= 8'h10 ;
			data[97017] <= 8'h10 ;
			data[97018] <= 8'h10 ;
			data[97019] <= 8'h10 ;
			data[97020] <= 8'h10 ;
			data[97021] <= 8'h10 ;
			data[97022] <= 8'h10 ;
			data[97023] <= 8'h10 ;
			data[97024] <= 8'h10 ;
			data[97025] <= 8'h10 ;
			data[97026] <= 8'h10 ;
			data[97027] <= 8'h10 ;
			data[97028] <= 8'h10 ;
			data[97029] <= 8'h10 ;
			data[97030] <= 8'h10 ;
			data[97031] <= 8'h10 ;
			data[97032] <= 8'h10 ;
			data[97033] <= 8'h10 ;
			data[97034] <= 8'h10 ;
			data[97035] <= 8'h10 ;
			data[97036] <= 8'h10 ;
			data[97037] <= 8'h10 ;
			data[97038] <= 8'h10 ;
			data[97039] <= 8'h10 ;
			data[97040] <= 8'h10 ;
			data[97041] <= 8'h10 ;
			data[97042] <= 8'h10 ;
			data[97043] <= 8'h10 ;
			data[97044] <= 8'h10 ;
			data[97045] <= 8'h10 ;
			data[97046] <= 8'h10 ;
			data[97047] <= 8'h10 ;
			data[97048] <= 8'h10 ;
			data[97049] <= 8'h10 ;
			data[97050] <= 8'h10 ;
			data[97051] <= 8'h10 ;
			data[97052] <= 8'h10 ;
			data[97053] <= 8'h10 ;
			data[97054] <= 8'h10 ;
			data[97055] <= 8'h10 ;
			data[97056] <= 8'h10 ;
			data[97057] <= 8'h10 ;
			data[97058] <= 8'h10 ;
			data[97059] <= 8'h10 ;
			data[97060] <= 8'h10 ;
			data[97061] <= 8'h10 ;
			data[97062] <= 8'h10 ;
			data[97063] <= 8'h10 ;
			data[97064] <= 8'h10 ;
			data[97065] <= 8'h10 ;
			data[97066] <= 8'h10 ;
			data[97067] <= 8'h10 ;
			data[97068] <= 8'h10 ;
			data[97069] <= 8'h10 ;
			data[97070] <= 8'h10 ;
			data[97071] <= 8'h10 ;
			data[97072] <= 8'h10 ;
			data[97073] <= 8'h10 ;
			data[97074] <= 8'h10 ;
			data[97075] <= 8'h10 ;
			data[97076] <= 8'h10 ;
			data[97077] <= 8'h10 ;
			data[97078] <= 8'h10 ;
			data[97079] <= 8'h10 ;
			data[97080] <= 8'h10 ;
			data[97081] <= 8'h10 ;
			data[97082] <= 8'h10 ;
			data[97083] <= 8'h10 ;
			data[97084] <= 8'h10 ;
			data[97085] <= 8'h10 ;
			data[97086] <= 8'h10 ;
			data[97087] <= 8'h10 ;
			data[97088] <= 8'h10 ;
			data[97089] <= 8'h10 ;
			data[97090] <= 8'h10 ;
			data[97091] <= 8'h10 ;
			data[97092] <= 8'h10 ;
			data[97093] <= 8'h10 ;
			data[97094] <= 8'h10 ;
			data[97095] <= 8'h10 ;
			data[97096] <= 8'h10 ;
			data[97097] <= 8'h10 ;
			data[97098] <= 8'h10 ;
			data[97099] <= 8'h10 ;
			data[97100] <= 8'h10 ;
			data[97101] <= 8'h10 ;
			data[97102] <= 8'h10 ;
			data[97103] <= 8'h10 ;
			data[97104] <= 8'h10 ;
			data[97105] <= 8'h10 ;
			data[97106] <= 8'h10 ;
			data[97107] <= 8'h10 ;
			data[97108] <= 8'h10 ;
			data[97109] <= 8'h10 ;
			data[97110] <= 8'h10 ;
			data[97111] <= 8'h10 ;
			data[97112] <= 8'h10 ;
			data[97113] <= 8'h10 ;
			data[97114] <= 8'h10 ;
			data[97115] <= 8'h10 ;
			data[97116] <= 8'h10 ;
			data[97117] <= 8'h10 ;
			data[97118] <= 8'h10 ;
			data[97119] <= 8'h10 ;
			data[97120] <= 8'h10 ;
			data[97121] <= 8'h10 ;
			data[97122] <= 8'h10 ;
			data[97123] <= 8'h10 ;
			data[97124] <= 8'h10 ;
			data[97125] <= 8'h10 ;
			data[97126] <= 8'h10 ;
			data[97127] <= 8'h10 ;
			data[97128] <= 8'h10 ;
			data[97129] <= 8'h10 ;
			data[97130] <= 8'h10 ;
			data[97131] <= 8'h10 ;
			data[97132] <= 8'h10 ;
			data[97133] <= 8'h10 ;
			data[97134] <= 8'h10 ;
			data[97135] <= 8'h10 ;
			data[97136] <= 8'h10 ;
			data[97137] <= 8'h10 ;
			data[97138] <= 8'h10 ;
			data[97139] <= 8'h10 ;
			data[97140] <= 8'h10 ;
			data[97141] <= 8'h10 ;
			data[97142] <= 8'h10 ;
			data[97143] <= 8'h10 ;
			data[97144] <= 8'h10 ;
			data[97145] <= 8'h10 ;
			data[97146] <= 8'h10 ;
			data[97147] <= 8'h10 ;
			data[97148] <= 8'h10 ;
			data[97149] <= 8'h10 ;
			data[97150] <= 8'h10 ;
			data[97151] <= 8'h10 ;
			data[97152] <= 8'h10 ;
			data[97153] <= 8'h10 ;
			data[97154] <= 8'h10 ;
			data[97155] <= 8'h10 ;
			data[97156] <= 8'h10 ;
			data[97157] <= 8'h10 ;
			data[97158] <= 8'h10 ;
			data[97159] <= 8'h10 ;
			data[97160] <= 8'h10 ;
			data[97161] <= 8'h10 ;
			data[97162] <= 8'h10 ;
			data[97163] <= 8'h10 ;
			data[97164] <= 8'h10 ;
			data[97165] <= 8'h10 ;
			data[97166] <= 8'h10 ;
			data[97167] <= 8'h10 ;
			data[97168] <= 8'h10 ;
			data[97169] <= 8'h10 ;
			data[97170] <= 8'h10 ;
			data[97171] <= 8'h10 ;
			data[97172] <= 8'h10 ;
			data[97173] <= 8'h10 ;
			data[97174] <= 8'h10 ;
			data[97175] <= 8'h10 ;
			data[97176] <= 8'h10 ;
			data[97177] <= 8'h10 ;
			data[97178] <= 8'h10 ;
			data[97179] <= 8'h10 ;
			data[97180] <= 8'h10 ;
			data[97181] <= 8'h10 ;
			data[97182] <= 8'h10 ;
			data[97183] <= 8'h10 ;
			data[97184] <= 8'h10 ;
			data[97185] <= 8'h10 ;
			data[97186] <= 8'h10 ;
			data[97187] <= 8'h10 ;
			data[97188] <= 8'h10 ;
			data[97189] <= 8'h10 ;
			data[97190] <= 8'h10 ;
			data[97191] <= 8'h10 ;
			data[97192] <= 8'h10 ;
			data[97193] <= 8'h10 ;
			data[97194] <= 8'h10 ;
			data[97195] <= 8'h10 ;
			data[97196] <= 8'h10 ;
			data[97197] <= 8'h10 ;
			data[97198] <= 8'h10 ;
			data[97199] <= 8'h10 ;
			data[97200] <= 8'h10 ;
			data[97201] <= 8'h10 ;
			data[97202] <= 8'h10 ;
			data[97203] <= 8'h10 ;
			data[97204] <= 8'h10 ;
			data[97205] <= 8'h10 ;
			data[97206] <= 8'h10 ;
			data[97207] <= 8'h10 ;
			data[97208] <= 8'h10 ;
			data[97209] <= 8'h10 ;
			data[97210] <= 8'h10 ;
			data[97211] <= 8'h10 ;
			data[97212] <= 8'h10 ;
			data[97213] <= 8'h10 ;
			data[97214] <= 8'h10 ;
			data[97215] <= 8'h10 ;
			data[97216] <= 8'h10 ;
			data[97217] <= 8'h10 ;
			data[97218] <= 8'h10 ;
			data[97219] <= 8'h10 ;
			data[97220] <= 8'h10 ;
			data[97221] <= 8'h10 ;
			data[97222] <= 8'h10 ;
			data[97223] <= 8'h10 ;
			data[97224] <= 8'h10 ;
			data[97225] <= 8'h10 ;
			data[97226] <= 8'h10 ;
			data[97227] <= 8'h10 ;
			data[97228] <= 8'h10 ;
			data[97229] <= 8'h10 ;
			data[97230] <= 8'h10 ;
			data[97231] <= 8'h10 ;
			data[97232] <= 8'h10 ;
			data[97233] <= 8'h10 ;
			data[97234] <= 8'h10 ;
			data[97235] <= 8'h10 ;
			data[97236] <= 8'h10 ;
			data[97237] <= 8'h10 ;
			data[97238] <= 8'h10 ;
			data[97239] <= 8'h10 ;
			data[97240] <= 8'h10 ;
			data[97241] <= 8'h10 ;
			data[97242] <= 8'h10 ;
			data[97243] <= 8'h10 ;
			data[97244] <= 8'h10 ;
			data[97245] <= 8'h10 ;
			data[97246] <= 8'h10 ;
			data[97247] <= 8'h10 ;
			data[97248] <= 8'h10 ;
			data[97249] <= 8'h10 ;
			data[97250] <= 8'h10 ;
			data[97251] <= 8'h10 ;
			data[97252] <= 8'h10 ;
			data[97253] <= 8'h10 ;
			data[97254] <= 8'h10 ;
			data[97255] <= 8'h10 ;
			data[97256] <= 8'h10 ;
			data[97257] <= 8'h10 ;
			data[97258] <= 8'h10 ;
			data[97259] <= 8'h10 ;
			data[97260] <= 8'h10 ;
			data[97261] <= 8'h10 ;
			data[97262] <= 8'h10 ;
			data[97263] <= 8'h10 ;
			data[97264] <= 8'h10 ;
			data[97265] <= 8'h10 ;
			data[97266] <= 8'h10 ;
			data[97267] <= 8'h10 ;
			data[97268] <= 8'h10 ;
			data[97269] <= 8'h10 ;
			data[97270] <= 8'h10 ;
			data[97271] <= 8'h10 ;
			data[97272] <= 8'h10 ;
			data[97273] <= 8'h10 ;
			data[97274] <= 8'h10 ;
			data[97275] <= 8'h10 ;
			data[97276] <= 8'h10 ;
			data[97277] <= 8'h10 ;
			data[97278] <= 8'h10 ;
			data[97279] <= 8'h10 ;
			data[97280] <= 8'h10 ;
			data[97281] <= 8'h10 ;
			data[97282] <= 8'h10 ;
			data[97283] <= 8'h10 ;
			data[97284] <= 8'h10 ;
			data[97285] <= 8'h10 ;
			data[97286] <= 8'h10 ;
			data[97287] <= 8'h10 ;
			data[97288] <= 8'h10 ;
			data[97289] <= 8'h10 ;
			data[97290] <= 8'h10 ;
			data[97291] <= 8'h10 ;
			data[97292] <= 8'h10 ;
			data[97293] <= 8'h10 ;
			data[97294] <= 8'h10 ;
			data[97295] <= 8'h10 ;
			data[97296] <= 8'h10 ;
			data[97297] <= 8'h10 ;
			data[97298] <= 8'h10 ;
			data[97299] <= 8'h10 ;
			data[97300] <= 8'h10 ;
			data[97301] <= 8'h10 ;
			data[97302] <= 8'h10 ;
			data[97303] <= 8'h10 ;
			data[97304] <= 8'h10 ;
			data[97305] <= 8'h10 ;
			data[97306] <= 8'h10 ;
			data[97307] <= 8'h10 ;
			data[97308] <= 8'h10 ;
			data[97309] <= 8'h10 ;
			data[97310] <= 8'h10 ;
			data[97311] <= 8'h10 ;
			data[97312] <= 8'h10 ;
			data[97313] <= 8'h10 ;
			data[97314] <= 8'h10 ;
			data[97315] <= 8'h10 ;
			data[97316] <= 8'h10 ;
			data[97317] <= 8'h10 ;
			data[97318] <= 8'h10 ;
			data[97319] <= 8'h10 ;
			data[97320] <= 8'h10 ;
			data[97321] <= 8'h10 ;
			data[97322] <= 8'h10 ;
			data[97323] <= 8'h10 ;
			data[97324] <= 8'h10 ;
			data[97325] <= 8'h10 ;
			data[97326] <= 8'h10 ;
			data[97327] <= 8'h10 ;
			data[97328] <= 8'h10 ;
			data[97329] <= 8'h10 ;
			data[97330] <= 8'h10 ;
			data[97331] <= 8'h10 ;
			data[97332] <= 8'h10 ;
			data[97333] <= 8'h10 ;
			data[97334] <= 8'h10 ;
			data[97335] <= 8'h10 ;
			data[97336] <= 8'h10 ;
			data[97337] <= 8'h10 ;
			data[97338] <= 8'h10 ;
			data[97339] <= 8'h10 ;
			data[97340] <= 8'h10 ;
			data[97341] <= 8'h10 ;
			data[97342] <= 8'h10 ;
			data[97343] <= 8'h10 ;
			data[97344] <= 8'h10 ;
			data[97345] <= 8'h10 ;
			data[97346] <= 8'h10 ;
			data[97347] <= 8'h10 ;
			data[97348] <= 8'h10 ;
			data[97349] <= 8'h10 ;
			data[97350] <= 8'h10 ;
			data[97351] <= 8'h10 ;
			data[97352] <= 8'h10 ;
			data[97353] <= 8'h10 ;
			data[97354] <= 8'h10 ;
			data[97355] <= 8'h10 ;
			data[97356] <= 8'h10 ;
			data[97357] <= 8'h10 ;
			data[97358] <= 8'h10 ;
			data[97359] <= 8'h10 ;
			data[97360] <= 8'h10 ;
			data[97361] <= 8'h10 ;
			data[97362] <= 8'h10 ;
			data[97363] <= 8'h10 ;
			data[97364] <= 8'h10 ;
			data[97365] <= 8'h10 ;
			data[97366] <= 8'h10 ;
			data[97367] <= 8'h10 ;
			data[97368] <= 8'h10 ;
			data[97369] <= 8'h10 ;
			data[97370] <= 8'h10 ;
			data[97371] <= 8'h10 ;
			data[97372] <= 8'h10 ;
			data[97373] <= 8'h10 ;
			data[97374] <= 8'h10 ;
			data[97375] <= 8'h10 ;
			data[97376] <= 8'h10 ;
			data[97377] <= 8'h10 ;
			data[97378] <= 8'h10 ;
			data[97379] <= 8'h10 ;
			data[97380] <= 8'h10 ;
			data[97381] <= 8'h10 ;
			data[97382] <= 8'h10 ;
			data[97383] <= 8'h10 ;
			data[97384] <= 8'h10 ;
			data[97385] <= 8'h10 ;
			data[97386] <= 8'h10 ;
			data[97387] <= 8'h10 ;
			data[97388] <= 8'h10 ;
			data[97389] <= 8'h10 ;
			data[97390] <= 8'h10 ;
			data[97391] <= 8'h10 ;
			data[97392] <= 8'h10 ;
			data[97393] <= 8'h10 ;
			data[97394] <= 8'h10 ;
			data[97395] <= 8'h10 ;
			data[97396] <= 8'h10 ;
			data[97397] <= 8'h10 ;
			data[97398] <= 8'h10 ;
			data[97399] <= 8'h10 ;
			data[97400] <= 8'h10 ;
			data[97401] <= 8'h10 ;
			data[97402] <= 8'h10 ;
			data[97403] <= 8'h10 ;
			data[97404] <= 8'h10 ;
			data[97405] <= 8'h10 ;
			data[97406] <= 8'h10 ;
			data[97407] <= 8'h10 ;
			data[97408] <= 8'h10 ;
			data[97409] <= 8'h10 ;
			data[97410] <= 8'h10 ;
			data[97411] <= 8'h10 ;
			data[97412] <= 8'h10 ;
			data[97413] <= 8'h10 ;
			data[97414] <= 8'h10 ;
			data[97415] <= 8'h10 ;
			data[97416] <= 8'h10 ;
			data[97417] <= 8'h10 ;
			data[97418] <= 8'h10 ;
			data[97419] <= 8'h10 ;
			data[97420] <= 8'h10 ;
			data[97421] <= 8'h10 ;
			data[97422] <= 8'h10 ;
			data[97423] <= 8'h10 ;
			data[97424] <= 8'h10 ;
			data[97425] <= 8'h10 ;
			data[97426] <= 8'h10 ;
			data[97427] <= 8'h10 ;
			data[97428] <= 8'h10 ;
			data[97429] <= 8'h10 ;
			data[97430] <= 8'h10 ;
			data[97431] <= 8'h10 ;
			data[97432] <= 8'h10 ;
			data[97433] <= 8'h10 ;
			data[97434] <= 8'h10 ;
			data[97435] <= 8'h10 ;
			data[97436] <= 8'h10 ;
			data[97437] <= 8'h10 ;
			data[97438] <= 8'h10 ;
			data[97439] <= 8'h10 ;
			data[97440] <= 8'h10 ;
			data[97441] <= 8'h10 ;
			data[97442] <= 8'h10 ;
			data[97443] <= 8'h10 ;
			data[97444] <= 8'h10 ;
			data[97445] <= 8'h10 ;
			data[97446] <= 8'h10 ;
			data[97447] <= 8'h10 ;
			data[97448] <= 8'h10 ;
			data[97449] <= 8'h10 ;
			data[97450] <= 8'h10 ;
			data[97451] <= 8'h10 ;
			data[97452] <= 8'h10 ;
			data[97453] <= 8'h10 ;
			data[97454] <= 8'h10 ;
			data[97455] <= 8'h10 ;
			data[97456] <= 8'h10 ;
			data[97457] <= 8'h10 ;
			data[97458] <= 8'h10 ;
			data[97459] <= 8'h10 ;
			data[97460] <= 8'h10 ;
			data[97461] <= 8'h10 ;
			data[97462] <= 8'h10 ;
			data[97463] <= 8'h10 ;
			data[97464] <= 8'h10 ;
			data[97465] <= 8'h10 ;
			data[97466] <= 8'h10 ;
			data[97467] <= 8'h10 ;
			data[97468] <= 8'h10 ;
			data[97469] <= 8'h10 ;
			data[97470] <= 8'h10 ;
			data[97471] <= 8'h10 ;
			data[97472] <= 8'h10 ;
			data[97473] <= 8'h10 ;
			data[97474] <= 8'h10 ;
			data[97475] <= 8'h10 ;
			data[97476] <= 8'h10 ;
			data[97477] <= 8'h10 ;
			data[97478] <= 8'h10 ;
			data[97479] <= 8'h10 ;
			data[97480] <= 8'h10 ;
			data[97481] <= 8'h10 ;
			data[97482] <= 8'h10 ;
			data[97483] <= 8'h10 ;
			data[97484] <= 8'h10 ;
			data[97485] <= 8'h10 ;
			data[97486] <= 8'h10 ;
			data[97487] <= 8'h10 ;
			data[97488] <= 8'h10 ;
			data[97489] <= 8'h10 ;
			data[97490] <= 8'h10 ;
			data[97491] <= 8'h10 ;
			data[97492] <= 8'h10 ;
			data[97493] <= 8'h10 ;
			data[97494] <= 8'h10 ;
			data[97495] <= 8'h10 ;
			data[97496] <= 8'h10 ;
			data[97497] <= 8'h10 ;
			data[97498] <= 8'h10 ;
			data[97499] <= 8'h10 ;
			data[97500] <= 8'h10 ;
			data[97501] <= 8'h10 ;
			data[97502] <= 8'h10 ;
			data[97503] <= 8'h10 ;
			data[97504] <= 8'h10 ;
			data[97505] <= 8'h10 ;
			data[97506] <= 8'h10 ;
			data[97507] <= 8'h10 ;
			data[97508] <= 8'h10 ;
			data[97509] <= 8'h10 ;
			data[97510] <= 8'h10 ;
			data[97511] <= 8'h10 ;
			data[97512] <= 8'h10 ;
			data[97513] <= 8'h10 ;
			data[97514] <= 8'h10 ;
			data[97515] <= 8'h10 ;
			data[97516] <= 8'h10 ;
			data[97517] <= 8'h10 ;
			data[97518] <= 8'h10 ;
			data[97519] <= 8'h10 ;
			data[97520] <= 8'h10 ;
			data[97521] <= 8'h10 ;
			data[97522] <= 8'h10 ;
			data[97523] <= 8'h10 ;
			data[97524] <= 8'h10 ;
			data[97525] <= 8'h10 ;
			data[97526] <= 8'h10 ;
			data[97527] <= 8'h10 ;
			data[97528] <= 8'h10 ;
			data[97529] <= 8'h10 ;
			data[97530] <= 8'h10 ;
			data[97531] <= 8'h10 ;
			data[97532] <= 8'h10 ;
			data[97533] <= 8'h10 ;
			data[97534] <= 8'h10 ;
			data[97535] <= 8'h10 ;
			data[97536] <= 8'h10 ;
			data[97537] <= 8'h10 ;
			data[97538] <= 8'h10 ;
			data[97539] <= 8'h10 ;
			data[97540] <= 8'h10 ;
			data[97541] <= 8'h10 ;
			data[97542] <= 8'h10 ;
			data[97543] <= 8'h10 ;
			data[97544] <= 8'h10 ;
			data[97545] <= 8'h10 ;
			data[97546] <= 8'h10 ;
			data[97547] <= 8'h10 ;
			data[97548] <= 8'h10 ;
			data[97549] <= 8'h10 ;
			data[97550] <= 8'h10 ;
			data[97551] <= 8'h10 ;
			data[97552] <= 8'h10 ;
			data[97553] <= 8'h10 ;
			data[97554] <= 8'h10 ;
			data[97555] <= 8'h10 ;
			data[97556] <= 8'h10 ;
			data[97557] <= 8'h10 ;
			data[97558] <= 8'h10 ;
			data[97559] <= 8'h10 ;
			data[97560] <= 8'h10 ;
			data[97561] <= 8'h10 ;
			data[97562] <= 8'h10 ;
			data[97563] <= 8'h10 ;
			data[97564] <= 8'h10 ;
			data[97565] <= 8'h10 ;
			data[97566] <= 8'h10 ;
			data[97567] <= 8'h10 ;
			data[97568] <= 8'h10 ;
			data[97569] <= 8'h10 ;
			data[97570] <= 8'h10 ;
			data[97571] <= 8'h10 ;
			data[97572] <= 8'h10 ;
			data[97573] <= 8'h10 ;
			data[97574] <= 8'h10 ;
			data[97575] <= 8'h10 ;
			data[97576] <= 8'h10 ;
			data[97577] <= 8'h10 ;
			data[97578] <= 8'h10 ;
			data[97579] <= 8'h10 ;
			data[97580] <= 8'h10 ;
			data[97581] <= 8'h10 ;
			data[97582] <= 8'h10 ;
			data[97583] <= 8'h10 ;
			data[97584] <= 8'h10 ;
			data[97585] <= 8'h10 ;
			data[97586] <= 8'h10 ;
			data[97587] <= 8'h10 ;
			data[97588] <= 8'h10 ;
			data[97589] <= 8'h10 ;
			data[97590] <= 8'h10 ;
			data[97591] <= 8'h10 ;
			data[97592] <= 8'h10 ;
			data[97593] <= 8'h10 ;
			data[97594] <= 8'h10 ;
			data[97595] <= 8'h10 ;
			data[97596] <= 8'h10 ;
			data[97597] <= 8'h10 ;
			data[97598] <= 8'h10 ;
			data[97599] <= 8'h10 ;
			data[97600] <= 8'h10 ;
			data[97601] <= 8'h10 ;
			data[97602] <= 8'h10 ;
			data[97603] <= 8'h10 ;
			data[97604] <= 8'h10 ;
			data[97605] <= 8'h10 ;
			data[97606] <= 8'h10 ;
			data[97607] <= 8'h10 ;
			data[97608] <= 8'h10 ;
			data[97609] <= 8'h10 ;
			data[97610] <= 8'h10 ;
			data[97611] <= 8'h10 ;
			data[97612] <= 8'h10 ;
			data[97613] <= 8'h10 ;
			data[97614] <= 8'h10 ;
			data[97615] <= 8'h10 ;
			data[97616] <= 8'h10 ;
			data[97617] <= 8'h10 ;
			data[97618] <= 8'h10 ;
			data[97619] <= 8'h10 ;
			data[97620] <= 8'h10 ;
			data[97621] <= 8'h10 ;
			data[97622] <= 8'h10 ;
			data[97623] <= 8'h10 ;
			data[97624] <= 8'h10 ;
			data[97625] <= 8'h10 ;
			data[97626] <= 8'h10 ;
			data[97627] <= 8'h10 ;
			data[97628] <= 8'h10 ;
			data[97629] <= 8'h10 ;
			data[97630] <= 8'h10 ;
			data[97631] <= 8'h10 ;
			data[97632] <= 8'h10 ;
			data[97633] <= 8'h10 ;
			data[97634] <= 8'h10 ;
			data[97635] <= 8'h10 ;
			data[97636] <= 8'h10 ;
			data[97637] <= 8'h10 ;
			data[97638] <= 8'h10 ;
			data[97639] <= 8'h10 ;
			data[97640] <= 8'h10 ;
			data[97641] <= 8'h10 ;
			data[97642] <= 8'h10 ;
			data[97643] <= 8'h10 ;
			data[97644] <= 8'h10 ;
			data[97645] <= 8'h10 ;
			data[97646] <= 8'h10 ;
			data[97647] <= 8'h10 ;
			data[97648] <= 8'h10 ;
			data[97649] <= 8'h10 ;
			data[97650] <= 8'h10 ;
			data[97651] <= 8'h10 ;
			data[97652] <= 8'h10 ;
			data[97653] <= 8'h10 ;
			data[97654] <= 8'h10 ;
			data[97655] <= 8'h10 ;
			data[97656] <= 8'h10 ;
			data[97657] <= 8'h10 ;
			data[97658] <= 8'h10 ;
			data[97659] <= 8'h10 ;
			data[97660] <= 8'h10 ;
			data[97661] <= 8'h10 ;
			data[97662] <= 8'h10 ;
			data[97663] <= 8'h10 ;
			data[97664] <= 8'h10 ;
			data[97665] <= 8'h10 ;
			data[97666] <= 8'h10 ;
			data[97667] <= 8'h10 ;
			data[97668] <= 8'h10 ;
			data[97669] <= 8'h10 ;
			data[97670] <= 8'h10 ;
			data[97671] <= 8'h10 ;
			data[97672] <= 8'h10 ;
			data[97673] <= 8'h10 ;
			data[97674] <= 8'h10 ;
			data[97675] <= 8'h10 ;
			data[97676] <= 8'h10 ;
			data[97677] <= 8'h10 ;
			data[97678] <= 8'h10 ;
			data[97679] <= 8'h10 ;
			data[97680] <= 8'h10 ;
			data[97681] <= 8'h10 ;
			data[97682] <= 8'h10 ;
			data[97683] <= 8'h10 ;
			data[97684] <= 8'h10 ;
			data[97685] <= 8'h10 ;
			data[97686] <= 8'h10 ;
			data[97687] <= 8'h10 ;
			data[97688] <= 8'h10 ;
			data[97689] <= 8'h10 ;
			data[97690] <= 8'h10 ;
			data[97691] <= 8'h10 ;
			data[97692] <= 8'h10 ;
			data[97693] <= 8'h10 ;
			data[97694] <= 8'h10 ;
			data[97695] <= 8'h10 ;
			data[97696] <= 8'h10 ;
			data[97697] <= 8'h10 ;
			data[97698] <= 8'h10 ;
			data[97699] <= 8'h10 ;
			data[97700] <= 8'h10 ;
			data[97701] <= 8'h10 ;
			data[97702] <= 8'h10 ;
			data[97703] <= 8'h10 ;
			data[97704] <= 8'h10 ;
			data[97705] <= 8'h10 ;
			data[97706] <= 8'h10 ;
			data[97707] <= 8'h10 ;
			data[97708] <= 8'h10 ;
			data[97709] <= 8'h10 ;
			data[97710] <= 8'h10 ;
			data[97711] <= 8'h10 ;
			data[97712] <= 8'h10 ;
			data[97713] <= 8'h10 ;
			data[97714] <= 8'h10 ;
			data[97715] <= 8'h10 ;
			data[97716] <= 8'h10 ;
			data[97717] <= 8'h10 ;
			data[97718] <= 8'h10 ;
			data[97719] <= 8'h10 ;
			data[97720] <= 8'h10 ;
			data[97721] <= 8'h10 ;
			data[97722] <= 8'h10 ;
			data[97723] <= 8'h10 ;
			data[97724] <= 8'h10 ;
			data[97725] <= 8'h10 ;
			data[97726] <= 8'h10 ;
			data[97727] <= 8'h10 ;
			data[97728] <= 8'h10 ;
			data[97729] <= 8'h10 ;
			data[97730] <= 8'h10 ;
			data[97731] <= 8'h10 ;
			data[97732] <= 8'h10 ;
			data[97733] <= 8'h10 ;
			data[97734] <= 8'h10 ;
			data[97735] <= 8'h10 ;
			data[97736] <= 8'h10 ;
			data[97737] <= 8'h10 ;
			data[97738] <= 8'h10 ;
			data[97739] <= 8'h10 ;
			data[97740] <= 8'h10 ;
			data[97741] <= 8'h10 ;
			data[97742] <= 8'h10 ;
			data[97743] <= 8'h10 ;
			data[97744] <= 8'h10 ;
			data[97745] <= 8'h10 ;
			data[97746] <= 8'h10 ;
			data[97747] <= 8'h10 ;
			data[97748] <= 8'h10 ;
			data[97749] <= 8'h10 ;
			data[97750] <= 8'h10 ;
			data[97751] <= 8'h10 ;
			data[97752] <= 8'h10 ;
			data[97753] <= 8'h10 ;
			data[97754] <= 8'h10 ;
			data[97755] <= 8'h10 ;
			data[97756] <= 8'h10 ;
			data[97757] <= 8'h10 ;
			data[97758] <= 8'h10 ;
			data[97759] <= 8'h10 ;
			data[97760] <= 8'h10 ;
			data[97761] <= 8'h10 ;
			data[97762] <= 8'h10 ;
			data[97763] <= 8'h10 ;
			data[97764] <= 8'h10 ;
			data[97765] <= 8'h10 ;
			data[97766] <= 8'h10 ;
			data[97767] <= 8'h10 ;
			data[97768] <= 8'h10 ;
			data[97769] <= 8'h10 ;
			data[97770] <= 8'h10 ;
			data[97771] <= 8'h10 ;
			data[97772] <= 8'h10 ;
			data[97773] <= 8'h10 ;
			data[97774] <= 8'h10 ;
			data[97775] <= 8'h10 ;
			data[97776] <= 8'h10 ;
			data[97777] <= 8'h10 ;
			data[97778] <= 8'h10 ;
			data[97779] <= 8'h10 ;
			data[97780] <= 8'h10 ;
			data[97781] <= 8'h10 ;
			data[97782] <= 8'h10 ;
			data[97783] <= 8'h10 ;
			data[97784] <= 8'h10 ;
			data[97785] <= 8'h10 ;
			data[97786] <= 8'h10 ;
			data[97787] <= 8'h10 ;
			data[97788] <= 8'h10 ;
			data[97789] <= 8'h10 ;
			data[97790] <= 8'h10 ;
			data[97791] <= 8'h10 ;
			data[97792] <= 8'h10 ;
			data[97793] <= 8'h10 ;
			data[97794] <= 8'h10 ;
			data[97795] <= 8'h10 ;
			data[97796] <= 8'h10 ;
			data[97797] <= 8'h10 ;
			data[97798] <= 8'h10 ;
			data[97799] <= 8'h10 ;
			data[97800] <= 8'h10 ;
			data[97801] <= 8'h10 ;
			data[97802] <= 8'h10 ;
			data[97803] <= 8'h10 ;
			data[97804] <= 8'h10 ;
			data[97805] <= 8'h10 ;
			data[97806] <= 8'h10 ;
			data[97807] <= 8'h10 ;
			data[97808] <= 8'h10 ;
			data[97809] <= 8'h10 ;
			data[97810] <= 8'h10 ;
			data[97811] <= 8'h10 ;
			data[97812] <= 8'h10 ;
			data[97813] <= 8'h10 ;
			data[97814] <= 8'h10 ;
			data[97815] <= 8'h10 ;
			data[97816] <= 8'h10 ;
			data[97817] <= 8'h10 ;
			data[97818] <= 8'h10 ;
			data[97819] <= 8'h10 ;
			data[97820] <= 8'h10 ;
			data[97821] <= 8'h10 ;
			data[97822] <= 8'h10 ;
			data[97823] <= 8'h10 ;
			data[97824] <= 8'h10 ;
			data[97825] <= 8'h10 ;
			data[97826] <= 8'h10 ;
			data[97827] <= 8'h10 ;
			data[97828] <= 8'h10 ;
			data[97829] <= 8'h10 ;
			data[97830] <= 8'h10 ;
			data[97831] <= 8'h10 ;
			data[97832] <= 8'h10 ;
			data[97833] <= 8'h10 ;
			data[97834] <= 8'h10 ;
			data[97835] <= 8'h10 ;
			data[97836] <= 8'h10 ;
			data[97837] <= 8'h10 ;
			data[97838] <= 8'h10 ;
			data[97839] <= 8'h10 ;
			data[97840] <= 8'h10 ;
			data[97841] <= 8'h10 ;
			data[97842] <= 8'h10 ;
			data[97843] <= 8'h10 ;
			data[97844] <= 8'h10 ;
			data[97845] <= 8'h10 ;
			data[97846] <= 8'h10 ;
			data[97847] <= 8'h10 ;
			data[97848] <= 8'h10 ;
			data[97849] <= 8'h10 ;
			data[97850] <= 8'h10 ;
			data[97851] <= 8'h10 ;
			data[97852] <= 8'h10 ;
			data[97853] <= 8'h10 ;
			data[97854] <= 8'h10 ;
			data[97855] <= 8'h10 ;
			data[97856] <= 8'h10 ;
			data[97857] <= 8'h10 ;
			data[97858] <= 8'h10 ;
			data[97859] <= 8'h10 ;
			data[97860] <= 8'h10 ;
			data[97861] <= 8'h10 ;
			data[97862] <= 8'h10 ;
			data[97863] <= 8'h10 ;
			data[97864] <= 8'h10 ;
			data[97865] <= 8'h10 ;
			data[97866] <= 8'h10 ;
			data[97867] <= 8'h10 ;
			data[97868] <= 8'h10 ;
			data[97869] <= 8'h10 ;
			data[97870] <= 8'h10 ;
			data[97871] <= 8'h10 ;
			data[97872] <= 8'h10 ;
			data[97873] <= 8'h10 ;
			data[97874] <= 8'h10 ;
			data[97875] <= 8'h10 ;
			data[97876] <= 8'h10 ;
			data[97877] <= 8'h10 ;
			data[97878] <= 8'h10 ;
			data[97879] <= 8'h10 ;
			data[97880] <= 8'h10 ;
			data[97881] <= 8'h10 ;
			data[97882] <= 8'h10 ;
			data[97883] <= 8'h10 ;
			data[97884] <= 8'h10 ;
			data[97885] <= 8'h10 ;
			data[97886] <= 8'h10 ;
			data[97887] <= 8'h10 ;
			data[97888] <= 8'h10 ;
			data[97889] <= 8'h10 ;
			data[97890] <= 8'h10 ;
			data[97891] <= 8'h10 ;
			data[97892] <= 8'h10 ;
			data[97893] <= 8'h10 ;
			data[97894] <= 8'h10 ;
			data[97895] <= 8'h10 ;
			data[97896] <= 8'h10 ;
			data[97897] <= 8'h10 ;
			data[97898] <= 8'h10 ;
			data[97899] <= 8'h10 ;
			data[97900] <= 8'h10 ;
			data[97901] <= 8'h10 ;
			data[97902] <= 8'h10 ;
			data[97903] <= 8'h10 ;
			data[97904] <= 8'h10 ;
			data[97905] <= 8'h10 ;
			data[97906] <= 8'h10 ;
			data[97907] <= 8'h10 ;
			data[97908] <= 8'h10 ;
			data[97909] <= 8'h10 ;
			data[97910] <= 8'h10 ;
			data[97911] <= 8'h10 ;
			data[97912] <= 8'h10 ;
			data[97913] <= 8'h10 ;
			data[97914] <= 8'h10 ;
			data[97915] <= 8'h10 ;
			data[97916] <= 8'h10 ;
			data[97917] <= 8'h10 ;
			data[97918] <= 8'h10 ;
			data[97919] <= 8'h10 ;
			data[97920] <= 8'h10 ;
			data[97921] <= 8'h10 ;
			data[97922] <= 8'h10 ;
			data[97923] <= 8'h10 ;
			data[97924] <= 8'h10 ;
			data[97925] <= 8'h10 ;
			data[97926] <= 8'h10 ;
			data[97927] <= 8'h10 ;
			data[97928] <= 8'h10 ;
			data[97929] <= 8'h10 ;
			data[97930] <= 8'h10 ;
			data[97931] <= 8'h10 ;
			data[97932] <= 8'h10 ;
			data[97933] <= 8'h10 ;
			data[97934] <= 8'h10 ;
			data[97935] <= 8'h10 ;
			data[97936] <= 8'h10 ;
			data[97937] <= 8'h10 ;
			data[97938] <= 8'h10 ;
			data[97939] <= 8'h10 ;
			data[97940] <= 8'h10 ;
			data[97941] <= 8'h10 ;
			data[97942] <= 8'h10 ;
			data[97943] <= 8'h10 ;
			data[97944] <= 8'h10 ;
			data[97945] <= 8'h10 ;
			data[97946] <= 8'h10 ;
			data[97947] <= 8'h10 ;
			data[97948] <= 8'h10 ;
			data[97949] <= 8'h10 ;
			data[97950] <= 8'h10 ;
			data[97951] <= 8'h10 ;
			data[97952] <= 8'h10 ;
			data[97953] <= 8'h10 ;
			data[97954] <= 8'h10 ;
			data[97955] <= 8'h10 ;
			data[97956] <= 8'h10 ;
			data[97957] <= 8'h10 ;
			data[97958] <= 8'h10 ;
			data[97959] <= 8'h10 ;
			data[97960] <= 8'h10 ;
			data[97961] <= 8'h10 ;
			data[97962] <= 8'h10 ;
			data[97963] <= 8'h10 ;
			data[97964] <= 8'h10 ;
			data[97965] <= 8'h10 ;
			data[97966] <= 8'h10 ;
			data[97967] <= 8'h10 ;
			data[97968] <= 8'h10 ;
			data[97969] <= 8'h10 ;
			data[97970] <= 8'h10 ;
			data[97971] <= 8'h10 ;
			data[97972] <= 8'h10 ;
			data[97973] <= 8'h10 ;
			data[97974] <= 8'h10 ;
			data[97975] <= 8'h10 ;
			data[97976] <= 8'h10 ;
			data[97977] <= 8'h10 ;
			data[97978] <= 8'h10 ;
			data[97979] <= 8'h10 ;
			data[97980] <= 8'h10 ;
			data[97981] <= 8'h10 ;
			data[97982] <= 8'h10 ;
			data[97983] <= 8'h10 ;
			data[97984] <= 8'h10 ;
			data[97985] <= 8'h10 ;
			data[97986] <= 8'h10 ;
			data[97987] <= 8'h10 ;
			data[97988] <= 8'h10 ;
			data[97989] <= 8'h10 ;
			data[97990] <= 8'h10 ;
			data[97991] <= 8'h10 ;
			data[97992] <= 8'h10 ;
			data[97993] <= 8'h10 ;
			data[97994] <= 8'h10 ;
			data[97995] <= 8'h10 ;
			data[97996] <= 8'h10 ;
			data[97997] <= 8'h10 ;
			data[97998] <= 8'h10 ;
			data[97999] <= 8'h10 ;
			data[98000] <= 8'h10 ;
			data[98001] <= 8'h10 ;
			data[98002] <= 8'h10 ;
			data[98003] <= 8'h10 ;
			data[98004] <= 8'h10 ;
			data[98005] <= 8'h10 ;
			data[98006] <= 8'h10 ;
			data[98007] <= 8'h10 ;
			data[98008] <= 8'h10 ;
			data[98009] <= 8'h10 ;
			data[98010] <= 8'h10 ;
			data[98011] <= 8'h10 ;
			data[98012] <= 8'h10 ;
			data[98013] <= 8'h10 ;
			data[98014] <= 8'h10 ;
			data[98015] <= 8'h10 ;
			data[98016] <= 8'h10 ;
			data[98017] <= 8'h10 ;
			data[98018] <= 8'h10 ;
			data[98019] <= 8'h10 ;
			data[98020] <= 8'h10 ;
			data[98021] <= 8'h10 ;
			data[98022] <= 8'h10 ;
			data[98023] <= 8'h10 ;
			data[98024] <= 8'h10 ;
			data[98025] <= 8'h10 ;
			data[98026] <= 8'h10 ;
			data[98027] <= 8'h10 ;
			data[98028] <= 8'h10 ;
			data[98029] <= 8'h10 ;
			data[98030] <= 8'h10 ;
			data[98031] <= 8'h10 ;
			data[98032] <= 8'h10 ;
			data[98033] <= 8'h10 ;
			data[98034] <= 8'h10 ;
			data[98035] <= 8'h10 ;
			data[98036] <= 8'h10 ;
			data[98037] <= 8'h10 ;
			data[98038] <= 8'h10 ;
			data[98039] <= 8'h10 ;
			data[98040] <= 8'h10 ;
			data[98041] <= 8'h10 ;
			data[98042] <= 8'h10 ;
			data[98043] <= 8'h10 ;
			data[98044] <= 8'h10 ;
			data[98045] <= 8'h10 ;
			data[98046] <= 8'h10 ;
			data[98047] <= 8'h10 ;
			data[98048] <= 8'h10 ;
			data[98049] <= 8'h10 ;
			data[98050] <= 8'h10 ;
			data[98051] <= 8'h10 ;
			data[98052] <= 8'h10 ;
			data[98053] <= 8'h10 ;
			data[98054] <= 8'h10 ;
			data[98055] <= 8'h10 ;
			data[98056] <= 8'h10 ;
			data[98057] <= 8'h10 ;
			data[98058] <= 8'h10 ;
			data[98059] <= 8'h10 ;
			data[98060] <= 8'h10 ;
			data[98061] <= 8'h10 ;
			data[98062] <= 8'h10 ;
			data[98063] <= 8'h10 ;
			data[98064] <= 8'h10 ;
			data[98065] <= 8'h10 ;
			data[98066] <= 8'h10 ;
			data[98067] <= 8'h10 ;
			data[98068] <= 8'h10 ;
			data[98069] <= 8'h10 ;
			data[98070] <= 8'h10 ;
			data[98071] <= 8'h10 ;
			data[98072] <= 8'h10 ;
			data[98073] <= 8'h10 ;
			data[98074] <= 8'h10 ;
			data[98075] <= 8'h10 ;
			data[98076] <= 8'h10 ;
			data[98077] <= 8'h10 ;
			data[98078] <= 8'h10 ;
			data[98079] <= 8'h10 ;
			data[98080] <= 8'h10 ;
			data[98081] <= 8'h10 ;
			data[98082] <= 8'h10 ;
			data[98083] <= 8'h10 ;
			data[98084] <= 8'h10 ;
			data[98085] <= 8'h10 ;
			data[98086] <= 8'h10 ;
			data[98087] <= 8'h10 ;
			data[98088] <= 8'h10 ;
			data[98089] <= 8'h10 ;
			data[98090] <= 8'h10 ;
			data[98091] <= 8'h10 ;
			data[98092] <= 8'h10 ;
			data[98093] <= 8'h10 ;
			data[98094] <= 8'h10 ;
			data[98095] <= 8'h10 ;
			data[98096] <= 8'h10 ;
			data[98097] <= 8'h10 ;
			data[98098] <= 8'h10 ;
			data[98099] <= 8'h10 ;
			data[98100] <= 8'h10 ;
			data[98101] <= 8'h10 ;
			data[98102] <= 8'h10 ;
			data[98103] <= 8'h10 ;
			data[98104] <= 8'h10 ;
			data[98105] <= 8'h10 ;
			data[98106] <= 8'h10 ;
			data[98107] <= 8'h10 ;
			data[98108] <= 8'h10 ;
			data[98109] <= 8'h10 ;
			data[98110] <= 8'h10 ;
			data[98111] <= 8'h10 ;
			data[98112] <= 8'h10 ;
			data[98113] <= 8'h10 ;
			data[98114] <= 8'h10 ;
			data[98115] <= 8'h10 ;
			data[98116] <= 8'h10 ;
			data[98117] <= 8'h10 ;
			data[98118] <= 8'h10 ;
			data[98119] <= 8'h10 ;
			data[98120] <= 8'h10 ;
			data[98121] <= 8'h10 ;
			data[98122] <= 8'h10 ;
			data[98123] <= 8'h10 ;
			data[98124] <= 8'h10 ;
			data[98125] <= 8'h10 ;
			data[98126] <= 8'h10 ;
			data[98127] <= 8'h10 ;
			data[98128] <= 8'h10 ;
			data[98129] <= 8'h10 ;
			data[98130] <= 8'h10 ;
			data[98131] <= 8'h10 ;
			data[98132] <= 8'h10 ;
			data[98133] <= 8'h10 ;
			data[98134] <= 8'h10 ;
			data[98135] <= 8'h10 ;
			data[98136] <= 8'h10 ;
			data[98137] <= 8'h10 ;
			data[98138] <= 8'h10 ;
			data[98139] <= 8'h10 ;
			data[98140] <= 8'h10 ;
			data[98141] <= 8'h10 ;
			data[98142] <= 8'h10 ;
			data[98143] <= 8'h10 ;
			data[98144] <= 8'h10 ;
			data[98145] <= 8'h10 ;
			data[98146] <= 8'h10 ;
			data[98147] <= 8'h10 ;
			data[98148] <= 8'h10 ;
			data[98149] <= 8'h10 ;
			data[98150] <= 8'h10 ;
			data[98151] <= 8'h10 ;
			data[98152] <= 8'h10 ;
			data[98153] <= 8'h10 ;
			data[98154] <= 8'h10 ;
			data[98155] <= 8'h10 ;
			data[98156] <= 8'h10 ;
			data[98157] <= 8'h10 ;
			data[98158] <= 8'h10 ;
			data[98159] <= 8'h10 ;
			data[98160] <= 8'h10 ;
			data[98161] <= 8'h10 ;
			data[98162] <= 8'h10 ;
			data[98163] <= 8'h10 ;
			data[98164] <= 8'h10 ;
			data[98165] <= 8'h10 ;
			data[98166] <= 8'h10 ;
			data[98167] <= 8'h10 ;
			data[98168] <= 8'h10 ;
			data[98169] <= 8'h10 ;
			data[98170] <= 8'h10 ;
			data[98171] <= 8'h10 ;
			data[98172] <= 8'h10 ;
			data[98173] <= 8'h10 ;
			data[98174] <= 8'h10 ;
			data[98175] <= 8'h10 ;
			data[98176] <= 8'h10 ;
			data[98177] <= 8'h10 ;
			data[98178] <= 8'h10 ;
			data[98179] <= 8'h10 ;
			data[98180] <= 8'h10 ;
			data[98181] <= 8'h10 ;
			data[98182] <= 8'h10 ;
			data[98183] <= 8'h10 ;
			data[98184] <= 8'h10 ;
			data[98185] <= 8'h10 ;
			data[98186] <= 8'h10 ;
			data[98187] <= 8'h10 ;
			data[98188] <= 8'h10 ;
			data[98189] <= 8'h10 ;
			data[98190] <= 8'h10 ;
			data[98191] <= 8'h10 ;
			data[98192] <= 8'h10 ;
			data[98193] <= 8'h10 ;
			data[98194] <= 8'h10 ;
			data[98195] <= 8'h10 ;
			data[98196] <= 8'h10 ;
			data[98197] <= 8'h10 ;
			data[98198] <= 8'h10 ;
			data[98199] <= 8'h10 ;
			data[98200] <= 8'h10 ;
			data[98201] <= 8'h10 ;
			data[98202] <= 8'h10 ;
			data[98203] <= 8'h10 ;
			data[98204] <= 8'h10 ;
			data[98205] <= 8'h10 ;
			data[98206] <= 8'h10 ;
			data[98207] <= 8'h10 ;
			data[98208] <= 8'h10 ;
			data[98209] <= 8'h10 ;
			data[98210] <= 8'h10 ;
			data[98211] <= 8'h10 ;
			data[98212] <= 8'h10 ;
			data[98213] <= 8'h10 ;
			data[98214] <= 8'h10 ;
			data[98215] <= 8'h10 ;
			data[98216] <= 8'h10 ;
			data[98217] <= 8'h10 ;
			data[98218] <= 8'h10 ;
			data[98219] <= 8'h10 ;
			data[98220] <= 8'h10 ;
			data[98221] <= 8'h10 ;
			data[98222] <= 8'h10 ;
			data[98223] <= 8'h10 ;
			data[98224] <= 8'h10 ;
			data[98225] <= 8'h10 ;
			data[98226] <= 8'h10 ;
			data[98227] <= 8'h10 ;
			data[98228] <= 8'h10 ;
			data[98229] <= 8'h10 ;
			data[98230] <= 8'h10 ;
			data[98231] <= 8'h10 ;
			data[98232] <= 8'h10 ;
			data[98233] <= 8'h10 ;
			data[98234] <= 8'h10 ;
			data[98235] <= 8'h10 ;
			data[98236] <= 8'h10 ;
			data[98237] <= 8'h10 ;
			data[98238] <= 8'h10 ;
			data[98239] <= 8'h10 ;
			data[98240] <= 8'h10 ;
			data[98241] <= 8'h10 ;
			data[98242] <= 8'h10 ;
			data[98243] <= 8'h10 ;
			data[98244] <= 8'h10 ;
			data[98245] <= 8'h10 ;
			data[98246] <= 8'h10 ;
			data[98247] <= 8'h10 ;
			data[98248] <= 8'h10 ;
			data[98249] <= 8'h10 ;
			data[98250] <= 8'h10 ;
			data[98251] <= 8'h10 ;
			data[98252] <= 8'h10 ;
			data[98253] <= 8'h10 ;
			data[98254] <= 8'h10 ;
			data[98255] <= 8'h10 ;
			data[98256] <= 8'h10 ;
			data[98257] <= 8'h10 ;
			data[98258] <= 8'h10 ;
			data[98259] <= 8'h10 ;
			data[98260] <= 8'h10 ;
			data[98261] <= 8'h10 ;
			data[98262] <= 8'h10 ;
			data[98263] <= 8'h10 ;
			data[98264] <= 8'h10 ;
			data[98265] <= 8'h10 ;
			data[98266] <= 8'h10 ;
			data[98267] <= 8'h10 ;
			data[98268] <= 8'h10 ;
			data[98269] <= 8'h10 ;
			data[98270] <= 8'h10 ;
			data[98271] <= 8'h10 ;
			data[98272] <= 8'h10 ;
			data[98273] <= 8'h10 ;
			data[98274] <= 8'h10 ;
			data[98275] <= 8'h10 ;
			data[98276] <= 8'h10 ;
			data[98277] <= 8'h10 ;
			data[98278] <= 8'h10 ;
			data[98279] <= 8'h10 ;
			data[98280] <= 8'h10 ;
			data[98281] <= 8'h10 ;
			data[98282] <= 8'h10 ;
			data[98283] <= 8'h10 ;
			data[98284] <= 8'h10 ;
			data[98285] <= 8'h10 ;
			data[98286] <= 8'h10 ;
			data[98287] <= 8'h10 ;
			data[98288] <= 8'h10 ;
			data[98289] <= 8'h10 ;
			data[98290] <= 8'h10 ;
			data[98291] <= 8'h10 ;
			data[98292] <= 8'h10 ;
			data[98293] <= 8'h10 ;
			data[98294] <= 8'h10 ;
			data[98295] <= 8'h10 ;
			data[98296] <= 8'h10 ;
			data[98297] <= 8'h10 ;
			data[98298] <= 8'h10 ;
			data[98299] <= 8'h10 ;
			data[98300] <= 8'h10 ;
			data[98301] <= 8'h10 ;
			data[98302] <= 8'h10 ;
			data[98303] <= 8'h10 ;
			data[98304] <= 8'h10 ;
			data[98305] <= 8'h10 ;
			data[98306] <= 8'h10 ;
			data[98307] <= 8'h10 ;
			data[98308] <= 8'h10 ;
			data[98309] <= 8'h10 ;
			data[98310] <= 8'h10 ;
			data[98311] <= 8'h10 ;
			data[98312] <= 8'h10 ;
			data[98313] <= 8'h10 ;
			data[98314] <= 8'h10 ;
			data[98315] <= 8'h10 ;
			data[98316] <= 8'h10 ;
			data[98317] <= 8'h10 ;
			data[98318] <= 8'h10 ;
			data[98319] <= 8'h10 ;
			data[98320] <= 8'h10 ;
			data[98321] <= 8'h10 ;
			data[98322] <= 8'h10 ;
			data[98323] <= 8'h10 ;
			data[98324] <= 8'h10 ;
			data[98325] <= 8'h10 ;
			data[98326] <= 8'h10 ;
			data[98327] <= 8'h10 ;
			data[98328] <= 8'h10 ;
			data[98329] <= 8'h10 ;
			data[98330] <= 8'h10 ;
			data[98331] <= 8'h10 ;
			data[98332] <= 8'h10 ;
			data[98333] <= 8'h10 ;
			data[98334] <= 8'h10 ;
			data[98335] <= 8'h10 ;
			data[98336] <= 8'h10 ;
			data[98337] <= 8'h10 ;
			data[98338] <= 8'h10 ;
			data[98339] <= 8'h10 ;
			data[98340] <= 8'h10 ;
			data[98341] <= 8'h10 ;
			data[98342] <= 8'h10 ;
			data[98343] <= 8'h10 ;
			data[98344] <= 8'h10 ;
			data[98345] <= 8'h10 ;
			data[98346] <= 8'h10 ;
			data[98347] <= 8'h10 ;
			data[98348] <= 8'h10 ;
			data[98349] <= 8'h10 ;
			data[98350] <= 8'h10 ;
			data[98351] <= 8'h10 ;
			data[98352] <= 8'h10 ;
			data[98353] <= 8'h10 ;
			data[98354] <= 8'h10 ;
			data[98355] <= 8'h10 ;
			data[98356] <= 8'h10 ;
			data[98357] <= 8'h10 ;
			data[98358] <= 8'h10 ;
			data[98359] <= 8'h10 ;
			data[98360] <= 8'h10 ;
			data[98361] <= 8'h10 ;
			data[98362] <= 8'h10 ;
			data[98363] <= 8'h10 ;
			data[98364] <= 8'h10 ;
			data[98365] <= 8'h10 ;
			data[98366] <= 8'h10 ;
			data[98367] <= 8'h10 ;
			data[98368] <= 8'h10 ;
			data[98369] <= 8'h10 ;
			data[98370] <= 8'h10 ;
			data[98371] <= 8'h10 ;
			data[98372] <= 8'h10 ;
			data[98373] <= 8'h10 ;
			data[98374] <= 8'h10 ;
			data[98375] <= 8'h10 ;
			data[98376] <= 8'h10 ;
			data[98377] <= 8'h10 ;
			data[98378] <= 8'h10 ;
			data[98379] <= 8'h10 ;
			data[98380] <= 8'h10 ;
			data[98381] <= 8'h10 ;
			data[98382] <= 8'h10 ;
			data[98383] <= 8'h10 ;
			data[98384] <= 8'h10 ;
			data[98385] <= 8'h10 ;
			data[98386] <= 8'h10 ;
			data[98387] <= 8'h10 ;
			data[98388] <= 8'h10 ;
			data[98389] <= 8'h10 ;
			data[98390] <= 8'h10 ;
			data[98391] <= 8'h10 ;
			data[98392] <= 8'h10 ;
			data[98393] <= 8'h10 ;
			data[98394] <= 8'h10 ;
			data[98395] <= 8'h10 ;
			data[98396] <= 8'h10 ;
			data[98397] <= 8'h10 ;
			data[98398] <= 8'h10 ;
			data[98399] <= 8'h10 ;
			data[98400] <= 8'h10 ;
			data[98401] <= 8'h10 ;
			data[98402] <= 8'h10 ;
			data[98403] <= 8'h10 ;
			data[98404] <= 8'h10 ;
			data[98405] <= 8'h10 ;
			data[98406] <= 8'h10 ;
			data[98407] <= 8'h10 ;
			data[98408] <= 8'h10 ;
			data[98409] <= 8'h10 ;
			data[98410] <= 8'h10 ;
			data[98411] <= 8'h10 ;
			data[98412] <= 8'h10 ;
			data[98413] <= 8'h10 ;
			data[98414] <= 8'h10 ;
			data[98415] <= 8'h10 ;
			data[98416] <= 8'h10 ;
			data[98417] <= 8'h10 ;
			data[98418] <= 8'h10 ;
			data[98419] <= 8'h10 ;
			data[98420] <= 8'h10 ;
			data[98421] <= 8'h10 ;
			data[98422] <= 8'h10 ;
			data[98423] <= 8'h10 ;
			data[98424] <= 8'h10 ;
			data[98425] <= 8'h10 ;
			data[98426] <= 8'h10 ;
			data[98427] <= 8'h10 ;
			data[98428] <= 8'h10 ;
			data[98429] <= 8'h10 ;
			data[98430] <= 8'h10 ;
			data[98431] <= 8'h10 ;
			data[98432] <= 8'h10 ;
			data[98433] <= 8'h10 ;
			data[98434] <= 8'h10 ;
			data[98435] <= 8'h10 ;
			data[98436] <= 8'h10 ;
			data[98437] <= 8'h10 ;
			data[98438] <= 8'h10 ;
			data[98439] <= 8'h10 ;
			data[98440] <= 8'h10 ;
			data[98441] <= 8'h10 ;
			data[98442] <= 8'h10 ;
			data[98443] <= 8'h10 ;
			data[98444] <= 8'h10 ;
			data[98445] <= 8'h10 ;
			data[98446] <= 8'h10 ;
			data[98447] <= 8'h10 ;
			data[98448] <= 8'h10 ;
			data[98449] <= 8'h10 ;
			data[98450] <= 8'h10 ;
			data[98451] <= 8'h10 ;
			data[98452] <= 8'h10 ;
			data[98453] <= 8'h10 ;
			data[98454] <= 8'h10 ;
			data[98455] <= 8'h10 ;
			data[98456] <= 8'h10 ;
			data[98457] <= 8'h10 ;
			data[98458] <= 8'h10 ;
			data[98459] <= 8'h10 ;
			data[98460] <= 8'h10 ;
			data[98461] <= 8'h10 ;
			data[98462] <= 8'h10 ;
			data[98463] <= 8'h10 ;
			data[98464] <= 8'h10 ;
			data[98465] <= 8'h10 ;
			data[98466] <= 8'h10 ;
			data[98467] <= 8'h10 ;
			data[98468] <= 8'h10 ;
			data[98469] <= 8'h10 ;
			data[98470] <= 8'h10 ;
			data[98471] <= 8'h10 ;
			data[98472] <= 8'h10 ;
			data[98473] <= 8'h10 ;
			data[98474] <= 8'h10 ;
			data[98475] <= 8'h10 ;
			data[98476] <= 8'h10 ;
			data[98477] <= 8'h10 ;
			data[98478] <= 8'h10 ;
			data[98479] <= 8'h10 ;
			data[98480] <= 8'h10 ;
			data[98481] <= 8'h10 ;
			data[98482] <= 8'h10 ;
			data[98483] <= 8'h10 ;
			data[98484] <= 8'h10 ;
			data[98485] <= 8'h10 ;
			data[98486] <= 8'h10 ;
			data[98487] <= 8'h10 ;
			data[98488] <= 8'h10 ;
			data[98489] <= 8'h10 ;
			data[98490] <= 8'h10 ;
			data[98491] <= 8'h10 ;
			data[98492] <= 8'h10 ;
			data[98493] <= 8'h10 ;
			data[98494] <= 8'h10 ;
			data[98495] <= 8'h10 ;
			data[98496] <= 8'h10 ;
			data[98497] <= 8'h10 ;
			data[98498] <= 8'h10 ;
			data[98499] <= 8'h10 ;
			data[98500] <= 8'h10 ;
			data[98501] <= 8'h10 ;
			data[98502] <= 8'h10 ;
			data[98503] <= 8'h10 ;
			data[98504] <= 8'h10 ;
			data[98505] <= 8'h10 ;
			data[98506] <= 8'h10 ;
			data[98507] <= 8'h10 ;
			data[98508] <= 8'h10 ;
			data[98509] <= 8'h10 ;
			data[98510] <= 8'h10 ;
			data[98511] <= 8'h10 ;
			data[98512] <= 8'h10 ;
			data[98513] <= 8'h10 ;
			data[98514] <= 8'h10 ;
			data[98515] <= 8'h10 ;
			data[98516] <= 8'h10 ;
			data[98517] <= 8'h10 ;
			data[98518] <= 8'h10 ;
			data[98519] <= 8'h10 ;
			data[98520] <= 8'h10 ;
			data[98521] <= 8'h10 ;
			data[98522] <= 8'h10 ;
			data[98523] <= 8'h10 ;
			data[98524] <= 8'h10 ;
			data[98525] <= 8'h10 ;
			data[98526] <= 8'h10 ;
			data[98527] <= 8'h10 ;
			data[98528] <= 8'h10 ;
			data[98529] <= 8'h10 ;
			data[98530] <= 8'h10 ;
			data[98531] <= 8'h10 ;
			data[98532] <= 8'h10 ;
			data[98533] <= 8'h10 ;
			data[98534] <= 8'h10 ;
			data[98535] <= 8'h10 ;
			data[98536] <= 8'h10 ;
			data[98537] <= 8'h10 ;
			data[98538] <= 8'h10 ;
			data[98539] <= 8'h10 ;
			data[98540] <= 8'h10 ;
			data[98541] <= 8'h10 ;
			data[98542] <= 8'h10 ;
			data[98543] <= 8'h10 ;
			data[98544] <= 8'h10 ;
			data[98545] <= 8'h10 ;
			data[98546] <= 8'h10 ;
			data[98547] <= 8'h10 ;
			data[98548] <= 8'h10 ;
			data[98549] <= 8'h10 ;
			data[98550] <= 8'h10 ;
			data[98551] <= 8'h10 ;
			data[98552] <= 8'h10 ;
			data[98553] <= 8'h10 ;
			data[98554] <= 8'h10 ;
			data[98555] <= 8'h10 ;
			data[98556] <= 8'h10 ;
			data[98557] <= 8'h10 ;
			data[98558] <= 8'h10 ;
			data[98559] <= 8'h10 ;
			data[98560] <= 8'h10 ;
			data[98561] <= 8'h10 ;
			data[98562] <= 8'h10 ;
			data[98563] <= 8'h10 ;
			data[98564] <= 8'h10 ;
			data[98565] <= 8'h10 ;
			data[98566] <= 8'h10 ;
			data[98567] <= 8'h10 ;
			data[98568] <= 8'h10 ;
			data[98569] <= 8'h10 ;
			data[98570] <= 8'h10 ;
			data[98571] <= 8'h10 ;
			data[98572] <= 8'h10 ;
			data[98573] <= 8'h10 ;
			data[98574] <= 8'h10 ;
			data[98575] <= 8'h10 ;
			data[98576] <= 8'h10 ;
			data[98577] <= 8'h10 ;
			data[98578] <= 8'h10 ;
			data[98579] <= 8'h10 ;
			data[98580] <= 8'h10 ;
			data[98581] <= 8'h10 ;
			data[98582] <= 8'h10 ;
			data[98583] <= 8'h10 ;
			data[98584] <= 8'h10 ;
			data[98585] <= 8'h10 ;
			data[98586] <= 8'h10 ;
			data[98587] <= 8'h10 ;
			data[98588] <= 8'h10 ;
			data[98589] <= 8'h10 ;
			data[98590] <= 8'h10 ;
			data[98591] <= 8'h10 ;
			data[98592] <= 8'h10 ;
			data[98593] <= 8'h10 ;
			data[98594] <= 8'h10 ;
			data[98595] <= 8'h10 ;
			data[98596] <= 8'h10 ;
			data[98597] <= 8'h10 ;
			data[98598] <= 8'h10 ;
			data[98599] <= 8'h10 ;
			data[98600] <= 8'h10 ;
			data[98601] <= 8'h10 ;
			data[98602] <= 8'h10 ;
			data[98603] <= 8'h10 ;
			data[98604] <= 8'h10 ;
			data[98605] <= 8'h10 ;
			data[98606] <= 8'h10 ;
			data[98607] <= 8'h10 ;
			data[98608] <= 8'h10 ;
			data[98609] <= 8'h10 ;
			data[98610] <= 8'h10 ;
			data[98611] <= 8'h10 ;
			data[98612] <= 8'h10 ;
			data[98613] <= 8'h10 ;
			data[98614] <= 8'h10 ;
			data[98615] <= 8'h10 ;
			data[98616] <= 8'h10 ;
			data[98617] <= 8'h10 ;
			data[98618] <= 8'h10 ;
			data[98619] <= 8'h10 ;
			data[98620] <= 8'h10 ;
			data[98621] <= 8'h10 ;
			data[98622] <= 8'h10 ;
			data[98623] <= 8'h10 ;
			data[98624] <= 8'h10 ;
			data[98625] <= 8'h10 ;
			data[98626] <= 8'h10 ;
			data[98627] <= 8'h10 ;
			data[98628] <= 8'h10 ;
			data[98629] <= 8'h10 ;
			data[98630] <= 8'h10 ;
			data[98631] <= 8'h10 ;
			data[98632] <= 8'h10 ;
			data[98633] <= 8'h10 ;
			data[98634] <= 8'h10 ;
			data[98635] <= 8'h10 ;
			data[98636] <= 8'h10 ;
			data[98637] <= 8'h10 ;
			data[98638] <= 8'h10 ;
			data[98639] <= 8'h10 ;
			data[98640] <= 8'h10 ;
			data[98641] <= 8'h10 ;
			data[98642] <= 8'h10 ;
			data[98643] <= 8'h10 ;
			data[98644] <= 8'h10 ;
			data[98645] <= 8'h10 ;
			data[98646] <= 8'h10 ;
			data[98647] <= 8'h10 ;
			data[98648] <= 8'h10 ;
			data[98649] <= 8'h10 ;
			data[98650] <= 8'h10 ;
			data[98651] <= 8'h10 ;
			data[98652] <= 8'h10 ;
			data[98653] <= 8'h10 ;
			data[98654] <= 8'h10 ;
			data[98655] <= 8'h10 ;
			data[98656] <= 8'h10 ;
			data[98657] <= 8'h10 ;
			data[98658] <= 8'h10 ;
			data[98659] <= 8'h10 ;
			data[98660] <= 8'h10 ;
			data[98661] <= 8'h10 ;
			data[98662] <= 8'h10 ;
			data[98663] <= 8'h10 ;
			data[98664] <= 8'h10 ;
			data[98665] <= 8'h10 ;
			data[98666] <= 8'h10 ;
			data[98667] <= 8'h10 ;
			data[98668] <= 8'h10 ;
			data[98669] <= 8'h10 ;
			data[98670] <= 8'h10 ;
			data[98671] <= 8'h10 ;
			data[98672] <= 8'h10 ;
			data[98673] <= 8'h10 ;
			data[98674] <= 8'h10 ;
			data[98675] <= 8'h10 ;
			data[98676] <= 8'h10 ;
			data[98677] <= 8'h10 ;
			data[98678] <= 8'h10 ;
			data[98679] <= 8'h10 ;
			data[98680] <= 8'h10 ;
			data[98681] <= 8'h10 ;
			data[98682] <= 8'h10 ;
			data[98683] <= 8'h10 ;
			data[98684] <= 8'h10 ;
			data[98685] <= 8'h10 ;
			data[98686] <= 8'h10 ;
			data[98687] <= 8'h10 ;
			data[98688] <= 8'h10 ;
			data[98689] <= 8'h10 ;
			data[98690] <= 8'h10 ;
			data[98691] <= 8'h10 ;
			data[98692] <= 8'h10 ;
			data[98693] <= 8'h10 ;
			data[98694] <= 8'h10 ;
			data[98695] <= 8'h10 ;
			data[98696] <= 8'h10 ;
			data[98697] <= 8'h10 ;
			data[98698] <= 8'h10 ;
			data[98699] <= 8'h10 ;
			data[98700] <= 8'h10 ;
			data[98701] <= 8'h10 ;
			data[98702] <= 8'h10 ;
			data[98703] <= 8'h10 ;
			data[98704] <= 8'h10 ;
			data[98705] <= 8'h10 ;
			data[98706] <= 8'h10 ;
			data[98707] <= 8'h10 ;
			data[98708] <= 8'h10 ;
			data[98709] <= 8'h10 ;
			data[98710] <= 8'h10 ;
			data[98711] <= 8'h10 ;
			data[98712] <= 8'h10 ;
			data[98713] <= 8'h10 ;
			data[98714] <= 8'h10 ;
			data[98715] <= 8'h10 ;
			data[98716] <= 8'h10 ;
			data[98717] <= 8'h10 ;
			data[98718] <= 8'h10 ;
			data[98719] <= 8'h10 ;
			data[98720] <= 8'h10 ;
			data[98721] <= 8'h10 ;
			data[98722] <= 8'h10 ;
			data[98723] <= 8'h10 ;
			data[98724] <= 8'h10 ;
			data[98725] <= 8'h10 ;
			data[98726] <= 8'h10 ;
			data[98727] <= 8'h10 ;
			data[98728] <= 8'h10 ;
			data[98729] <= 8'h10 ;
			data[98730] <= 8'h10 ;
			data[98731] <= 8'h10 ;
			data[98732] <= 8'h10 ;
			data[98733] <= 8'h10 ;
			data[98734] <= 8'h10 ;
			data[98735] <= 8'h10 ;
			data[98736] <= 8'h10 ;
			data[98737] <= 8'h10 ;
			data[98738] <= 8'h10 ;
			data[98739] <= 8'h10 ;
			data[98740] <= 8'h10 ;
			data[98741] <= 8'h10 ;
			data[98742] <= 8'h10 ;
			data[98743] <= 8'h10 ;
			data[98744] <= 8'h10 ;
			data[98745] <= 8'h10 ;
			data[98746] <= 8'h10 ;
			data[98747] <= 8'h10 ;
			data[98748] <= 8'h10 ;
			data[98749] <= 8'h10 ;
			data[98750] <= 8'h10 ;
			data[98751] <= 8'h10 ;
			data[98752] <= 8'h10 ;
			data[98753] <= 8'h10 ;
			data[98754] <= 8'h10 ;
			data[98755] <= 8'h10 ;
			data[98756] <= 8'h10 ;
			data[98757] <= 8'h10 ;
			data[98758] <= 8'h10 ;
			data[98759] <= 8'h10 ;
			data[98760] <= 8'h10 ;
			data[98761] <= 8'h10 ;
			data[98762] <= 8'h10 ;
			data[98763] <= 8'h10 ;
			data[98764] <= 8'h10 ;
			data[98765] <= 8'h10 ;
			data[98766] <= 8'h10 ;
			data[98767] <= 8'h10 ;
			data[98768] <= 8'h10 ;
			data[98769] <= 8'h10 ;
			data[98770] <= 8'h10 ;
			data[98771] <= 8'h10 ;
			data[98772] <= 8'h10 ;
			data[98773] <= 8'h10 ;
			data[98774] <= 8'h10 ;
			data[98775] <= 8'h10 ;
			data[98776] <= 8'h10 ;
			data[98777] <= 8'h10 ;
			data[98778] <= 8'h10 ;
			data[98779] <= 8'h10 ;
			data[98780] <= 8'h10 ;
			data[98781] <= 8'h10 ;
			data[98782] <= 8'h10 ;
			data[98783] <= 8'h10 ;
			data[98784] <= 8'h10 ;
			data[98785] <= 8'h10 ;
			data[98786] <= 8'h10 ;
			data[98787] <= 8'h10 ;
			data[98788] <= 8'h10 ;
			data[98789] <= 8'h10 ;
			data[98790] <= 8'h10 ;
			data[98791] <= 8'h10 ;
			data[98792] <= 8'h10 ;
			data[98793] <= 8'h10 ;
			data[98794] <= 8'h10 ;
			data[98795] <= 8'h10 ;
			data[98796] <= 8'h10 ;
			data[98797] <= 8'h10 ;
			data[98798] <= 8'h10 ;
			data[98799] <= 8'h10 ;
			data[98800] <= 8'h10 ;
			data[98801] <= 8'h10 ;
			data[98802] <= 8'h10 ;
			data[98803] <= 8'h10 ;
			data[98804] <= 8'h10 ;
			data[98805] <= 8'h10 ;
			data[98806] <= 8'h10 ;
			data[98807] <= 8'h10 ;
			data[98808] <= 8'h10 ;
			data[98809] <= 8'h10 ;
			data[98810] <= 8'h10 ;
			data[98811] <= 8'h10 ;
			data[98812] <= 8'h10 ;
			data[98813] <= 8'h10 ;
			data[98814] <= 8'h10 ;
			data[98815] <= 8'h10 ;
			data[98816] <= 8'h10 ;
			data[98817] <= 8'h10 ;
			data[98818] <= 8'h10 ;
			data[98819] <= 8'h10 ;
			data[98820] <= 8'h10 ;
			data[98821] <= 8'h10 ;
			data[98822] <= 8'h10 ;
			data[98823] <= 8'h10 ;
			data[98824] <= 8'h10 ;
			data[98825] <= 8'h10 ;
			data[98826] <= 8'h10 ;
			data[98827] <= 8'h10 ;
			data[98828] <= 8'h10 ;
			data[98829] <= 8'h10 ;
			data[98830] <= 8'h10 ;
			data[98831] <= 8'h10 ;
			data[98832] <= 8'h10 ;
			data[98833] <= 8'h10 ;
			data[98834] <= 8'h10 ;
			data[98835] <= 8'h10 ;
			data[98836] <= 8'h10 ;
			data[98837] <= 8'h10 ;
			data[98838] <= 8'h10 ;
			data[98839] <= 8'h10 ;
			data[98840] <= 8'h10 ;
			data[98841] <= 8'h10 ;
			data[98842] <= 8'h10 ;
			data[98843] <= 8'h10 ;
			data[98844] <= 8'h10 ;
			data[98845] <= 8'h10 ;
			data[98846] <= 8'h10 ;
			data[98847] <= 8'h10 ;
			data[98848] <= 8'h10 ;
			data[98849] <= 8'h10 ;
			data[98850] <= 8'h10 ;
			data[98851] <= 8'h10 ;
			data[98852] <= 8'h10 ;
			data[98853] <= 8'h10 ;
			data[98854] <= 8'h10 ;
			data[98855] <= 8'h10 ;
			data[98856] <= 8'h10 ;
			data[98857] <= 8'h10 ;
			data[98858] <= 8'h10 ;
			data[98859] <= 8'h10 ;
			data[98860] <= 8'h10 ;
			data[98861] <= 8'h10 ;
			data[98862] <= 8'h10 ;
			data[98863] <= 8'h10 ;
			data[98864] <= 8'h10 ;
			data[98865] <= 8'h10 ;
			data[98866] <= 8'h10 ;
			data[98867] <= 8'h10 ;
			data[98868] <= 8'h10 ;
			data[98869] <= 8'h10 ;
			data[98870] <= 8'h10 ;
			data[98871] <= 8'h10 ;
			data[98872] <= 8'h10 ;
			data[98873] <= 8'h10 ;
			data[98874] <= 8'h10 ;
			data[98875] <= 8'h10 ;
			data[98876] <= 8'h10 ;
			data[98877] <= 8'h10 ;
			data[98878] <= 8'h10 ;
			data[98879] <= 8'h10 ;
			data[98880] <= 8'h10 ;
			data[98881] <= 8'h10 ;
			data[98882] <= 8'h10 ;
			data[98883] <= 8'h10 ;
			data[98884] <= 8'h10 ;
			data[98885] <= 8'h10 ;
			data[98886] <= 8'h10 ;
			data[98887] <= 8'h10 ;
			data[98888] <= 8'h10 ;
			data[98889] <= 8'h10 ;
			data[98890] <= 8'h10 ;
			data[98891] <= 8'h10 ;
			data[98892] <= 8'h10 ;
			data[98893] <= 8'h10 ;
			data[98894] <= 8'h10 ;
			data[98895] <= 8'h10 ;
			data[98896] <= 8'h10 ;
			data[98897] <= 8'h10 ;
			data[98898] <= 8'h10 ;
			data[98899] <= 8'h10 ;
			data[98900] <= 8'h10 ;
			data[98901] <= 8'h10 ;
			data[98902] <= 8'h10 ;
			data[98903] <= 8'h10 ;
			data[98904] <= 8'h10 ;
			data[98905] <= 8'h10 ;
			data[98906] <= 8'h10 ;
			data[98907] <= 8'h10 ;
			data[98908] <= 8'h10 ;
			data[98909] <= 8'h10 ;
			data[98910] <= 8'h10 ;
			data[98911] <= 8'h10 ;
			data[98912] <= 8'h10 ;
			data[98913] <= 8'h10 ;
			data[98914] <= 8'h10 ;
			data[98915] <= 8'h10 ;
			data[98916] <= 8'h10 ;
			data[98917] <= 8'h10 ;
			data[98918] <= 8'h10 ;
			data[98919] <= 8'h10 ;
			data[98920] <= 8'h10 ;
			data[98921] <= 8'h10 ;
			data[98922] <= 8'h10 ;
			data[98923] <= 8'h10 ;
			data[98924] <= 8'h10 ;
			data[98925] <= 8'h10 ;
			data[98926] <= 8'h10 ;
			data[98927] <= 8'h10 ;
			data[98928] <= 8'h10 ;
			data[98929] <= 8'h10 ;
			data[98930] <= 8'h10 ;
			data[98931] <= 8'h10 ;
			data[98932] <= 8'h10 ;
			data[98933] <= 8'h10 ;
			data[98934] <= 8'h10 ;
			data[98935] <= 8'h10 ;
			data[98936] <= 8'h10 ;
			data[98937] <= 8'h10 ;
			data[98938] <= 8'h10 ;
			data[98939] <= 8'h10 ;
			data[98940] <= 8'h10 ;
			data[98941] <= 8'h10 ;
			data[98942] <= 8'h10 ;
			data[98943] <= 8'h10 ;
			data[98944] <= 8'h10 ;
			data[98945] <= 8'h10 ;
			data[98946] <= 8'h10 ;
			data[98947] <= 8'h10 ;
			data[98948] <= 8'h10 ;
			data[98949] <= 8'h10 ;
			data[98950] <= 8'h10 ;
			data[98951] <= 8'h10 ;
			data[98952] <= 8'h10 ;
			data[98953] <= 8'h10 ;
			data[98954] <= 8'h10 ;
			data[98955] <= 8'h10 ;
			data[98956] <= 8'h10 ;
			data[98957] <= 8'h10 ;
			data[98958] <= 8'h10 ;
			data[98959] <= 8'h10 ;
			data[98960] <= 8'h10 ;
			data[98961] <= 8'h10 ;
			data[98962] <= 8'h10 ;
			data[98963] <= 8'h10 ;
			data[98964] <= 8'h10 ;
			data[98965] <= 8'h10 ;
			data[98966] <= 8'h10 ;
			data[98967] <= 8'h10 ;
			data[98968] <= 8'h10 ;
			data[98969] <= 8'h10 ;
			data[98970] <= 8'h10 ;
			data[98971] <= 8'h10 ;
			data[98972] <= 8'h10 ;
			data[98973] <= 8'h10 ;
			data[98974] <= 8'h10 ;
			data[98975] <= 8'h10 ;
			data[98976] <= 8'h10 ;
			data[98977] <= 8'h10 ;
			data[98978] <= 8'h10 ;
			data[98979] <= 8'h10 ;
			data[98980] <= 8'h10 ;
			data[98981] <= 8'h10 ;
			data[98982] <= 8'h10 ;
			data[98983] <= 8'h10 ;
			data[98984] <= 8'h10 ;
			data[98985] <= 8'h10 ;
			data[98986] <= 8'h10 ;
			data[98987] <= 8'h10 ;
			data[98988] <= 8'h10 ;
			data[98989] <= 8'h10 ;
			data[98990] <= 8'h10 ;
			data[98991] <= 8'h10 ;
			data[98992] <= 8'h10 ;
			data[98993] <= 8'h10 ;
			data[98994] <= 8'h10 ;
			data[98995] <= 8'h10 ;
			data[98996] <= 8'h10 ;
			data[98997] <= 8'h10 ;
			data[98998] <= 8'h10 ;
			data[98999] <= 8'h10 ;
			data[99000] <= 8'h10 ;
			data[99001] <= 8'h10 ;
			data[99002] <= 8'h10 ;
			data[99003] <= 8'h10 ;
			data[99004] <= 8'h10 ;
			data[99005] <= 8'h10 ;
			data[99006] <= 8'h10 ;
			data[99007] <= 8'h10 ;
			data[99008] <= 8'h10 ;
			data[99009] <= 8'h10 ;
			data[99010] <= 8'h10 ;
			data[99011] <= 8'h10 ;
			data[99012] <= 8'h10 ;
			data[99013] <= 8'h10 ;
			data[99014] <= 8'h10 ;
			data[99015] <= 8'h10 ;
			data[99016] <= 8'h10 ;
			data[99017] <= 8'h10 ;
			data[99018] <= 8'h10 ;
			data[99019] <= 8'h10 ;
			data[99020] <= 8'h10 ;
			data[99021] <= 8'h10 ;
			data[99022] <= 8'h10 ;
			data[99023] <= 8'h10 ;
			data[99024] <= 8'h10 ;
			data[99025] <= 8'h10 ;
			data[99026] <= 8'h10 ;
			data[99027] <= 8'h10 ;
			data[99028] <= 8'h10 ;
			data[99029] <= 8'h10 ;
			data[99030] <= 8'h10 ;
			data[99031] <= 8'h10 ;
			data[99032] <= 8'h10 ;
			data[99033] <= 8'h10 ;
			data[99034] <= 8'h10 ;
			data[99035] <= 8'h10 ;
			data[99036] <= 8'h10 ;
			data[99037] <= 8'h10 ;
			data[99038] <= 8'h10 ;
			data[99039] <= 8'h10 ;
			data[99040] <= 8'h10 ;
			data[99041] <= 8'h10 ;
			data[99042] <= 8'h10 ;
			data[99043] <= 8'h10 ;
			data[99044] <= 8'h10 ;
			data[99045] <= 8'h10 ;
			data[99046] <= 8'h10 ;
			data[99047] <= 8'h10 ;
			data[99048] <= 8'h10 ;
			data[99049] <= 8'h10 ;
			data[99050] <= 8'h10 ;
			data[99051] <= 8'h10 ;
			data[99052] <= 8'h10 ;
			data[99053] <= 8'h10 ;
			data[99054] <= 8'h10 ;
			data[99055] <= 8'h10 ;
			data[99056] <= 8'h10 ;
			data[99057] <= 8'h10 ;
			data[99058] <= 8'h10 ;
			data[99059] <= 8'h10 ;
			data[99060] <= 8'h10 ;
			data[99061] <= 8'h10 ;
			data[99062] <= 8'h10 ;
			data[99063] <= 8'h10 ;
			data[99064] <= 8'h10 ;
			data[99065] <= 8'h10 ;
			data[99066] <= 8'h10 ;
			data[99067] <= 8'h10 ;
			data[99068] <= 8'h10 ;
			data[99069] <= 8'h10 ;
			data[99070] <= 8'h10 ;
			data[99071] <= 8'h10 ;
			data[99072] <= 8'h10 ;
			data[99073] <= 8'h10 ;
			data[99074] <= 8'h10 ;
			data[99075] <= 8'h10 ;
			data[99076] <= 8'h10 ;
			data[99077] <= 8'h10 ;
			data[99078] <= 8'h10 ;
			data[99079] <= 8'h10 ;
			data[99080] <= 8'h10 ;
			data[99081] <= 8'h10 ;
			data[99082] <= 8'h10 ;
			data[99083] <= 8'h10 ;
			data[99084] <= 8'h10 ;
			data[99085] <= 8'h10 ;
			data[99086] <= 8'h10 ;
			data[99087] <= 8'h10 ;
			data[99088] <= 8'h10 ;
			data[99089] <= 8'h10 ;
			data[99090] <= 8'h10 ;
			data[99091] <= 8'h10 ;
			data[99092] <= 8'h10 ;
			data[99093] <= 8'h10 ;
			data[99094] <= 8'h10 ;
			data[99095] <= 8'h10 ;
			data[99096] <= 8'h10 ;
			data[99097] <= 8'h10 ;
			data[99098] <= 8'h10 ;
			data[99099] <= 8'h10 ;
			data[99100] <= 8'h10 ;
			data[99101] <= 8'h10 ;
			data[99102] <= 8'h10 ;
			data[99103] <= 8'h10 ;
			data[99104] <= 8'h10 ;
			data[99105] <= 8'h10 ;
			data[99106] <= 8'h10 ;
			data[99107] <= 8'h10 ;
			data[99108] <= 8'h10 ;
			data[99109] <= 8'h10 ;
			data[99110] <= 8'h10 ;
			data[99111] <= 8'h10 ;
			data[99112] <= 8'h10 ;
			data[99113] <= 8'h10 ;
			data[99114] <= 8'h10 ;
			data[99115] <= 8'h10 ;
			data[99116] <= 8'h10 ;
			data[99117] <= 8'h10 ;
			data[99118] <= 8'h10 ;
			data[99119] <= 8'h10 ;
			data[99120] <= 8'h10 ;
			data[99121] <= 8'h10 ;
			data[99122] <= 8'h10 ;
			data[99123] <= 8'h10 ;
			data[99124] <= 8'h10 ;
			data[99125] <= 8'h10 ;
			data[99126] <= 8'h10 ;
			data[99127] <= 8'h10 ;
			data[99128] <= 8'h10 ;
			data[99129] <= 8'h10 ;
			data[99130] <= 8'h10 ;
			data[99131] <= 8'h10 ;
			data[99132] <= 8'h10 ;
			data[99133] <= 8'h10 ;
			data[99134] <= 8'h10 ;
			data[99135] <= 8'h10 ;
			data[99136] <= 8'h10 ;
			data[99137] <= 8'h10 ;
			data[99138] <= 8'h10 ;
			data[99139] <= 8'h10 ;
			data[99140] <= 8'h10 ;
			data[99141] <= 8'h10 ;
			data[99142] <= 8'h10 ;
			data[99143] <= 8'h10 ;
			data[99144] <= 8'h10 ;
			data[99145] <= 8'h10 ;
			data[99146] <= 8'h10 ;
			data[99147] <= 8'h10 ;
			data[99148] <= 8'h10 ;
			data[99149] <= 8'h10 ;
			data[99150] <= 8'h10 ;
			data[99151] <= 8'h10 ;
			data[99152] <= 8'h10 ;
			data[99153] <= 8'h10 ;
			data[99154] <= 8'h10 ;
			data[99155] <= 8'h10 ;
			data[99156] <= 8'h10 ;
			data[99157] <= 8'h10 ;
			data[99158] <= 8'h10 ;
			data[99159] <= 8'h10 ;
			data[99160] <= 8'h10 ;
			data[99161] <= 8'h10 ;
			data[99162] <= 8'h10 ;
			data[99163] <= 8'h10 ;
			data[99164] <= 8'h10 ;
			data[99165] <= 8'h10 ;
			data[99166] <= 8'h10 ;
			data[99167] <= 8'h10 ;
			data[99168] <= 8'h10 ;
			data[99169] <= 8'h10 ;
			data[99170] <= 8'h10 ;
			data[99171] <= 8'h10 ;
			data[99172] <= 8'h10 ;
			data[99173] <= 8'h10 ;
			data[99174] <= 8'h10 ;
			data[99175] <= 8'h10 ;
			data[99176] <= 8'h10 ;
			data[99177] <= 8'h10 ;
			data[99178] <= 8'h10 ;
			data[99179] <= 8'h10 ;
			data[99180] <= 8'h10 ;
			data[99181] <= 8'h10 ;
			data[99182] <= 8'h10 ;
			data[99183] <= 8'h10 ;
			data[99184] <= 8'h10 ;
			data[99185] <= 8'h10 ;
			data[99186] <= 8'h10 ;
			data[99187] <= 8'h10 ;
			data[99188] <= 8'h10 ;
			data[99189] <= 8'h10 ;
			data[99190] <= 8'h10 ;
			data[99191] <= 8'h10 ;
			data[99192] <= 8'h10 ;
			data[99193] <= 8'h10 ;
			data[99194] <= 8'h10 ;
			data[99195] <= 8'h10 ;
			data[99196] <= 8'h10 ;
			data[99197] <= 8'h10 ;
			data[99198] <= 8'h10 ;
			data[99199] <= 8'h10 ;
			data[99200] <= 8'h10 ;
			data[99201] <= 8'h10 ;
			data[99202] <= 8'h10 ;
			data[99203] <= 8'h10 ;
			data[99204] <= 8'h10 ;
			data[99205] <= 8'h10 ;
			data[99206] <= 8'h10 ;
			data[99207] <= 8'h10 ;
			data[99208] <= 8'h10 ;
			data[99209] <= 8'h10 ;
			data[99210] <= 8'h10 ;
			data[99211] <= 8'h10 ;
			data[99212] <= 8'h10 ;
			data[99213] <= 8'h10 ;
			data[99214] <= 8'h10 ;
			data[99215] <= 8'h10 ;
			data[99216] <= 8'h10 ;
			data[99217] <= 8'h10 ;
			data[99218] <= 8'h10 ;
			data[99219] <= 8'h10 ;
			data[99220] <= 8'h10 ;
			data[99221] <= 8'h10 ;
			data[99222] <= 8'h10 ;
			data[99223] <= 8'h10 ;
			data[99224] <= 8'h10 ;
			data[99225] <= 8'h10 ;
			data[99226] <= 8'h10 ;
			data[99227] <= 8'h10 ;
			data[99228] <= 8'h10 ;
			data[99229] <= 8'h10 ;
			data[99230] <= 8'h10 ;
			data[99231] <= 8'h10 ;
			data[99232] <= 8'h10 ;
			data[99233] <= 8'h10 ;
			data[99234] <= 8'h10 ;
			data[99235] <= 8'h10 ;
			data[99236] <= 8'h10 ;
			data[99237] <= 8'h10 ;
			data[99238] <= 8'h10 ;
			data[99239] <= 8'h10 ;
			data[99240] <= 8'h10 ;
			data[99241] <= 8'h10 ;
			data[99242] <= 8'h10 ;
			data[99243] <= 8'h10 ;
			data[99244] <= 8'h10 ;
			data[99245] <= 8'h10 ;
			data[99246] <= 8'h10 ;
			data[99247] <= 8'h10 ;
			data[99248] <= 8'h10 ;
			data[99249] <= 8'h10 ;
			data[99250] <= 8'h10 ;
			data[99251] <= 8'h10 ;
			data[99252] <= 8'h10 ;
			data[99253] <= 8'h10 ;
			data[99254] <= 8'h10 ;
			data[99255] <= 8'h10 ;
			data[99256] <= 8'h10 ;
			data[99257] <= 8'h10 ;
			data[99258] <= 8'h10 ;
			data[99259] <= 8'h10 ;
			data[99260] <= 8'h10 ;
			data[99261] <= 8'h10 ;
			data[99262] <= 8'h10 ;
			data[99263] <= 8'h10 ;
			data[99264] <= 8'h10 ;
			data[99265] <= 8'h10 ;
			data[99266] <= 8'h10 ;
			data[99267] <= 8'h10 ;
			data[99268] <= 8'h10 ;
			data[99269] <= 8'h10 ;
			data[99270] <= 8'h10 ;
			data[99271] <= 8'h10 ;
			data[99272] <= 8'h10 ;
			data[99273] <= 8'h10 ;
			data[99274] <= 8'h10 ;
			data[99275] <= 8'h10 ;
			data[99276] <= 8'h10 ;
			data[99277] <= 8'h10 ;
			data[99278] <= 8'h10 ;
			data[99279] <= 8'h10 ;
			data[99280] <= 8'h10 ;
			data[99281] <= 8'h10 ;
			data[99282] <= 8'h10 ;
			data[99283] <= 8'h10 ;
			data[99284] <= 8'h10 ;
			data[99285] <= 8'h10 ;
			data[99286] <= 8'h10 ;
			data[99287] <= 8'h10 ;
			data[99288] <= 8'h10 ;
			data[99289] <= 8'h10 ;
			data[99290] <= 8'h10 ;
			data[99291] <= 8'h10 ;
			data[99292] <= 8'h10 ;
			data[99293] <= 8'h10 ;
			data[99294] <= 8'h10 ;
			data[99295] <= 8'h10 ;
			data[99296] <= 8'h10 ;
			data[99297] <= 8'h10 ;
			data[99298] <= 8'h10 ;
			data[99299] <= 8'h10 ;
			data[99300] <= 8'h10 ;
			data[99301] <= 8'h10 ;
			data[99302] <= 8'h10 ;
			data[99303] <= 8'h10 ;
			data[99304] <= 8'h10 ;
			data[99305] <= 8'h10 ;
			data[99306] <= 8'h10 ;
			data[99307] <= 8'h10 ;
			data[99308] <= 8'h10 ;
			data[99309] <= 8'h10 ;
			data[99310] <= 8'h10 ;
			data[99311] <= 8'h10 ;
			data[99312] <= 8'h10 ;
			data[99313] <= 8'h10 ;
			data[99314] <= 8'h10 ;
			data[99315] <= 8'h10 ;
			data[99316] <= 8'h10 ;
			data[99317] <= 8'h10 ;
			data[99318] <= 8'h10 ;
			data[99319] <= 8'h10 ;
			data[99320] <= 8'h10 ;
			data[99321] <= 8'h10 ;
			data[99322] <= 8'h10 ;
			data[99323] <= 8'h10 ;
			data[99324] <= 8'h10 ;
			data[99325] <= 8'h10 ;
			data[99326] <= 8'h10 ;
			data[99327] <= 8'h10 ;
			data[99328] <= 8'h10 ;
			data[99329] <= 8'h10 ;
			data[99330] <= 8'h10 ;
			data[99331] <= 8'h10 ;
			data[99332] <= 8'h10 ;
			data[99333] <= 8'h10 ;
			data[99334] <= 8'h10 ;
			data[99335] <= 8'h10 ;
			data[99336] <= 8'h10 ;
			data[99337] <= 8'h10 ;
			data[99338] <= 8'h10 ;
			data[99339] <= 8'h10 ;
			data[99340] <= 8'h10 ;
			data[99341] <= 8'h10 ;
			data[99342] <= 8'h10 ;
			data[99343] <= 8'h10 ;
			data[99344] <= 8'h10 ;
			data[99345] <= 8'h10 ;
			data[99346] <= 8'h10 ;
			data[99347] <= 8'h10 ;
			data[99348] <= 8'h10 ;
			data[99349] <= 8'h10 ;
			data[99350] <= 8'h10 ;
			data[99351] <= 8'h10 ;
			data[99352] <= 8'h10 ;
			data[99353] <= 8'h10 ;
			data[99354] <= 8'h10 ;
			data[99355] <= 8'h10 ;
			data[99356] <= 8'h10 ;
			data[99357] <= 8'h10 ;
			data[99358] <= 8'h10 ;
			data[99359] <= 8'h10 ;
			data[99360] <= 8'h10 ;
			data[99361] <= 8'h10 ;
			data[99362] <= 8'h10 ;
			data[99363] <= 8'h10 ;
			data[99364] <= 8'h10 ;
			data[99365] <= 8'h10 ;
			data[99366] <= 8'h10 ;
			data[99367] <= 8'h10 ;
			data[99368] <= 8'h10 ;
			data[99369] <= 8'h10 ;
			data[99370] <= 8'h10 ;
			data[99371] <= 8'h10 ;
			data[99372] <= 8'h10 ;
			data[99373] <= 8'h10 ;
			data[99374] <= 8'h10 ;
			data[99375] <= 8'h10 ;
			data[99376] <= 8'h10 ;
			data[99377] <= 8'h10 ;
			data[99378] <= 8'h10 ;
			data[99379] <= 8'h10 ;
			data[99380] <= 8'h10 ;
			data[99381] <= 8'h10 ;
			data[99382] <= 8'h10 ;
			data[99383] <= 8'h10 ;
			data[99384] <= 8'h10 ;
			data[99385] <= 8'h10 ;
			data[99386] <= 8'h10 ;
			data[99387] <= 8'h10 ;
			data[99388] <= 8'h10 ;
			data[99389] <= 8'h10 ;
			data[99390] <= 8'h10 ;
			data[99391] <= 8'h10 ;
			data[99392] <= 8'h10 ;
			data[99393] <= 8'h10 ;
			data[99394] <= 8'h10 ;
			data[99395] <= 8'h10 ;
			data[99396] <= 8'h10 ;
			data[99397] <= 8'h10 ;
			data[99398] <= 8'h10 ;
			data[99399] <= 8'h10 ;
			data[99400] <= 8'h10 ;
			data[99401] <= 8'h10 ;
			data[99402] <= 8'h10 ;
			data[99403] <= 8'h10 ;
			data[99404] <= 8'h10 ;
			data[99405] <= 8'h10 ;
			data[99406] <= 8'h10 ;
			data[99407] <= 8'h10 ;
			data[99408] <= 8'h10 ;
			data[99409] <= 8'h10 ;
			data[99410] <= 8'h10 ;
			data[99411] <= 8'h10 ;
			data[99412] <= 8'h10 ;
			data[99413] <= 8'h10 ;
			data[99414] <= 8'h10 ;
			data[99415] <= 8'h10 ;
			data[99416] <= 8'h10 ;
			data[99417] <= 8'h10 ;
			data[99418] <= 8'h10 ;
			data[99419] <= 8'h10 ;
			data[99420] <= 8'h10 ;
			data[99421] <= 8'h10 ;
			data[99422] <= 8'h10 ;
			data[99423] <= 8'h10 ;
			data[99424] <= 8'h10 ;
			data[99425] <= 8'h10 ;
			data[99426] <= 8'h10 ;
			data[99427] <= 8'h10 ;
			data[99428] <= 8'h10 ;
			data[99429] <= 8'h10 ;
			data[99430] <= 8'h10 ;
			data[99431] <= 8'h10 ;
			data[99432] <= 8'h10 ;
			data[99433] <= 8'h10 ;
			data[99434] <= 8'h10 ;
			data[99435] <= 8'h10 ;
			data[99436] <= 8'h10 ;
			data[99437] <= 8'h10 ;
			data[99438] <= 8'h10 ;
			data[99439] <= 8'h10 ;
			data[99440] <= 8'h10 ;
			data[99441] <= 8'h10 ;
			data[99442] <= 8'h10 ;
			data[99443] <= 8'h10 ;
			data[99444] <= 8'h10 ;
			data[99445] <= 8'h10 ;
			data[99446] <= 8'h10 ;
			data[99447] <= 8'h10 ;
			data[99448] <= 8'h10 ;
			data[99449] <= 8'h10 ;
			data[99450] <= 8'h10 ;
			data[99451] <= 8'h10 ;
			data[99452] <= 8'h10 ;
			data[99453] <= 8'h10 ;
			data[99454] <= 8'h10 ;
			data[99455] <= 8'h10 ;
			data[99456] <= 8'h10 ;
			data[99457] <= 8'h10 ;
			data[99458] <= 8'h10 ;
			data[99459] <= 8'h10 ;
			data[99460] <= 8'h10 ;
			data[99461] <= 8'h10 ;
			data[99462] <= 8'h10 ;
			data[99463] <= 8'h10 ;
			data[99464] <= 8'h10 ;
			data[99465] <= 8'h10 ;
			data[99466] <= 8'h10 ;
			data[99467] <= 8'h10 ;
			data[99468] <= 8'h10 ;
			data[99469] <= 8'h10 ;
			data[99470] <= 8'h10 ;
			data[99471] <= 8'h10 ;
			data[99472] <= 8'h10 ;
			data[99473] <= 8'h10 ;
			data[99474] <= 8'h10 ;
			data[99475] <= 8'h10 ;
			data[99476] <= 8'h10 ;
			data[99477] <= 8'h10 ;
			data[99478] <= 8'h10 ;
			data[99479] <= 8'h10 ;
			data[99480] <= 8'h10 ;
			data[99481] <= 8'h10 ;
			data[99482] <= 8'h10 ;
			data[99483] <= 8'h10 ;
			data[99484] <= 8'h10 ;
			data[99485] <= 8'h10 ;
			data[99486] <= 8'h10 ;
			data[99487] <= 8'h10 ;
			data[99488] <= 8'h10 ;
			data[99489] <= 8'h10 ;
			data[99490] <= 8'h10 ;
			data[99491] <= 8'h10 ;
			data[99492] <= 8'h10 ;
			data[99493] <= 8'h10 ;
			data[99494] <= 8'h10 ;
			data[99495] <= 8'h10 ;
			data[99496] <= 8'h10 ;
			data[99497] <= 8'h10 ;
			data[99498] <= 8'h10 ;
			data[99499] <= 8'h10 ;
			data[99500] <= 8'h10 ;
			data[99501] <= 8'h10 ;
			data[99502] <= 8'h10 ;
			data[99503] <= 8'h10 ;
			data[99504] <= 8'h10 ;
			data[99505] <= 8'h10 ;
			data[99506] <= 8'h10 ;
			data[99507] <= 8'h10 ;
			data[99508] <= 8'h10 ;
			data[99509] <= 8'h10 ;
			data[99510] <= 8'h10 ;
			data[99511] <= 8'h10 ;
			data[99512] <= 8'h10 ;
			data[99513] <= 8'h10 ;
			data[99514] <= 8'h10 ;
			data[99515] <= 8'h10 ;
			data[99516] <= 8'h10 ;
			data[99517] <= 8'h10 ;
			data[99518] <= 8'h10 ;
			data[99519] <= 8'h10 ;
			data[99520] <= 8'h10 ;
			data[99521] <= 8'h10 ;
			data[99522] <= 8'h10 ;
			data[99523] <= 8'h10 ;
			data[99524] <= 8'h10 ;
			data[99525] <= 8'h10 ;
			data[99526] <= 8'h10 ;
			data[99527] <= 8'h10 ;
			data[99528] <= 8'h10 ;
			data[99529] <= 8'h10 ;
			data[99530] <= 8'h10 ;
			data[99531] <= 8'h10 ;
			data[99532] <= 8'h10 ;
			data[99533] <= 8'h10 ;
			data[99534] <= 8'h10 ;
			data[99535] <= 8'h10 ;
			data[99536] <= 8'h10 ;
			data[99537] <= 8'h10 ;
			data[99538] <= 8'h10 ;
			data[99539] <= 8'h10 ;
			data[99540] <= 8'h10 ;
			data[99541] <= 8'h10 ;
			data[99542] <= 8'h10 ;
			data[99543] <= 8'h10 ;
			data[99544] <= 8'h10 ;
			data[99545] <= 8'h10 ;
			data[99546] <= 8'h10 ;
			data[99547] <= 8'h10 ;
			data[99548] <= 8'h10 ;
			data[99549] <= 8'h10 ;
			data[99550] <= 8'h10 ;
			data[99551] <= 8'h10 ;
			data[99552] <= 8'h10 ;
			data[99553] <= 8'h10 ;
			data[99554] <= 8'h10 ;
			data[99555] <= 8'h10 ;
			data[99556] <= 8'h10 ;
			data[99557] <= 8'h10 ;
			data[99558] <= 8'h10 ;
			data[99559] <= 8'h10 ;
			data[99560] <= 8'h10 ;
			data[99561] <= 8'h10 ;
			data[99562] <= 8'h10 ;
			data[99563] <= 8'h10 ;
			data[99564] <= 8'h10 ;
			data[99565] <= 8'h10 ;
			data[99566] <= 8'h10 ;
			data[99567] <= 8'h10 ;
			data[99568] <= 8'h10 ;
			data[99569] <= 8'h10 ;
			data[99570] <= 8'h10 ;
			data[99571] <= 8'h10 ;
			data[99572] <= 8'h10 ;
			data[99573] <= 8'h10 ;
			data[99574] <= 8'h10 ;
			data[99575] <= 8'h10 ;
			data[99576] <= 8'h10 ;
			data[99577] <= 8'h10 ;
			data[99578] <= 8'h10 ;
			data[99579] <= 8'h10 ;
			data[99580] <= 8'h10 ;
			data[99581] <= 8'h10 ;
			data[99582] <= 8'h10 ;
			data[99583] <= 8'h10 ;
			data[99584] <= 8'h10 ;
			data[99585] <= 8'h10 ;
			data[99586] <= 8'h10 ;
			data[99587] <= 8'h10 ;
			data[99588] <= 8'h10 ;
			data[99589] <= 8'h10 ;
			data[99590] <= 8'h10 ;
			data[99591] <= 8'h10 ;
			data[99592] <= 8'h10 ;
			data[99593] <= 8'h10 ;
			data[99594] <= 8'h10 ;
			data[99595] <= 8'h10 ;
			data[99596] <= 8'h10 ;
			data[99597] <= 8'h10 ;
			data[99598] <= 8'h10 ;
			data[99599] <= 8'h10 ;
			data[99600] <= 8'h10 ;
			data[99601] <= 8'h10 ;
			data[99602] <= 8'h10 ;
			data[99603] <= 8'h10 ;
			data[99604] <= 8'h10 ;
			data[99605] <= 8'h10 ;
			data[99606] <= 8'h10 ;
			data[99607] <= 8'h10 ;
			data[99608] <= 8'h10 ;
			data[99609] <= 8'h10 ;
			data[99610] <= 8'h10 ;
			data[99611] <= 8'h10 ;
			data[99612] <= 8'h10 ;
			data[99613] <= 8'h10 ;
			data[99614] <= 8'h10 ;
			data[99615] <= 8'h10 ;
			data[99616] <= 8'h10 ;
			data[99617] <= 8'h10 ;
			data[99618] <= 8'h10 ;
			data[99619] <= 8'h10 ;
			data[99620] <= 8'h10 ;
			data[99621] <= 8'h10 ;
			data[99622] <= 8'h10 ;
			data[99623] <= 8'h10 ;
			data[99624] <= 8'h10 ;
			data[99625] <= 8'h10 ;
			data[99626] <= 8'h10 ;
			data[99627] <= 8'h10 ;
			data[99628] <= 8'h10 ;
			data[99629] <= 8'h10 ;
			data[99630] <= 8'h10 ;
			data[99631] <= 8'h10 ;
			data[99632] <= 8'h10 ;
			data[99633] <= 8'h10 ;
			data[99634] <= 8'h10 ;
			data[99635] <= 8'h10 ;
			data[99636] <= 8'h10 ;
			data[99637] <= 8'h10 ;
			data[99638] <= 8'h10 ;
			data[99639] <= 8'h10 ;
			data[99640] <= 8'h10 ;
			data[99641] <= 8'h10 ;
			data[99642] <= 8'h10 ;
			data[99643] <= 8'h10 ;
			data[99644] <= 8'h10 ;
			data[99645] <= 8'h10 ;
			data[99646] <= 8'h10 ;
			data[99647] <= 8'h10 ;
			data[99648] <= 8'h10 ;
			data[99649] <= 8'h10 ;
			data[99650] <= 8'h10 ;
			data[99651] <= 8'h10 ;
			data[99652] <= 8'h10 ;
			data[99653] <= 8'h10 ;
			data[99654] <= 8'h10 ;
			data[99655] <= 8'h10 ;
			data[99656] <= 8'h10 ;
			data[99657] <= 8'h10 ;
			data[99658] <= 8'h10 ;
			data[99659] <= 8'h10 ;
			data[99660] <= 8'h10 ;
			data[99661] <= 8'h10 ;
			data[99662] <= 8'h10 ;
			data[99663] <= 8'h10 ;
			data[99664] <= 8'h10 ;
			data[99665] <= 8'h10 ;
			data[99666] <= 8'h10 ;
			data[99667] <= 8'h10 ;
			data[99668] <= 8'h10 ;
			data[99669] <= 8'h10 ;
			data[99670] <= 8'h10 ;
			data[99671] <= 8'h10 ;
			data[99672] <= 8'h10 ;
			data[99673] <= 8'h10 ;
			data[99674] <= 8'h10 ;
			data[99675] <= 8'h10 ;
			data[99676] <= 8'h10 ;
			data[99677] <= 8'h10 ;
			data[99678] <= 8'h10 ;
			data[99679] <= 8'h10 ;
			data[99680] <= 8'h10 ;
			data[99681] <= 8'h10 ;
			data[99682] <= 8'h10 ;
			data[99683] <= 8'h10 ;
			data[99684] <= 8'h10 ;
			data[99685] <= 8'h10 ;
			data[99686] <= 8'h10 ;
			data[99687] <= 8'h10 ;
			data[99688] <= 8'h10 ;
			data[99689] <= 8'h10 ;
			data[99690] <= 8'h10 ;
			data[99691] <= 8'h10 ;
			data[99692] <= 8'h10 ;
			data[99693] <= 8'h10 ;
			data[99694] <= 8'h10 ;
			data[99695] <= 8'h10 ;
			data[99696] <= 8'h10 ;
			data[99697] <= 8'h10 ;
			data[99698] <= 8'h10 ;
			data[99699] <= 8'h10 ;
			data[99700] <= 8'h10 ;
			data[99701] <= 8'h10 ;
			data[99702] <= 8'h10 ;
			data[99703] <= 8'h10 ;
			data[99704] <= 8'h10 ;
			data[99705] <= 8'h10 ;
			data[99706] <= 8'h10 ;
			data[99707] <= 8'h10 ;
			data[99708] <= 8'h10 ;
			data[99709] <= 8'h10 ;
			data[99710] <= 8'h10 ;
			data[99711] <= 8'h10 ;
			data[99712] <= 8'h10 ;
			data[99713] <= 8'h10 ;
			data[99714] <= 8'h10 ;
			data[99715] <= 8'h10 ;
			data[99716] <= 8'h10 ;
			data[99717] <= 8'h10 ;
			data[99718] <= 8'h10 ;
			data[99719] <= 8'h10 ;
			data[99720] <= 8'h10 ;
			data[99721] <= 8'h10 ;
			data[99722] <= 8'h10 ;
			data[99723] <= 8'h10 ;
			data[99724] <= 8'h10 ;
			data[99725] <= 8'h10 ;
			data[99726] <= 8'h10 ;
			data[99727] <= 8'h10 ;
			data[99728] <= 8'h10 ;
			data[99729] <= 8'h10 ;
			data[99730] <= 8'h10 ;
			data[99731] <= 8'h10 ;
			data[99732] <= 8'h10 ;
			data[99733] <= 8'h10 ;
			data[99734] <= 8'h10 ;
			data[99735] <= 8'h10 ;
			data[99736] <= 8'h10 ;
			data[99737] <= 8'h10 ;
			data[99738] <= 8'h10 ;
			data[99739] <= 8'h10 ;
			data[99740] <= 8'h10 ;
			data[99741] <= 8'h10 ;
			data[99742] <= 8'h10 ;
			data[99743] <= 8'h10 ;
			data[99744] <= 8'h10 ;
			data[99745] <= 8'h10 ;
			data[99746] <= 8'h10 ;
			data[99747] <= 8'h10 ;
			data[99748] <= 8'h10 ;
			data[99749] <= 8'h10 ;
			data[99750] <= 8'h10 ;
			data[99751] <= 8'h10 ;
			data[99752] <= 8'h10 ;
			data[99753] <= 8'h10 ;
			data[99754] <= 8'h10 ;
			data[99755] <= 8'h10 ;
			data[99756] <= 8'h10 ;
			data[99757] <= 8'h10 ;
			data[99758] <= 8'h10 ;
			data[99759] <= 8'h10 ;
			data[99760] <= 8'h10 ;
			data[99761] <= 8'h10 ;
			data[99762] <= 8'h10 ;
			data[99763] <= 8'h10 ;
			data[99764] <= 8'h10 ;
			data[99765] <= 8'h10 ;
			data[99766] <= 8'h10 ;
			data[99767] <= 8'h10 ;
			data[99768] <= 8'h10 ;
			data[99769] <= 8'h10 ;
			data[99770] <= 8'h10 ;
			data[99771] <= 8'h10 ;
			data[99772] <= 8'h10 ;
			data[99773] <= 8'h10 ;
			data[99774] <= 8'h10 ;
			data[99775] <= 8'h10 ;
			data[99776] <= 8'h10 ;
			data[99777] <= 8'h10 ;
			data[99778] <= 8'h10 ;
			data[99779] <= 8'h10 ;
			data[99780] <= 8'h10 ;
			data[99781] <= 8'h10 ;
			data[99782] <= 8'h10 ;
			data[99783] <= 8'h10 ;
			data[99784] <= 8'h10 ;
			data[99785] <= 8'h10 ;
			data[99786] <= 8'h10 ;
			data[99787] <= 8'h10 ;
			data[99788] <= 8'h10 ;
			data[99789] <= 8'h10 ;
			data[99790] <= 8'h10 ;
			data[99791] <= 8'h10 ;
			data[99792] <= 8'h10 ;
			data[99793] <= 8'h10 ;
			data[99794] <= 8'h10 ;
			data[99795] <= 8'h10 ;
			data[99796] <= 8'h10 ;
			data[99797] <= 8'h10 ;
			data[99798] <= 8'h10 ;
			data[99799] <= 8'h10 ;
			data[99800] <= 8'h10 ;
			data[99801] <= 8'h10 ;
			data[99802] <= 8'h10 ;
			data[99803] <= 8'h10 ;
			data[99804] <= 8'h10 ;
			data[99805] <= 8'h10 ;
			data[99806] <= 8'h10 ;
			data[99807] <= 8'h10 ;
			data[99808] <= 8'h10 ;
			data[99809] <= 8'h10 ;
			data[99810] <= 8'h10 ;
			data[99811] <= 8'h10 ;
			data[99812] <= 8'h10 ;
			data[99813] <= 8'h10 ;
			data[99814] <= 8'h10 ;
			data[99815] <= 8'h10 ;
			data[99816] <= 8'h10 ;
			data[99817] <= 8'h10 ;
			data[99818] <= 8'h10 ;
			data[99819] <= 8'h10 ;
			data[99820] <= 8'h10 ;
			data[99821] <= 8'h10 ;
			data[99822] <= 8'h10 ;
			data[99823] <= 8'h10 ;
			data[99824] <= 8'h10 ;
			data[99825] <= 8'h10 ;
			data[99826] <= 8'h10 ;
			data[99827] <= 8'h10 ;
			data[99828] <= 8'h10 ;
			data[99829] <= 8'h10 ;
			data[99830] <= 8'h10 ;
			data[99831] <= 8'h10 ;
			data[99832] <= 8'h10 ;
			data[99833] <= 8'h10 ;
			data[99834] <= 8'h10 ;
			data[99835] <= 8'h10 ;
			data[99836] <= 8'h10 ;
			data[99837] <= 8'h10 ;
			data[99838] <= 8'h10 ;
			data[99839] <= 8'h10 ;
			data[99840] <= 8'h10 ;
			data[99841] <= 8'h10 ;
			data[99842] <= 8'h10 ;
			data[99843] <= 8'h10 ;
			data[99844] <= 8'h10 ;
			data[99845] <= 8'h10 ;
			data[99846] <= 8'h10 ;
			data[99847] <= 8'h10 ;
			data[99848] <= 8'h10 ;
			data[99849] <= 8'h10 ;
			data[99850] <= 8'h10 ;
			data[99851] <= 8'h10 ;
			data[99852] <= 8'h10 ;
			data[99853] <= 8'h10 ;
			data[99854] <= 8'h10 ;
			data[99855] <= 8'h10 ;
			data[99856] <= 8'h10 ;
			data[99857] <= 8'h10 ;
			data[99858] <= 8'h10 ;
			data[99859] <= 8'h10 ;
			data[99860] <= 8'h10 ;
			data[99861] <= 8'h10 ;
			data[99862] <= 8'h10 ;
			data[99863] <= 8'h10 ;
			data[99864] <= 8'h10 ;
			data[99865] <= 8'h10 ;
			data[99866] <= 8'h10 ;
			data[99867] <= 8'h10 ;
			data[99868] <= 8'h10 ;
			data[99869] <= 8'h10 ;
			data[99870] <= 8'h10 ;
			data[99871] <= 8'h10 ;
			data[99872] <= 8'h10 ;
			data[99873] <= 8'h10 ;
			data[99874] <= 8'h10 ;
			data[99875] <= 8'h10 ;
			data[99876] <= 8'h10 ;
			data[99877] <= 8'h10 ;
			data[99878] <= 8'h10 ;
			data[99879] <= 8'h10 ;
			data[99880] <= 8'h10 ;
			data[99881] <= 8'h10 ;
			data[99882] <= 8'h10 ;
			data[99883] <= 8'h10 ;
			data[99884] <= 8'h10 ;
			data[99885] <= 8'h10 ;
			data[99886] <= 8'h10 ;
			data[99887] <= 8'h10 ;
			data[99888] <= 8'h10 ;
			data[99889] <= 8'h10 ;
			data[99890] <= 8'h10 ;
			data[99891] <= 8'h10 ;
			data[99892] <= 8'h10 ;
			data[99893] <= 8'h10 ;
			data[99894] <= 8'h10 ;
			data[99895] <= 8'h10 ;
			data[99896] <= 8'h10 ;
			data[99897] <= 8'h10 ;
			data[99898] <= 8'h10 ;
			data[99899] <= 8'h10 ;
			data[99900] <= 8'h10 ;
			data[99901] <= 8'h10 ;
			data[99902] <= 8'h10 ;
			data[99903] <= 8'h10 ;
			data[99904] <= 8'h10 ;
			data[99905] <= 8'h10 ;
			data[99906] <= 8'h10 ;
			data[99907] <= 8'h10 ;
			data[99908] <= 8'h10 ;
			data[99909] <= 8'h10 ;
			data[99910] <= 8'h10 ;
			data[99911] <= 8'h10 ;
			data[99912] <= 8'h10 ;
			data[99913] <= 8'h10 ;
			data[99914] <= 8'h10 ;
			data[99915] <= 8'h10 ;
			data[99916] <= 8'h10 ;
			data[99917] <= 8'h10 ;
			data[99918] <= 8'h10 ;
			data[99919] <= 8'h10 ;
			data[99920] <= 8'h10 ;
			data[99921] <= 8'h10 ;
			data[99922] <= 8'h10 ;
			data[99923] <= 8'h10 ;
			data[99924] <= 8'h10 ;
			data[99925] <= 8'h10 ;
			data[99926] <= 8'h10 ;
			data[99927] <= 8'h10 ;
			data[99928] <= 8'h10 ;
			data[99929] <= 8'h10 ;
			data[99930] <= 8'h10 ;
			data[99931] <= 8'h10 ;
			data[99932] <= 8'h10 ;
			data[99933] <= 8'h10 ;
			data[99934] <= 8'h10 ;
			data[99935] <= 8'h10 ;
			data[99936] <= 8'h10 ;
			data[99937] <= 8'h10 ;
			data[99938] <= 8'h10 ;
			data[99939] <= 8'h10 ;
			data[99940] <= 8'h10 ;
			data[99941] <= 8'h10 ;
			data[99942] <= 8'h10 ;
			data[99943] <= 8'h10 ;
			data[99944] <= 8'h10 ;
			data[99945] <= 8'h10 ;
			data[99946] <= 8'h10 ;
			data[99947] <= 8'h10 ;
			data[99948] <= 8'h10 ;
			data[99949] <= 8'h10 ;
			data[99950] <= 8'h10 ;
			data[99951] <= 8'h10 ;
			data[99952] <= 8'h10 ;
			data[99953] <= 8'h10 ;
			data[99954] <= 8'h10 ;
			data[99955] <= 8'h10 ;
			data[99956] <= 8'h10 ;
			data[99957] <= 8'h10 ;
			data[99958] <= 8'h10 ;
			data[99959] <= 8'h10 ;
			data[99960] <= 8'h10 ;
			data[99961] <= 8'h10 ;
			data[99962] <= 8'h10 ;
			data[99963] <= 8'h10 ;
			data[99964] <= 8'h10 ;
			data[99965] <= 8'h10 ;
			data[99966] <= 8'h10 ;
			data[99967] <= 8'h10 ;
			data[99968] <= 8'h10 ;
			data[99969] <= 8'h10 ;
			data[99970] <= 8'h10 ;
			data[99971] <= 8'h10 ;
			data[99972] <= 8'h10 ;
			data[99973] <= 8'h10 ;
			data[99974] <= 8'h10 ;
			data[99975] <= 8'h10 ;
			data[99976] <= 8'h10 ;
			data[99977] <= 8'h10 ;
			data[99978] <= 8'h10 ;
			data[99979] <= 8'h10 ;
			data[99980] <= 8'h10 ;
			data[99981] <= 8'h10 ;
			data[99982] <= 8'h10 ;
			data[99983] <= 8'h10 ;
			data[99984] <= 8'h10 ;
			data[99985] <= 8'h10 ;
			data[99986] <= 8'h10 ;
			data[99987] <= 8'h10 ;
			data[99988] <= 8'h10 ;
			data[99989] <= 8'h10 ;
			data[99990] <= 8'h10 ;
			data[99991] <= 8'h10 ;
			data[99992] <= 8'h10 ;
			data[99993] <= 8'h10 ;
			data[99994] <= 8'h10 ;
			data[99995] <= 8'h10 ;
			data[99996] <= 8'h10 ;
			data[99997] <= 8'h10 ;
			data[99998] <= 8'h10 ;
			data[99999] <= 8'h10 ;
			data[100000] <= 8'h10 ;
			data[100001] <= 8'h10 ;
			data[100002] <= 8'h10 ;
			data[100003] <= 8'h10 ;
			data[100004] <= 8'h10 ;
			data[100005] <= 8'h10 ;
			data[100006] <= 8'h10 ;
			data[100007] <= 8'h10 ;
			data[100008] <= 8'h10 ;
			data[100009] <= 8'h10 ;
			data[100010] <= 8'h10 ;
			data[100011] <= 8'h10 ;
			data[100012] <= 8'h10 ;
			data[100013] <= 8'h10 ;
			data[100014] <= 8'h10 ;
			data[100015] <= 8'h10 ;
			data[100016] <= 8'h10 ;
			data[100017] <= 8'h10 ;
			data[100018] <= 8'h10 ;
			data[100019] <= 8'h10 ;
			data[100020] <= 8'h10 ;
			data[100021] <= 8'h10 ;
			data[100022] <= 8'h10 ;
			data[100023] <= 8'h10 ;
			data[100024] <= 8'h10 ;
			data[100025] <= 8'h10 ;
			data[100026] <= 8'h10 ;
			data[100027] <= 8'h10 ;
			data[100028] <= 8'h10 ;
			data[100029] <= 8'h10 ;
			data[100030] <= 8'h10 ;
			data[100031] <= 8'h10 ;
			data[100032] <= 8'h10 ;
			data[100033] <= 8'h10 ;
			data[100034] <= 8'h10 ;
			data[100035] <= 8'h10 ;
			data[100036] <= 8'h10 ;
			data[100037] <= 8'h10 ;
			data[100038] <= 8'h10 ;
			data[100039] <= 8'h10 ;
			data[100040] <= 8'h10 ;
			data[100041] <= 8'h10 ;
			data[100042] <= 8'h10 ;
			data[100043] <= 8'h10 ;
			data[100044] <= 8'h10 ;
			data[100045] <= 8'h10 ;
			data[100046] <= 8'h10 ;
			data[100047] <= 8'h10 ;
			data[100048] <= 8'h10 ;
			data[100049] <= 8'h10 ;
			data[100050] <= 8'h10 ;
			data[100051] <= 8'h10 ;
			data[100052] <= 8'h10 ;
			data[100053] <= 8'h10 ;
			data[100054] <= 8'h10 ;
			data[100055] <= 8'h10 ;
			data[100056] <= 8'h10 ;
			data[100057] <= 8'h10 ;
			data[100058] <= 8'h10 ;
			data[100059] <= 8'h10 ;
			data[100060] <= 8'h10 ;
			data[100061] <= 8'h10 ;
			data[100062] <= 8'h10 ;
			data[100063] <= 8'h10 ;
			data[100064] <= 8'h10 ;
			data[100065] <= 8'h10 ;
			data[100066] <= 8'h10 ;
			data[100067] <= 8'h10 ;
			data[100068] <= 8'h10 ;
			data[100069] <= 8'h10 ;
			data[100070] <= 8'h10 ;
			data[100071] <= 8'h10 ;
			data[100072] <= 8'h10 ;
			data[100073] <= 8'h10 ;
			data[100074] <= 8'h10 ;
			data[100075] <= 8'h10 ;
			data[100076] <= 8'h10 ;
			data[100077] <= 8'h10 ;
			data[100078] <= 8'h10 ;
			data[100079] <= 8'h10 ;
			data[100080] <= 8'h10 ;
			data[100081] <= 8'h10 ;
			data[100082] <= 8'h10 ;
			data[100083] <= 8'h10 ;
			data[100084] <= 8'h10 ;
			data[100085] <= 8'h10 ;
			data[100086] <= 8'h10 ;
			data[100087] <= 8'h10 ;
			data[100088] <= 8'h10 ;
			data[100089] <= 8'h10 ;
			data[100090] <= 8'h10 ;
			data[100091] <= 8'h10 ;
			data[100092] <= 8'h10 ;
			data[100093] <= 8'h10 ;
			data[100094] <= 8'h10 ;
			data[100095] <= 8'h10 ;
			data[100096] <= 8'h10 ;
			data[100097] <= 8'h10 ;
			data[100098] <= 8'h10 ;
			data[100099] <= 8'h10 ;
			data[100100] <= 8'h10 ;
			data[100101] <= 8'h10 ;
			data[100102] <= 8'h10 ;
			data[100103] <= 8'h10 ;
			data[100104] <= 8'h10 ;
			data[100105] <= 8'h10 ;
			data[100106] <= 8'h10 ;
			data[100107] <= 8'h10 ;
			data[100108] <= 8'h10 ;
			data[100109] <= 8'h10 ;
			data[100110] <= 8'h10 ;
			data[100111] <= 8'h10 ;
			data[100112] <= 8'h10 ;
			data[100113] <= 8'h10 ;
			data[100114] <= 8'h10 ;
			data[100115] <= 8'h10 ;
			data[100116] <= 8'h10 ;
			data[100117] <= 8'h10 ;
			data[100118] <= 8'h10 ;
			data[100119] <= 8'h10 ;
			data[100120] <= 8'h10 ;
			data[100121] <= 8'h10 ;
			data[100122] <= 8'h10 ;
			data[100123] <= 8'h10 ;
			data[100124] <= 8'h10 ;
			data[100125] <= 8'h10 ;
			data[100126] <= 8'h10 ;
			data[100127] <= 8'h10 ;
			data[100128] <= 8'h10 ;
			data[100129] <= 8'h10 ;
			data[100130] <= 8'h10 ;
			data[100131] <= 8'h10 ;
			data[100132] <= 8'h10 ;
			data[100133] <= 8'h10 ;
			data[100134] <= 8'h10 ;
			data[100135] <= 8'h10 ;
			data[100136] <= 8'h10 ;
			data[100137] <= 8'h10 ;
			data[100138] <= 8'h10 ;
			data[100139] <= 8'h10 ;
			data[100140] <= 8'h10 ;
			data[100141] <= 8'h10 ;
			data[100142] <= 8'h10 ;
			data[100143] <= 8'h10 ;
			data[100144] <= 8'h10 ;
			data[100145] <= 8'h10 ;
			data[100146] <= 8'h10 ;
			data[100147] <= 8'h10 ;
			data[100148] <= 8'h10 ;
			data[100149] <= 8'h10 ;
			data[100150] <= 8'h10 ;
			data[100151] <= 8'h10 ;
			data[100152] <= 8'h10 ;
			data[100153] <= 8'h10 ;
			data[100154] <= 8'h10 ;
			data[100155] <= 8'h10 ;
			data[100156] <= 8'h10 ;
			data[100157] <= 8'h10 ;
			data[100158] <= 8'h10 ;
			data[100159] <= 8'h10 ;
			data[100160] <= 8'h10 ;
			data[100161] <= 8'h10 ;
			data[100162] <= 8'h10 ;
			data[100163] <= 8'h10 ;
			data[100164] <= 8'h10 ;
			data[100165] <= 8'h10 ;
			data[100166] <= 8'h10 ;
			data[100167] <= 8'h10 ;
			data[100168] <= 8'h10 ;
			data[100169] <= 8'h10 ;
			data[100170] <= 8'h10 ;
			data[100171] <= 8'h10 ;
			data[100172] <= 8'h10 ;
			data[100173] <= 8'h10 ;
			data[100174] <= 8'h10 ;
			data[100175] <= 8'h10 ;
			data[100176] <= 8'h10 ;
			data[100177] <= 8'h10 ;
			data[100178] <= 8'h10 ;
			data[100179] <= 8'h10 ;
			data[100180] <= 8'h10 ;
			data[100181] <= 8'h10 ;
			data[100182] <= 8'h10 ;
			data[100183] <= 8'h10 ;
			data[100184] <= 8'h10 ;
			data[100185] <= 8'h10 ;
			data[100186] <= 8'h10 ;
			data[100187] <= 8'h10 ;
			data[100188] <= 8'h10 ;
			data[100189] <= 8'h10 ;
			data[100190] <= 8'h10 ;
			data[100191] <= 8'h10 ;
			data[100192] <= 8'h10 ;
			data[100193] <= 8'h10 ;
			data[100194] <= 8'h10 ;
			data[100195] <= 8'h10 ;
			data[100196] <= 8'h10 ;
			data[100197] <= 8'h10 ;
			data[100198] <= 8'h10 ;
			data[100199] <= 8'h10 ;
			data[100200] <= 8'h10 ;
			data[100201] <= 8'h10 ;
			data[100202] <= 8'h10 ;
			data[100203] <= 8'h10 ;
			data[100204] <= 8'h10 ;
			data[100205] <= 8'h10 ;
			data[100206] <= 8'h10 ;
			data[100207] <= 8'h10 ;
			data[100208] <= 8'h10 ;
			data[100209] <= 8'h10 ;
			data[100210] <= 8'h10 ;
			data[100211] <= 8'h10 ;
			data[100212] <= 8'h10 ;
			data[100213] <= 8'h10 ;
			data[100214] <= 8'h10 ;
			data[100215] <= 8'h10 ;
			data[100216] <= 8'h10 ;
			data[100217] <= 8'h10 ;
			data[100218] <= 8'h10 ;
			data[100219] <= 8'h10 ;
			data[100220] <= 8'h10 ;
			data[100221] <= 8'h10 ;
			data[100222] <= 8'h10 ;
			data[100223] <= 8'h10 ;
			data[100224] <= 8'h10 ;
			data[100225] <= 8'h10 ;
			data[100226] <= 8'h10 ;
			data[100227] <= 8'h10 ;
			data[100228] <= 8'h10 ;
			data[100229] <= 8'h10 ;
			data[100230] <= 8'h10 ;
			data[100231] <= 8'h10 ;
			data[100232] <= 8'h10 ;
			data[100233] <= 8'h10 ;
			data[100234] <= 8'h10 ;
			data[100235] <= 8'h10 ;
			data[100236] <= 8'h10 ;
			data[100237] <= 8'h10 ;
			data[100238] <= 8'h10 ;
			data[100239] <= 8'h10 ;
			data[100240] <= 8'h10 ;
			data[100241] <= 8'h10 ;
			data[100242] <= 8'h10 ;
			data[100243] <= 8'h10 ;
			data[100244] <= 8'h10 ;
			data[100245] <= 8'h10 ;
			data[100246] <= 8'h10 ;
			data[100247] <= 8'h10 ;
			data[100248] <= 8'h10 ;
			data[100249] <= 8'h10 ;
			data[100250] <= 8'h10 ;
			data[100251] <= 8'h10 ;
			data[100252] <= 8'h10 ;
			data[100253] <= 8'h10 ;
			data[100254] <= 8'h10 ;
			data[100255] <= 8'h10 ;
			data[100256] <= 8'h10 ;
			data[100257] <= 8'h10 ;
			data[100258] <= 8'h10 ;
			data[100259] <= 8'h10 ;
			data[100260] <= 8'h10 ;
			data[100261] <= 8'h10 ;
			data[100262] <= 8'h10 ;
			data[100263] <= 8'h10 ;
			data[100264] <= 8'h10 ;
			data[100265] <= 8'h10 ;
			data[100266] <= 8'h10 ;
			data[100267] <= 8'h10 ;
			data[100268] <= 8'h10 ;
			data[100269] <= 8'h10 ;
			data[100270] <= 8'h10 ;
			data[100271] <= 8'h10 ;
			data[100272] <= 8'h10 ;
			data[100273] <= 8'h10 ;
			data[100274] <= 8'h10 ;
			data[100275] <= 8'h10 ;
			data[100276] <= 8'h10 ;
			data[100277] <= 8'h10 ;
			data[100278] <= 8'h10 ;
			data[100279] <= 8'h10 ;
			data[100280] <= 8'h10 ;
			data[100281] <= 8'h10 ;
			data[100282] <= 8'h10 ;
			data[100283] <= 8'h10 ;
			data[100284] <= 8'h10 ;
			data[100285] <= 8'h10 ;
			data[100286] <= 8'h10 ;
			data[100287] <= 8'h10 ;
			data[100288] <= 8'h10 ;
			data[100289] <= 8'h10 ;
			data[100290] <= 8'h10 ;
			data[100291] <= 8'h10 ;
			data[100292] <= 8'h10 ;
			data[100293] <= 8'h10 ;
			data[100294] <= 8'h10 ;
			data[100295] <= 8'h10 ;
			data[100296] <= 8'h10 ;
			data[100297] <= 8'h10 ;
			data[100298] <= 8'h10 ;
			data[100299] <= 8'h10 ;
			data[100300] <= 8'h10 ;
			data[100301] <= 8'h10 ;
		end
		
		if ( enRead )
		begin
			dataOUT1 <= data[addr] ;
			dataOUT2 <= data[addr+1] ;
			dataOUT3 <= data[addr+2] ;
			dataOUT4 <= data[addr+3] ;
			dataOUT5 <= data[addr+4] ;
			dataOUT6 <= data[addr+5] ;
			dataOUT7 <= data[addr+6] ;
			dataOUT8 <= data[addr+7] ;
			dataOUT9 <= data[addr+8] ;
			dataOUT10 <= data[addr+9] ;
			dataOUT11 <= data[addr+10] ;
			dataOUT12 <= data[addr+11] ;
			dataOUT13 <= data[addr+12] ;
			dataOUT14 <= data[addr+13] ;
			dataOUT15 <= data[addr+14] ;
			dataOUT16 <= data[addr+15] ;
			dataOUT17 <= data[addr+16] ;
			dataOUT18 <= data[addr+17] ;
			dataOUT19 <= data[addr+18] ;
			dataOUT20 <= data[addr+19] ;
			dataOUT21 <= data[addr+20] ;
			dataOUT22 <= data[addr+21] ;
			dataOUT23 <= data[addr+22] ;
			dataOUT24 <= data[addr+23] ;
			dataOUT25 <= data[addr+24] ;
			dataOUT26 <= data[addr+25] ;
			dataOUT27 <= data[addr+26] ;
			dataOUT28 <= data[addr+27] ;
			dataOUT29 <= data[addr+28] ;
			dataOUT30 <= data[addr+29] ;
			dataOUT31 <= data[addr+30] ;
			dataOUT32 <= data[addr+31] ;
			dataOUT33 <= data[addr+32] ;
			dataOUT34 <= data[addr+33] ;
			dataOUT35 <= data[addr+34] ;
			dataOUT36 <= data[addr+35] ;
			dataOUT37 <= data[addr+36] ;
			dataOUT38 <= data[addr+37] ;
			dataOUT39 <= data[addr+38] ;
			dataOUT40 <= data[addr+39] ;
			dataOUT41 <= data[addr+40] ;
			dataOUT42 <= data[addr+41] ;
			dataOUT43 <= data[addr+42] ;
			dataOUT44 <= data[addr+43] ;
			dataOUT45 <= data[addr+44] ;
			dataOUT46 <= data[addr+45] ;
			dataOUT47 <= data[addr+46] ;
			dataOUT48 <= data[addr+47] ;
			dataOUT49 <= data[addr+48] ;
			dataOUT50 <= data[addr+49] ;
		end 
		else 
		begin 
			dataOUT1 <= 8'hzz ;
			dataOUT2 <= 8'hzz ;
			dataOUT3 <= 8'hzz ;
			dataOUT4 <= 8'hzz ;
			dataOUT5 <= 8'hzz ;
			dataOUT6 <= 8'hzz ;
			dataOUT7 <= 8'hzz ;
			dataOUT8 <= 8'hzz ;
			dataOUT9 <= 8'hzz ;
			dataOUT10 <= 8'hzz ;
			dataOUT11 <= 8'hzz ;
			dataOUT12 <= 8'hzz ;
			dataOUT13 <= 8'hzz ;
			dataOUT14 <= 8'hzz ;
			dataOUT15 <= 8'hzz ;
			dataOUT16 <= 8'hzz ;
			dataOUT17 <= 8'hzz ;
			dataOUT18 <= 8'hzz ;
			dataOUT19 <= 8'hzz ;
			dataOUT20 <= 8'hzz ;
			dataOUT21 <= 8'hzz ;
			dataOUT22 <= 8'hzz ;
			dataOUT23 <= 8'hzz ;
			dataOUT24 <= 8'hzz ;
			dataOUT25 <= 8'hzz ;
			dataOUT26 <= 8'hzz ;
			dataOUT27 <= 8'hzz ;
			dataOUT28 <= 8'hzz ;
			dataOUT29 <= 8'hzz ;
			dataOUT30 <= 8'hzz ;
			dataOUT31 <= 8'hzz ;
			dataOUT32 <= 8'hzz ;
			dataOUT33 <= 8'hzz ;
			dataOUT34 <= 8'hzz ;
			dataOUT35 <= 8'hzz ;
			dataOUT36 <= 8'hzz ;
			dataOUT37 <= 8'hzz ;
			dataOUT38 <= 8'hzz ;
			dataOUT39 <= 8'hzz ;
			dataOUT40 <= 8'hzz ;
			dataOUT41 <= 8'hzz ;
			dataOUT42 <= 8'hzz ;
			dataOUT43 <= 8'hzz ;
			dataOUT44 <= 8'hzz ;
			dataOUT45 <= 8'hzz ;
			dataOUT46 <= 8'hzz ;
			dataOUT47 <= 8'hzz ;
			dataOUT48 <= 8'hzz ;
			dataOUT49 <= 8'hzz ;
			dataOUT50 <= 8'hzz ;
		end 
	end 
   
endmodule