`timescale 1ns/10ps

module nnctrl50_tb ;
	reg clock, reset ;
	reg [7:0] in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19,  in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50 ;

	nnctrl50 t ( reset, clock, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19,  in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50 ) ;

	initial // reset、clock
	begin
		clock = 0 ;
		reset = 0 ;
		#100
		reset = 1 ;
		#100
		reset = 0 ;
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h01 ; in2 = 8'h01 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h00 ; in2 = 8'h00 ; in3 = 8'h01 ; in4 = 8'h01 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
		#200 begin 
			in1 = 8'h10 ; in2 = 8'h00 ; in3 = 8'h00 ; in4 = 8'h00 ; in5 = 8'h00 ; in6 = 8'h00 ; in7 = 8'h00 ; in8 = 8'h00 ; in9 = 8'h00 ; in10 = 8'h00 ; in11 = 8'h00 ; in12 = 8'h00 ; in13 = 8'h00 ; in14 = 8'h00 ; in15 = 8'h00 ; in16 = 8'h00 ; in17 = 8'h00 ; in18 = 8'h00 ; in19 = 8'h00 ;  in20 = 8'h00 ; in21 = 8'h00 ; in22 = 8'h00 ; in23 = 8'h00 ; in24 = 8'h00 ; in25 = 8'h00 ; in26 = 8'h00 ; in27 = 8'h00 ; in28 = 8'h00 ; in29 = 8'h00 ; in30 = 8'h00 ; in31 = 8'h00 ; in32 = 8'h00 ; in33 = 8'h00 ; in34 = 8'h00 ; in35 = 8'h00 ; in36 = 8'h00 ; in37 = 8'h00 ; in38 = 8'h00 ; in39 = 8'h00 ; in40 = 8'h00 ; in41 = 8'h00 ; in42 = 8'h00 ; in43 = 8'h00 ; in44 = 8'h00 ; in45 = 8'h00 ; in46 = 8'h00 ; in47 = 8'h00 ; in48 = 8'h00 ; in49 = 8'h00 ; in50 = 8'h00 ;
		end
	end
	always #100 clock = clock + 1; 


endmodule